module pre_norm_addsub_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [7:0] A ;
input [7:0] B ;
output [7:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire [8:0] carry ;
// instances
  FADDX1 U2_6(.A(A[6:6]),.B(n3),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n4),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n5),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n6),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n7),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n8),.CI(n1),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_7(.IN1(A[7:7]),.IN2(n2),.IN3(carry[7:7]),.Q(DIFF[7:7]));
  INVX0 U1(.INP(B[1:1]),.ZN(n8));
  INVX0 U2(.INP(B[2:2]),.ZN(n7));
  INVX0 U3(.INP(B[3:3]),.ZN(n6));
  AND2X1 U4(.IN1(A[0:0]),.IN2(n9),.Q(n1));
  INVX0 U5(.INP(B[4:4]),.ZN(n5));
  INVX0 U6(.INP(B[5:5]),.ZN(n4));
  INVX0 U7(.INP(B[6:6]),.ZN(n3));
  INVX0 U8(.INP(B[0:0]),.ZN(n9));
  INVX0 U9(.INP(B[7:7]),.ZN(n2));
  XOR2X1 U10(.IN1(A[0:0]),.IN2(n9),.Q(DIFF[0:0]));
endmodule
module pre_norm_addsub_DW01_sub_1_inj (A,B,CI,DIFF,CO);
input [7:0] A ;
input [7:0] B ;
output [7:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire [8:0] carry ;
// instances
  FADDX1 U2_6(.A(A[6:6]),.B(n4),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n5),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n6),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n7),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n8),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n9),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_7(.IN1(A[7:7]),.IN2(n3),.IN3(carry[7:7]),.Q(DIFF[7:7]));
  INVX0 U1(.INP(B[2:2]),.ZN(n8));
  INVX0 U2(.INP(B[3:3]),.ZN(n7));
  INVX0 U3(.INP(B[1:1]),.ZN(n9));
  NAND2X1 U4(.IN1(n1),.IN2(n2),.QN(carry[1:1]));
  INVX0 U5(.INP(A[0:0]),.ZN(n1));
  INVX0 U6(.INP(B[4:4]),.ZN(n6));
  INVX0 U7(.INP(B[5:5]),.ZN(n5));
  INVX0 U8(.INP(B[6:6]),.ZN(n4));
  INVX0 U9(.INP(n10),.ZN(n2));
  INVX0 U10(.INP(B[0:0]),.ZN(n10));
  INVX0 U11(.INP(B[7:7]),.ZN(n3));
  XOR2X1 U12(.IN1(n2),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module pre_norm_addsub_DW01_sub_2_inj (A,B,CI,DIFF,CO);
input [7:0] A ;
input [7:0] B ;
output [7:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire [8:0] carry ;
// instances
  FADDX1 U2_6(.A(A[6:6]),.B(n3),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n5),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n6),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n7),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n8),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n9),.CI(n1),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_7(.IN1(A[7:7]),.IN2(n4),.IN3(carry[7:7]),.Q(DIFF[7:7]));
  INVX0 U1(.INP(B[1:1]),.ZN(n9));
  INVX0 U2(.INP(B[2:2]),.ZN(n8));
  INVX0 U3(.INP(B[3:3]),.ZN(n7));
  AND2X1 U4(.IN1(A[0:0]),.IN2(n2),.Q(n1));
  INVX0 U5(.INP(B[5:5]),.ZN(n5));
  INVX0 U6(.INP(B[4:4]),.ZN(n6));
  XOR2X1 U7(.IN1(A[0:0]),.IN2(n2),.Q(DIFF[0:0]));
  INVX0 U8(.INP(B[0:0]),.ZN(n2));
  INVX0 U9(.INP(B[6:6]),.ZN(n3));
  INVX0 U10(.INP(B[7:7]),.ZN(n4));
endmodule
module pre_norm_addsub_DW01_sub_3_inj (A,B,CI,DIFF,CO);
input [7:0] A ;
input [7:0] B ;
output [7:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire [8:0] carry ;
// instances
  FADDX1 U2_6(.A(A[6:6]),.B(n4),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n6),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n7),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n8),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n9),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n10),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_7(.IN1(A[7:7]),.IN2(n5),.IN3(carry[7:7]),.Q(DIFF[7:7]));
  INVX0 U1(.INP(n3),.ZN(n2));
  INVX0 U2(.INP(B[2:2]),.ZN(n9));
  INVX0 U3(.INP(B[3:3]),.ZN(n8));
  NAND2X1 U4(.IN1(n1),.IN2(n2),.QN(carry[1:1]));
  INVX0 U5(.INP(B[1:1]),.ZN(n10));
  INVX0 U6(.INP(A[0:0]),.ZN(n1));
  INVX0 U7(.INP(B[5:5]),.ZN(n6));
  INVX0 U8(.INP(B[4:4]),.ZN(n7));
  XOR2X1 U9(.IN1(n2),.IN2(A[0:0]),.Q(DIFF[0:0]));
  INVX0 U10(.INP(B[0:0]),.ZN(n3));
  INVX0 U11(.INP(B[6:6]),.ZN(n4));
  INVX0 U12(.INP(B[7:7]),.ZN(n5));
endmodule
module pre_norm_addsub_inj (clk_i,opa_i,opb_i,fracta_28_o,fractb_28_o,exp_o);
input [31:0] opa_i ;
input [31:0] opb_i ;
output [27:0] fracta_28_o ;
output [27:0] fractb_28_o ;
output [7:0] exp_o ;
input clk_i ;
wire N109 ;
wire N124 ;
wire N125 ;
wire N126 ;
wire N127 ;
wire N128 ;
wire N129 ;
wire N130 ;
wire N131 ;
wire N139 ;
wire N140 ;
wire N141 ;
wire N142 ;
wire N143 ;
wire N144 ;
wire N145 ;
wire N146 ;
wire N155 ;
wire N156 ;
wire N157 ;
wire N158 ;
wire N159 ;
wire N160 ;
wire N161 ;
wire N162 ;
wire N163 ;
wire N164 ;
wire N165 ;
wire N166 ;
wire N167 ;
wire N168 ;
wire N169 ;
wire N170 ;
wire N179 ;
wire N180 ;
wire N181 ;
wire N182 ;
wire N183 ;
wire N184 ;
wire N185 ;
wire N186 ;
wire N187 ;
wire N188 ;
wire N189 ;
wire N190 ;
wire N191 ;
wire N192 ;
wire N193 ;
wire N194 ;
wire N231 ;
wire N236 ;
wire N238 ;
wire N246 ;
wire N247 ;
wire N248 ;
wire N249 ;
wire N252 ;
wire N253 ;
wire N254 ;
wire N263 ;
wire N264 ;
wire N265 ;
wire N266 ;
wire N267 ;
wire N269 ;
wire N270 ;
wire N271 ;
wire N272 ;
wire N280 ;
wire N281 ;
wire N282 ;
wire N283 ;
wire N284 ;
wire N285 ;
wire N286 ;
wire N287 ;
wire N288 ;
wire N289 ;
wire N290 ;
wire N297 ;
wire N298 ;
wire N299 ;
wire N300 ;
wire N301 ;
wire N302 ;
wire N303 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N308 ;
wire N314 ;
wire N315 ;
wire N316 ;
wire N317 ;
wire N318 ;
wire N319 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N324 ;
wire N325 ;
wire N331 ;
wire N332 ;
wire N333 ;
wire N334 ;
wire N335 ;
wire N336 ;
wire N337 ;
wire N338 ;
wire N339 ;
wire N340 ;
wire N341 ;
wire N342 ;
wire N348 ;
wire N349 ;
wire N350 ;
wire N351 ;
wire N352 ;
wire N353 ;
wire N354 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N365 ;
wire N366 ;
wire N367 ;
wire N368 ;
wire N369 ;
wire N370 ;
wire N371 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N382 ;
wire N383 ;
wire N384 ;
wire N385 ;
wire N386 ;
wire N387 ;
wire N388 ;
wire N389 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N399 ;
wire N400 ;
wire N401 ;
wire N402 ;
wire N403 ;
wire N404 ;
wire N405 ;
wire N406 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N416 ;
wire N417 ;
wire N418 ;
wire N419 ;
wire N420 ;
wire N421 ;
wire N422 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N433 ;
wire N434 ;
wire N435 ;
wire N436 ;
wire N437 ;
wire N438 ;
wire N439 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N450 ;
wire N451 ;
wire N452 ;
wire N453 ;
wire N454 ;
wire N455 ;
wire N456 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N467 ;
wire N468 ;
wire N469 ;
wire N470 ;
wire N471 ;
wire N472 ;
wire N473 ;
wire N474 ;
wire N475 ;
wire N476 ;
wire N477 ;
wire N478 ;
wire N484 ;
wire N485 ;
wire N486 ;
wire N487 ;
wire N488 ;
wire N489 ;
wire N490 ;
wire N491 ;
wire N492 ;
wire N493 ;
wire N494 ;
wire N495 ;
wire N501 ;
wire N502 ;
wire N503 ;
wire N504 ;
wire N505 ;
wire N506 ;
wire N507 ;
wire N508 ;
wire N509 ;
wire N510 ;
wire N511 ;
wire N512 ;
wire N518 ;
wire N519 ;
wire N520 ;
wire N521 ;
wire N522 ;
wire N523 ;
wire N524 ;
wire N525 ;
wire N526 ;
wire N527 ;
wire N528 ;
wire N529 ;
wire N535 ;
wire N536 ;
wire N537 ;
wire N538 ;
wire N539 ;
wire N540 ;
wire N541 ;
wire N542 ;
wire N543 ;
wire N544 ;
wire N545 ;
wire N546 ;
wire N552 ;
wire N553 ;
wire N554 ;
wire N555 ;
wire N556 ;
wire N557 ;
wire N558 ;
wire N559 ;
wire N560 ;
wire N561 ;
wire N562 ;
wire N563 ;
wire N569 ;
wire N570 ;
wire N571 ;
wire N572 ;
wire N573 ;
wire N574 ;
wire N575 ;
wire N576 ;
wire N577 ;
wire N578 ;
wire N579 ;
wire N580 ;
wire N586 ;
wire N587 ;
wire N588 ;
wire N589 ;
wire N590 ;
wire N591 ;
wire N592 ;
wire N593 ;
wire N594 ;
wire N595 ;
wire N596 ;
wire N597 ;
wire N603 ;
wire N604 ;
wire N605 ;
wire N606 ;
wire N607 ;
wire N608 ;
wire N609 ;
wire N610 ;
wire N611 ;
wire N612 ;
wire N613 ;
wire N614 ;
wire N619 ;
wire N620 ;
wire N621 ;
wire N622 ;
wire N623 ;
wire N624 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire \add_105_I28_L14036_C161/carry[5]  ;
wire \add_105_I28_L14036_C161/carry[4]  ;
wire \add_105_I28_L14036_C161/carry[3]  ;
wire \add_105_I28_L14036_C161/carry[2]  ;
wire \add_105_I27_L14036_C161/carry[5]  ;
wire \add_105_I27_L14036_C161/carry[4]  ;
wire \add_105_I27_L14036_C161/carry[3]  ;
wire \add_105_I27_L14036_C161/carry[2]  ;
wire \add_105_I26_L14036_C161/carry[5]  ;
wire \add_105_I26_L14036_C161/carry[4]  ;
wire \add_105_I26_L14036_C161/carry[3]  ;
wire \add_105_I26_L14036_C161/carry[2]  ;
wire \add_105_I25_L14036_C161/carry[5]  ;
wire \add_105_I25_L14036_C161/carry[4]  ;
wire \add_105_I25_L14036_C161/carry[3]  ;
wire \add_105_I25_L14036_C161/carry[2]  ;
wire \add_105_I24_L14036_C161/carry[5]  ;
wire \add_105_I24_L14036_C161/carry[4]  ;
wire \add_105_I24_L14036_C161/carry[3]  ;
wire \add_105_I24_L14036_C161/carry[2]  ;
wire \add_105_I23_L14036_C161/carry[5]  ;
wire \add_105_I23_L14036_C161/carry[4]  ;
wire \add_105_I23_L14036_C161/carry[3]  ;
wire \add_105_I23_L14036_C161/carry[2]  ;
wire \add_105_I22_L14036_C161/carry[5]  ;
wire \add_105_I22_L14036_C161/carry[4]  ;
wire \add_105_I22_L14036_C161/carry[3]  ;
wire \add_105_I22_L14036_C161/carry[2]  ;
wire \add_105_I21_L14036_C161/carry[5]  ;
wire \add_105_I21_L14036_C161/carry[4]  ;
wire \add_105_I21_L14036_C161/carry[3]  ;
wire \add_105_I21_L14036_C161/carry[2]  ;
wire \add_105_I20_L14036_C161/carry[5]  ;
wire \add_105_I20_L14036_C161/carry[4]  ;
wire \add_105_I20_L14036_C161/carry[3]  ;
wire \add_105_I20_L14036_C161/carry[2]  ;
wire \add_105_I19_L14036_C161/carry[5]  ;
wire \add_105_I19_L14036_C161/carry[4]  ;
wire \add_105_I19_L14036_C161/carry[3]  ;
wire \add_105_I19_L14036_C161/carry[2]  ;
wire \add_105_I18_L14036_C161/carry[5]  ;
wire \add_105_I18_L14036_C161/carry[4]  ;
wire \add_105_I18_L14036_C161/carry[3]  ;
wire \add_105_I18_L14036_C161/carry[2]  ;
wire \add_105_I17_L14036_C161/carry[5]  ;
wire \add_105_I17_L14036_C161/carry[4]  ;
wire \add_105_I17_L14036_C161/carry[3]  ;
wire \add_105_I17_L14036_C161/carry[2]  ;
wire \add_105_I16_L14036_C161/carry[5]  ;
wire \add_105_I16_L14036_C161/carry[4]  ;
wire \add_105_I16_L14036_C161/carry[3]  ;
wire \add_105_I16_L14036_C161/carry[2]  ;
wire \add_105_I15_L14036_C161/carry[5]  ;
wire \add_105_I15_L14036_C161/carry[4]  ;
wire \add_105_I15_L14036_C161/carry[3]  ;
wire \add_105_I15_L14036_C161/carry[2]  ;
wire \add_105_I14_L14036_C161/carry[5]  ;
wire \add_105_I14_L14036_C161/carry[4]  ;
wire \add_105_I14_L14036_C161/carry[3]  ;
wire \add_105_I14_L14036_C161/carry[2]  ;
wire \add_105_I13_L14036_C161/carry[5]  ;
wire \add_105_I13_L14036_C161/carry[4]  ;
wire \add_105_I13_L14036_C161/carry[3]  ;
wire \add_105_I13_L14036_C161/carry[2]  ;
wire \add_105_I12_L14036_C161/carry[5]  ;
wire \add_105_I12_L14036_C161/carry[4]  ;
wire \add_105_I12_L14036_C161/carry[3]  ;
wire \add_105_I12_L14036_C161/carry[2]  ;
wire \add_105_I11_L14036_C161/carry[5]  ;
wire \add_105_I11_L14036_C161/carry[4]  ;
wire \add_105_I11_L14036_C161/carry[3]  ;
wire \add_105_I11_L14036_C161/carry[2]  ;
wire \add_105_I10_L14036_C161/carry[5]  ;
wire \add_105_I10_L14036_C161/carry[4]  ;
wire \add_105_I10_L14036_C161/carry[3]  ;
wire \add_105_I10_L14036_C161/carry[2]  ;
wire \add_105_I9_L14036_C161/carry[5]  ;
wire \add_105_I9_L14036_C161/carry[4]  ;
wire \add_105_I9_L14036_C161/carry[3]  ;
wire \add_105_I9_L14036_C161/carry[2]  ;
wire \add_105_I8_L14036_C161/carry[4]  ;
wire \add_105_I8_L14036_C161/carry[3]  ;
wire \add_105_I8_L14036_C161/carry[2]  ;
wire \add_105_I7_L14036_C161/carry[2]  ;
wire \add_105_I7_L14036_C161/carry[3]  ;
wire \add_105_I6_L14036_C161/carry[2]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n152 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n381 ;
wire n382 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n404 ;
wire n405 ;
wire n406 ;
wire n407 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n416 ;
wire n417 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire [7:0] s_exp_o ;
wire [26:0] s_fracta_28_o ;
wire [26:0] s_fractb_28_o ;
wire [7:0] s_exp_diff ;
wire [26:3] s_fract_sm_28 ;
wire [26:0] s_fract_shr_28 ;
wire [5:0] s_rzeros ;
// instances
  DFFX1 desc0(.D(N131),.CLK(clk_i),.Q(s_exp_o[7:7]));
  DFFX1 desc1(.D(s_exp_o[7:7]),.CLK(clk_i),.Q(exp_o[7:7]));
  DFFX1 desc2(.D(N130),.CLK(clk_i),.Q(s_exp_o[6:6]));
  DFFX1 desc3(.D(s_exp_o[6:6]),.CLK(clk_i),.Q(exp_o[6:6]));
  DFFX1 desc4(.D(N129),.CLK(clk_i),.Q(s_exp_o[5:5]));
  DFFX1 desc5(.D(s_exp_o[5:5]),.CLK(clk_i),.Q(exp_o[5:5]));
  DFFX1 desc6(.D(N128),.CLK(clk_i),.Q(s_exp_o[4:4]));
  DFFX1 desc7(.D(s_exp_o[4:4]),.CLK(clk_i),.Q(exp_o[4:4]));
  DFFX1 desc8(.D(N127),.CLK(clk_i),.Q(s_exp_o[3:3]));
  DFFX1 desc9(.D(s_exp_o[3:3]),.CLK(clk_i),.Q(exp_o[3:3]));
  DFFX1 desc10(.D(N126),.CLK(clk_i),.Q(s_exp_o[2:2]));
  DFFX1 desc11(.D(s_exp_o[2:2]),.CLK(clk_i),.Q(exp_o[2:2]));
  DFFX1 desc12(.D(N125),.CLK(clk_i),.Q(s_exp_o[1:1]));
  DFFX1 desc13(.D(s_exp_o[1:1]),.CLK(clk_i),.Q(exp_o[1:1]));
  DFFX1 desc14(.D(N124),.CLK(clk_i),.Q(s_exp_o[0:0]));
  DFFX1 desc15(.D(s_exp_o[0:0]),.CLK(clk_i),.Q(exp_o[0:0]));
  DFFX1 desc16(.D(N194),.CLK(clk_i),.Q(s_exp_diff[7:7]));
  DFFX1 desc17(.D(N193),.CLK(clk_i),.Q(s_exp_diff[6:6]));
  DFFX1 desc18(.D(N192),.CLK(clk_i),.Q(s_exp_diff[5:5]));
  DFFX1 desc19(.D(N191),.CLK(clk_i),.Q(s_exp_diff[4:4]));
  DFFX1 desc20(.D(N190),.CLK(clk_i),.Q(s_exp_diff[3:3]),.QN(n2));
  DFFX1 desc21(.D(N189),.CLK(clk_i),.Q(s_exp_diff[2:2]),.QN(n5));
  DFFX1 desc22(.D(N188),.CLK(clk_i),.Q(s_exp_diff[1:1]),.QN(n4));
  DFFX1 desc23(.D(N187),.CLK(clk_i),.Q(s_exp_diff[0:0]),.QN(n3));
  DFFSSRX1 desc24(.D(n46),.RSTB(s_fract_shr_28[1:1]),.SETB(1'b1),.CLK(clk_i),.Q(fractb_28_o[1:1]));
  DFFSSRX1 desc25(.D(n32),.RSTB(s_fract_shr_28[1:1]),.SETB(1'b1),.CLK(clk_i),.Q(fracta_28_o[1:1]));
  DFFSSRX1 desc26(.D(n46),.RSTB(s_fract_shr_28[2:2]),.SETB(1'b1),.CLK(clk_i),.Q(fractb_28_o[2:2]));
  DFFSSRX1 desc27(.D(n32),.RSTB(s_fract_shr_28[2:2]),.SETB(1'b1),.CLK(clk_i),.Q(fracta_28_o[2:2]));
  DFFX1 desc28(.D(s_fracta_28_o[3:3]),.CLK(clk_i),.Q(fracta_28_o[3:3]));
  DFFX1 desc29(.D(s_fractb_28_o[3:3]),.CLK(clk_i),.Q(fractb_28_o[3:3]));
  DFFX1 desc30(.D(s_fracta_28_o[4:4]),.CLK(clk_i),.Q(fracta_28_o[4:4]));
  DFFX1 desc31(.D(s_fractb_28_o[4:4]),.CLK(clk_i),.Q(fractb_28_o[4:4]));
  DFFX1 desc32(.D(s_fracta_28_o[5:5]),.CLK(clk_i),.Q(fracta_28_o[5:5]));
  DFFX1 desc33(.D(s_fractb_28_o[5:5]),.CLK(clk_i),.Q(fractb_28_o[5:5]));
  DFFX1 desc34(.D(s_fracta_28_o[6:6]),.CLK(clk_i),.Q(fracta_28_o[6:6]));
  DFFX1 desc35(.D(s_fractb_28_o[6:6]),.CLK(clk_i),.Q(fractb_28_o[6:6]));
  DFFX1 desc36(.D(s_fracta_28_o[7:7]),.CLK(clk_i),.Q(fracta_28_o[7:7]));
  DFFX1 desc37(.D(s_fractb_28_o[7:7]),.CLK(clk_i),.Q(fractb_28_o[7:7]));
  DFFX1 desc38(.D(s_fracta_28_o[8:8]),.CLK(clk_i),.Q(fracta_28_o[8:8]));
  DFFX1 desc39(.D(s_fractb_28_o[8:8]),.CLK(clk_i),.Q(fractb_28_o[8:8]));
  DFFX1 desc40(.D(s_fracta_28_o[9:9]),.CLK(clk_i),.Q(fracta_28_o[9:9]));
  DFFX1 desc41(.D(s_fractb_28_o[9:9]),.CLK(clk_i),.Q(fractb_28_o[9:9]));
  DFFX1 desc42(.D(s_fracta_28_o[10:10]),.CLK(clk_i),.Q(fracta_28_o[10:10]));
  DFFX1 desc43(.D(s_fractb_28_o[10:10]),.CLK(clk_i),.Q(fractb_28_o[10:10]));
  DFFX1 desc44(.D(s_fracta_28_o[11:11]),.CLK(clk_i),.Q(fracta_28_o[11:11]));
  DFFX1 desc45(.D(s_fractb_28_o[11:11]),.CLK(clk_i),.Q(fractb_28_o[11:11]));
  DFFX1 desc46(.D(s_fracta_28_o[12:12]),.CLK(clk_i),.Q(fracta_28_o[12:12]));
  DFFX1 desc47(.D(s_fractb_28_o[12:12]),.CLK(clk_i),.Q(fractb_28_o[12:12]));
  DFFX1 desc48(.D(s_fracta_28_o[13:13]),.CLK(clk_i),.Q(fracta_28_o[13:13]));
  DFFX1 desc49(.D(s_fractb_28_o[13:13]),.CLK(clk_i),.Q(fractb_28_o[13:13]));
  DFFX1 desc50(.D(s_fracta_28_o[14:14]),.CLK(clk_i),.Q(fracta_28_o[14:14]));
  DFFX1 desc51(.D(s_fractb_28_o[14:14]),.CLK(clk_i),.Q(fractb_28_o[14:14]));
  DFFX1 desc52(.D(s_fracta_28_o[15:15]),.CLK(clk_i),.Q(fracta_28_o[15:15]));
  DFFX1 desc53(.D(s_fractb_28_o[15:15]),.CLK(clk_i),.Q(fractb_28_o[15:15]));
  DFFX1 desc54(.D(s_fracta_28_o[16:16]),.CLK(clk_i),.Q(fracta_28_o[16:16]));
  DFFX1 desc55(.D(s_fractb_28_o[16:16]),.CLK(clk_i),.Q(fractb_28_o[16:16]));
  DFFX1 desc56(.D(s_fracta_28_o[17:17]),.CLK(clk_i),.Q(fracta_28_o[17:17]));
  DFFX1 desc57(.D(s_fractb_28_o[17:17]),.CLK(clk_i),.Q(fractb_28_o[17:17]));
  DFFX1 desc58(.D(s_fracta_28_o[18:18]),.CLK(clk_i),.Q(fracta_28_o[18:18]));
  DFFX1 desc59(.D(s_fractb_28_o[18:18]),.CLK(clk_i),.Q(fractb_28_o[18:18]));
  DFFX1 desc60(.D(s_fracta_28_o[19:19]),.CLK(clk_i),.Q(fracta_28_o[19:19]));
  DFFX1 desc61(.D(s_fractb_28_o[19:19]),.CLK(clk_i),.Q(fractb_28_o[19:19]));
  DFFX1 desc62(.D(s_fracta_28_o[20:20]),.CLK(clk_i),.Q(fracta_28_o[20:20]));
  DFFX1 desc63(.D(s_fractb_28_o[20:20]),.CLK(clk_i),.Q(fractb_28_o[20:20]));
  DFFX1 desc64(.D(s_fracta_28_o[21:21]),.CLK(clk_i),.Q(fracta_28_o[21:21]));
  DFFX1 desc65(.D(s_fractb_28_o[21:21]),.CLK(clk_i),.Q(fractb_28_o[21:21]));
  DFFX1 desc66(.D(s_fracta_28_o[22:22]),.CLK(clk_i),.Q(fracta_28_o[22:22]));
  DFFX1 desc67(.D(s_fractb_28_o[22:22]),.CLK(clk_i),.Q(fractb_28_o[22:22]));
  DFFX1 desc68(.D(s_fracta_28_o[23:23]),.CLK(clk_i),.Q(fracta_28_o[23:23]));
  DFFX1 desc69(.D(s_fractb_28_o[23:23]),.CLK(clk_i),.Q(fractb_28_o[23:23]));
  DFFX1 desc70(.D(s_fracta_28_o[24:24]),.CLK(clk_i),.Q(fracta_28_o[24:24]));
  DFFX1 desc71(.D(s_fractb_28_o[24:24]),.CLK(clk_i),.Q(fractb_28_o[24:24]));
  DFFX1 desc72(.D(s_fracta_28_o[25:25]),.CLK(clk_i),.Q(fracta_28_o[25:25]));
  DFFX1 desc73(.D(s_fractb_28_o[25:25]),.CLK(clk_i),.Q(fractb_28_o[25:25]));
  DFFX1 desc74(.D(s_fracta_28_o[26:26]),.CLK(clk_i),.Q(fracta_28_o[26:26]));
  DFFX1 desc75(.D(s_fractb_28_o[26:26]),.CLK(clk_i),.Q(fractb_28_o[26:26]));
  DFFX1 desc76(.D(s_fractb_28_o[0:0]),.CLK(clk_i),.Q(fractb_28_o[0:0]));
  DFFX1 desc77(.D(s_fracta_28_o[0:0]),.CLK(clk_i),.Q(fracta_28_o[0:0]));
  AOI222X1 U143(.IN1(N376),.IN2(n120),.IN3(N325),.IN4(n121),.IN5(N342),.IN6(n122),.QN(n119));
  AOI22X1 U144(.IN1(N393),.IN2(n123),.IN3(N410),.IN4(n124),.QN(n118));
  AOI222X1 U145(.IN1(n125),.IN2(n6),.IN3(n281),.IN4(n126),.IN5(n127),.IN6(N359),.QN(n117));
  OA221X1 U146(.IN1(n91),.IN2(n130),.IN3(n92),.IN4(n131),.IN5(n132),.Q(n129));
  OA22X1 U147(.IN1(n133),.IN2(n95),.IN3(n94),.IN4(n134),.Q(n132));
  OA222X1 U148(.IN1(n93),.IN2(n135),.IN3(n90),.IN4(n136),.IN5(n137),.IN6(n138),.Q(n128));
  AO222X1 U149(.IN1(n141),.IN2(N597),.IN3(n142),.IN4(N580),.IN5(n143),.IN6(N563),.Q(n140));
  AO221X1 U150(.IN1(N624),.IN2(n144),.IN3(n145),.IN4(N614),.IN5(n146),.Q(n139));
  AO22X1 U151(.IN1(n147),.IN2(N546),.IN3(N529),.IN4(n148),.Q(n146));
  AOI222X1 U154(.IN1(N375),.IN2(n120),.IN3(N324),.IN4(n121),.IN5(N341),.IN6(n122),.QN(n154));
  AOI222X1 U155(.IN1(n281),.IN2(n155),.IN3(n123),.IN4(N392),.IN5(n124),.IN6(N409),.QN(n153));
  OA221X1 U156(.IN1(n97),.IN2(n130),.IN3(n98),.IN4(n131),.IN5(n158),.Q(n157));
  OA22X1 U157(.IN1(n133),.IN2(n101),.IN3(n100),.IN4(n134),.Q(n158));
  OA222X1 U158(.IN1(n99),.IN2(n135),.IN3(n96),.IN4(n136),.IN5(n159),.IN6(n138),.Q(n156));
  AO222X1 U159(.IN1(n141),.IN2(N596),.IN3(n142),.IN4(N579),.IN5(n143),.IN6(N562),.Q(n161));
  AO221X1 U160(.IN1(N623),.IN2(n144),.IN3(n145),.IN4(N613),.IN5(n162),.Q(n160));
  AO22X1 U161(.IN1(n147),.IN2(N545),.IN3(N528),.IN4(n148),.Q(n162));
  AOI22X1 U163(.IN1(n11),.IN2(n149),.IN3(N307),.IN4(n150),.QN(n151));
  AOI222X1 U165(.IN1(N374),.IN2(n120),.IN3(N323),.IN4(n121),.IN5(N340),.IN6(n122),.QN(n167));
  AOI222X1 U166(.IN1(n281),.IN2(n168),.IN3(n123),.IN4(N391),.IN5(n124),.IN6(N408),.QN(n166));
  OA221X1 U167(.IN1(n103),.IN2(n130),.IN3(n104),.IN4(n131),.IN5(n171),.Q(n170));
  OA22X1 U168(.IN1(n133),.IN2(n107),.IN3(n106),.IN4(n134),.Q(n171));
  OA222X1 U169(.IN1(n105),.IN2(n135),.IN3(n102),.IN4(n136),.IN5(n172),.IN6(n138),.Q(n169));
  AO222X1 U170(.IN1(n141),.IN2(N595),.IN3(n142),.IN4(N578),.IN5(n143),.IN6(N561),.Q(n174));
  AO221X1 U171(.IN1(N622),.IN2(n144),.IN3(n145),.IN4(N612),.IN5(n175),.Q(n173));
  AO22X1 U172(.IN1(n147),.IN2(N544),.IN3(N527),.IN4(n148),.Q(n175));
  AOI222X1 U173(.IN1(N289),.IN2(n125),.IN3(N357),.IN4(n127),.IN5(n8),.IN6(n163),.QN(n165));
  AOI22X1 U174(.IN1(N272),.IN2(n149),.IN3(N306),.IN4(n150),.QN(n164));
  NAND4X0 U175(.IN1(n177),.IN2(n178),.IN3(n179),.IN4(n180),.QN(s_rzeros[2:2]));
  AOI221X1 U176(.IN1(N407),.IN2(n124),.IN3(N390),.IN4(n123),.IN5(n181),.QN(n180));
  AO222X1 U177(.IN1(N373),.IN2(n120),.IN3(N322),.IN4(n121),.IN5(N339),.IN6(n122),.Q(n181));
  AOI22X1 U178(.IN1(N305),.IN2(n150),.IN3(N231),.IN4(n182),.QN(n179));
  AO221X1 U179(.IN1(N288),.IN2(n125),.IN3(N254),.IN4(n163),.IN5(n183),.Q(n182));
  AO21X1 U180(.IN1(N271),.IN2(n149),.IN3(n278),.Q(n183));
  AO21X1 U181(.IN1(n187),.IN2(n188),.IN3(n176),.Q(n178));
  OA221X1 U182(.IN1(n267),.IN2(n130),.IN3(n268),.IN4(n131),.IN5(n189),.Q(n188));
  OA22X1 U183(.IN1(n133),.IN2(n271),.IN3(n270),.IN4(n134),.Q(n189));
  OA222X1 U184(.IN1(n269),.IN2(n135),.IN3(n266),.IN4(n136),.IN5(n190),.IN6(n138),.Q(n187));
  AO222X1 U185(.IN1(n141),.IN2(N594),.IN3(n142),.IN4(N577),.IN5(n143),.IN6(N560),.Q(n192));
  AO221X1 U186(.IN1(N621),.IN2(n144),.IN3(n145),.IN4(N611),.IN5(n193),.Q(n191));
  AO22X1 U187(.IN1(n147),.IN2(N543),.IN3(N526),.IN4(n148),.Q(n193));
  AO221X1 U189(.IN1(n279),.IN2(n195),.IN3(n163),.IN4(N253),.IN5(s_fract_sm_28[3:3]),.Q(n194));
  NAND4X0 U190(.IN1(n196),.IN2(n197),.IN3(n198),.IN4(n199),.QN(n195));
  AOI221X1 U191(.IN1(N389),.IN2(n123),.IN3(N372),.IN4(n120),.IN5(n200),.QN(n199));
  AO22X1 U192(.IN1(N321),.IN2(n121),.IN3(N338),.IN4(n122),.Q(n200));
  AOI22X1 U193(.IN1(N355),.IN2(n127),.IN3(n280),.IN4(N304),.QN(n198));
  AO21X1 U194(.IN1(n201),.IN2(n202),.IN3(n176),.Q(n196));
  OA221X1 U195(.IN1(n273),.IN2(n130),.IN3(n274),.IN4(n131),.IN5(n203),.Q(n202));
  OA22X1 U196(.IN1(n133),.IN2(n277),.IN3(n276),.IN4(n134),.Q(n203));
  OA222X1 U197(.IN1(n275),.IN2(n135),.IN3(n272),.IN4(n136),.IN5(n204),.IN6(n138),.Q(n201));
  AO222X1 U198(.IN1(n141),.IN2(N593),.IN3(n142),.IN4(N576),.IN5(n143),.IN6(N559),.Q(n206));
  AO221X1 U199(.IN1(N620),.IN2(n144),.IN3(n145),.IN4(N610),.IN5(n207),.Q(n205));
  AO22X1 U200(.IN1(n147),.IN2(N542),.IN3(N525),.IN4(n148),.Q(n207));
  AO221X1 U201(.IN1(n125),.IN2(N286),.IN3(n149),.IN4(N269),.IN5(n208),.Q(s_rzeros[0:0]));
  AO221X1 U202(.IN1(n279),.IN2(n209),.IN3(n163),.IN4(N252),.IN5(s_fract_sm_28[3:3]),.Q(n208));
  AND2X1 U203(.IN1(n184),.IN2(n210),.Q(n163));
  NAND4X0 U204(.IN1(n211),.IN2(n212),.IN3(n213),.IN4(n214),.QN(n209));
  AOI221X1 U205(.IN1(N388),.IN2(n123),.IN3(N371),.IN4(n120),.IN5(n215),.QN(n214));
  AO22X1 U206(.IN1(N320),.IN2(n121),.IN3(N337),.IN4(n122),.Q(n215));
  AND2X1 U207(.IN1(n186),.IN2(n216),.Q(n121));
  AND2X1 U208(.IN1(n282),.IN2(n218),.Q(n120));
  AOI22X1 U209(.IN1(N354),.IN2(n127),.IN3(n280),.IN4(N303),.QN(n213));
  AND2X1 U210(.IN1(n217),.IN2(n220),.Q(n127));
  AND2X1 U211(.IN1(n219),.IN2(n176),.Q(n124));
  AO21X1 U212(.IN1(n221),.IN2(n222),.IN3(n176),.Q(n211));
  OA221X1 U213(.IN1(N501),.IN2(n130),.IN3(N484),.IN4(n131),.IN5(n223),.Q(n222));
  OA22X1 U214(.IN1(n133),.IN2(N433),.IN3(N450),.IN4(n134),.Q(n223));
  OR2X1 U215(.IN1(n226),.IN2(n227),.Q(n130));
  OA222X1 U216(.IN1(N467),.IN2(n135),.IN3(N518),.IN4(n136),.IN5(n228),.IN6(n138),.Q(n221));
  AO222X1 U217(.IN1(n141),.IN2(N592),.IN3(n142),.IN4(N575),.IN5(n143),.IN6(N558),.Q(n230));
  AND2X1 U218(.IN1(n231),.IN2(n232),.Q(n143));
  AND2X1 U219(.IN1(n233),.IN2(n234),.Q(n141));
  AO221X1 U220(.IN1(N619),.IN2(n144),.IN3(n145),.IN4(N609),.IN5(n235),.Q(n229));
  AO22X1 U221(.IN1(n147),.IN2(N541),.IN3(N524),.IN4(n148),.Q(n235));
  OR2X1 U222(.IN1(n224),.IN2(n225),.Q(n135));
  AND2X1 U223(.IN1(n236),.IN2(n185),.Q(n125));
  AO22X1 U224(.IN1(s_fract_shr_28[9:9]),.IN2(n46),.IN3(opb_i[6:6]),.IN4(n32),.Q(s_fractb_28_o[9:9]));
  AO22X1 U225(.IN1(s_fract_shr_28[8:8]),.IN2(n46),.IN3(opb_i[5:5]),.IN4(n32),.Q(s_fractb_28_o[8:8]));
  AO22X1 U226(.IN1(s_fract_shr_28[7:7]),.IN2(n46),.IN3(opb_i[4:4]),.IN4(n32),.Q(s_fractb_28_o[7:7]));
  AO22X1 U227(.IN1(s_fract_shr_28[6:6]),.IN2(n46),.IN3(opb_i[3:3]),.IN4(n32),.Q(s_fractb_28_o[6:6]));
  AO22X1 U228(.IN1(s_fract_shr_28[5:5]),.IN2(n45),.IN3(opb_i[2:2]),.IN4(n32),.Q(s_fractb_28_o[5:5]));
  AO22X1 U229(.IN1(s_fract_shr_28[4:4]),.IN2(n45),.IN3(opb_i[1:1]),.IN4(n32),.Q(s_fractb_28_o[4:4]));
  AO22X1 U230(.IN1(s_fract_shr_28[3:3]),.IN2(n45),.IN3(opb_i[0:0]),.IN4(n32),.Q(s_fractb_28_o[3:3]));
  AO22X1 U231(.IN1(s_fract_shr_28[26:26]),.IN2(n45),.IN3(n237),.IN4(n32),.Q(s_fractb_28_o[26:26]));
  AO22X1 U232(.IN1(s_fract_shr_28[25:25]),.IN2(n45),.IN3(opb_i[22:22]),.IN4(n32),.Q(s_fractb_28_o[25:25]));
  AO22X1 U233(.IN1(s_fract_shr_28[24:24]),.IN2(n45),.IN3(opb_i[21:21]),.IN4(n32),.Q(s_fractb_28_o[24:24]));
  AO22X1 U234(.IN1(s_fract_shr_28[23:23]),.IN2(n45),.IN3(opb_i[20:20]),.IN4(n32),.Q(s_fractb_28_o[23:23]));
  AO22X1 U235(.IN1(s_fract_shr_28[22:22]),.IN2(n45),.IN3(opb_i[19:19]),.IN4(n31),.Q(s_fractb_28_o[22:22]));
  AO22X1 U236(.IN1(s_fract_shr_28[21:21]),.IN2(n45),.IN3(opb_i[18:18]),.IN4(n31),.Q(s_fractb_28_o[21:21]));
  AO22X1 U237(.IN1(s_fract_shr_28[20:20]),.IN2(n45),.IN3(opb_i[17:17]),.IN4(n31),.Q(s_fractb_28_o[20:20]));
  AO22X1 U238(.IN1(s_fract_shr_28[19:19]),.IN2(n44),.IN3(opb_i[16:16]),.IN4(n31),.Q(s_fractb_28_o[19:19]));
  AO22X1 U239(.IN1(s_fract_shr_28[18:18]),.IN2(n44),.IN3(opb_i[15:15]),.IN4(n31),.Q(s_fractb_28_o[18:18]));
  AO22X1 U240(.IN1(s_fract_shr_28[17:17]),.IN2(n44),.IN3(opb_i[14:14]),.IN4(n31),.Q(s_fractb_28_o[17:17]));
  AO22X1 U241(.IN1(s_fract_shr_28[16:16]),.IN2(n44),.IN3(opb_i[13:13]),.IN4(n31),.Q(s_fractb_28_o[16:16]));
  AO22X1 U242(.IN1(s_fract_shr_28[15:15]),.IN2(n44),.IN3(opb_i[12:12]),.IN4(n31),.Q(s_fractb_28_o[15:15]));
  AO22X1 U243(.IN1(s_fract_shr_28[14:14]),.IN2(n44),.IN3(opb_i[11:11]),.IN4(n31),.Q(s_fractb_28_o[14:14]));
  AO22X1 U244(.IN1(s_fract_shr_28[13:13]),.IN2(n44),.IN3(opb_i[10:10]),.IN4(n31),.Q(s_fractb_28_o[13:13]));
  AO22X1 U245(.IN1(s_fract_shr_28[12:12]),.IN2(n44),.IN3(opb_i[9:9]),.IN4(n31),.Q(s_fractb_28_o[12:12]));
  AO22X1 U246(.IN1(s_fract_shr_28[11:11]),.IN2(n44),.IN3(opb_i[8:8]),.IN4(n31),.Q(s_fractb_28_o[11:11]));
  AO22X1 U247(.IN1(s_fract_shr_28[10:10]),.IN2(n44),.IN3(opb_i[7:7]),.IN4(n31),.Q(s_fractb_28_o[10:10]));
  AO22X1 U248(.IN1(opa_i[6:6]),.IN2(n43),.IN3(s_fract_shr_28[9:9]),.IN4(n31),.Q(s_fracta_28_o[9:9]));
  AO22X1 U249(.IN1(opa_i[5:5]),.IN2(n43),.IN3(s_fract_shr_28[8:8]),.IN4(n31),.Q(s_fracta_28_o[8:8]));
  AO22X1 U250(.IN1(opa_i[4:4]),.IN2(n43),.IN3(s_fract_shr_28[7:7]),.IN4(n31),.Q(s_fracta_28_o[7:7]));
  AO22X1 U251(.IN1(opa_i[3:3]),.IN2(n43),.IN3(s_fract_shr_28[6:6]),.IN4(n31),.Q(s_fracta_28_o[6:6]));
  AO22X1 U252(.IN1(opa_i[2:2]),.IN2(n43),.IN3(s_fract_shr_28[5:5]),.IN4(n31),.Q(s_fracta_28_o[5:5]));
  AO22X1 U253(.IN1(opa_i[1:1]),.IN2(n43),.IN3(s_fract_shr_28[4:4]),.IN4(n31),.Q(s_fracta_28_o[4:4]));
  AO22X1 U254(.IN1(n34),.IN2(opa_i[0:0]),.IN3(s_fract_shr_28[3:3]),.IN4(n31),.Q(s_fracta_28_o[3:3]));
  AO22X1 U255(.IN1(s_fract_shr_28[26:26]),.IN2(n32),.IN3(n34),.IN4(n239),.Q(s_fracta_28_o[26:26]));
  AO22X1 U256(.IN1(opa_i[22:22]),.IN2(n43),.IN3(s_fract_shr_28[25:25]),.IN4(n31),.Q(s_fracta_28_o[25:25]));
  AO22X1 U257(.IN1(opa_i[21:21]),.IN2(n43),.IN3(s_fract_shr_28[24:24]),.IN4(n31),.Q(s_fracta_28_o[24:24]));
  AO22X1 U258(.IN1(opa_i[20:20]),.IN2(n43),.IN3(s_fract_shr_28[23:23]),.IN4(n31),.Q(s_fracta_28_o[23:23]));
  AO22X1 U259(.IN1(opa_i[19:19]),.IN2(n43),.IN3(s_fract_shr_28[22:22]),.IN4(n31),.Q(s_fracta_28_o[22:22]));
  AO22X1 U260(.IN1(opa_i[18:18]),.IN2(n38),.IN3(s_fract_shr_28[21:21]),.IN4(n31),.Q(s_fracta_28_o[21:21]));
  AO22X1 U261(.IN1(opa_i[17:17]),.IN2(n38),.IN3(s_fract_shr_28[20:20]),.IN4(n31),.Q(s_fracta_28_o[20:20]));
  AO22X1 U262(.IN1(opa_i[16:16]),.IN2(n38),.IN3(s_fract_shr_28[19:19]),.IN4(n31),.Q(s_fracta_28_o[19:19]));
  AO22X1 U263(.IN1(opa_i[15:15]),.IN2(n38),.IN3(s_fract_shr_28[18:18]),.IN4(n31),.Q(s_fracta_28_o[18:18]));
  AO22X1 U264(.IN1(opa_i[14:14]),.IN2(n38),.IN3(s_fract_shr_28[17:17]),.IN4(n31),.Q(s_fracta_28_o[17:17]));
  AO22X1 U265(.IN1(opa_i[13:13]),.IN2(n38),.IN3(s_fract_shr_28[16:16]),.IN4(n31),.Q(s_fracta_28_o[16:16]));
  AO22X1 U266(.IN1(opa_i[12:12]),.IN2(n38),.IN3(s_fract_shr_28[15:15]),.IN4(n31),.Q(s_fracta_28_o[15:15]));
  AO22X1 U267(.IN1(opa_i[11:11]),.IN2(n38),.IN3(s_fract_shr_28[14:14]),.IN4(n31),.Q(s_fracta_28_o[14:14]));
  AO22X1 U268(.IN1(opa_i[10:10]),.IN2(n38),.IN3(s_fract_shr_28[13:13]),.IN4(n31),.Q(s_fracta_28_o[13:13]));
  AO22X1 U269(.IN1(opa_i[9:9]),.IN2(n37),.IN3(s_fract_shr_28[12:12]),.IN4(n31),.Q(s_fracta_28_o[12:12]));
  AO22X1 U270(.IN1(opa_i[8:8]),.IN2(n37),.IN3(s_fract_shr_28[11:11]),.IN4(n31),.Q(s_fracta_28_o[11:11]));
  AO22X1 U271(.IN1(opa_i[7:7]),.IN2(n37),.IN3(s_fract_shr_28[10:10]),.IN4(n31),.Q(s_fracta_28_o[10:10]));
  OR2X1 U273(.IN1(n138),.IN2(s_fract_sm_28[21:21]),.Q(n148));
  AO22X1 U274(.IN1(N608),.IN2(n305),.IN3(N597),.IN4(s_fract_sm_28[26:26]),.Q(N614));
  AO22X1 U275(.IN1(N607),.IN2(n305),.IN3(N596),.IN4(s_fract_sm_28[26:26]),.Q(N613));
  AO22X1 U276(.IN1(N606),.IN2(n305),.IN3(N595),.IN4(s_fract_sm_28[26:26]),.Q(N612));
  AO22X1 U277(.IN1(N605),.IN2(n305),.IN3(N594),.IN4(s_fract_sm_28[26:26]),.Q(N611));
  AO22X1 U278(.IN1(N604),.IN2(n305),.IN3(N593),.IN4(s_fract_sm_28[26:26]),.Q(N610));
  AO22X1 U279(.IN1(N603),.IN2(n305),.IN3(N592),.IN4(s_fract_sm_28[26:26]),.Q(N609));
  AO22X1 U280(.IN1(n239),.IN2(n32),.IN3(n34),.IN4(n237),.Q(s_fract_sm_28[26:26]));
  AO22X1 U281(.IN1(N591),.IN2(n304),.IN3(N580),.IN4(s_fract_sm_28[25:25]),.Q(N597));
  AO22X1 U282(.IN1(N590),.IN2(n304),.IN3(N579),.IN4(s_fract_sm_28[25:25]),.Q(N596));
  AO22X1 U283(.IN1(N589),.IN2(n304),.IN3(N578),.IN4(s_fract_sm_28[25:25]),.Q(N595));
  AO22X1 U284(.IN1(N588),.IN2(n304),.IN3(N577),.IN4(s_fract_sm_28[25:25]),.Q(N594));
  AO22X1 U285(.IN1(N587),.IN2(n304),.IN3(N576),.IN4(s_fract_sm_28[25:25]),.Q(N593));
  AO22X1 U286(.IN1(N586),.IN2(n304),.IN3(N575),.IN4(s_fract_sm_28[25:25]),.Q(N592));
  AO22X1 U288(.IN1(N574),.IN2(n303),.IN3(N563),.IN4(s_fract_sm_28[24:24]),.Q(N580));
  AO22X1 U289(.IN1(N573),.IN2(n303),.IN3(N562),.IN4(s_fract_sm_28[24:24]),.Q(N579));
  AO22X1 U290(.IN1(N572),.IN2(n303),.IN3(N561),.IN4(s_fract_sm_28[24:24]),.Q(N578));
  AO22X1 U291(.IN1(N571),.IN2(n303),.IN3(N560),.IN4(s_fract_sm_28[24:24]),.Q(N577));
  AO22X1 U292(.IN1(N570),.IN2(n303),.IN3(N559),.IN4(s_fract_sm_28[24:24]),.Q(N576));
  AO22X1 U293(.IN1(N569),.IN2(n303),.IN3(N558),.IN4(s_fract_sm_28[24:24]),.Q(N575));
  AO22X1 U295(.IN1(N557),.IN2(n302),.IN3(N546),.IN4(s_fract_sm_28[23:23]),.Q(N563));
  AO22X1 U296(.IN1(N556),.IN2(n302),.IN3(N545),.IN4(s_fract_sm_28[23:23]),.Q(N562));
  AO22X1 U297(.IN1(N555),.IN2(n302),.IN3(N544),.IN4(s_fract_sm_28[23:23]),.Q(N561));
  AO22X1 U298(.IN1(N554),.IN2(n302),.IN3(N543),.IN4(s_fract_sm_28[23:23]),.Q(N560));
  AO22X1 U299(.IN1(N553),.IN2(n302),.IN3(N542),.IN4(s_fract_sm_28[23:23]),.Q(N559));
  AO22X1 U300(.IN1(N552),.IN2(n302),.IN3(N541),.IN4(s_fract_sm_28[23:23]),.Q(N558));
  AO22X1 U302(.IN1(N540),.IN2(n301),.IN3(N529),.IN4(s_fract_sm_28[22:22]),.Q(N546));
  AO22X1 U303(.IN1(N539),.IN2(n301),.IN3(N528),.IN4(s_fract_sm_28[22:22]),.Q(N545));
  AO22X1 U304(.IN1(N538),.IN2(n301),.IN3(N527),.IN4(s_fract_sm_28[22:22]),.Q(N544));
  AO22X1 U305(.IN1(N537),.IN2(n301),.IN3(N526),.IN4(s_fract_sm_28[22:22]),.Q(N543));
  AO22X1 U306(.IN1(N536),.IN2(n301),.IN3(N525),.IN4(s_fract_sm_28[22:22]),.Q(N542));
  AO22X1 U307(.IN1(N535),.IN2(n301),.IN3(N524),.IN4(s_fract_sm_28[22:22]),.Q(N541));
  AO22X1 U309(.IN1(N523),.IN2(n300),.IN3(s_fract_sm_28[21:21]),.IN4(N512),.Q(N529));
  AO22X1 U310(.IN1(N522),.IN2(n300),.IN3(N511),.IN4(s_fract_sm_28[21:21]),.Q(N528));
  AO22X1 U311(.IN1(N521),.IN2(n300),.IN3(N510),.IN4(s_fract_sm_28[21:21]),.Q(N527));
  AO22X1 U312(.IN1(N520),.IN2(n300),.IN3(N509),.IN4(s_fract_sm_28[21:21]),.Q(N526));
  AO22X1 U313(.IN1(N519),.IN2(n300),.IN3(N508),.IN4(s_fract_sm_28[21:21]),.Q(N525));
  AO22X1 U314(.IN1(N518),.IN2(n300),.IN3(N507),.IN4(s_fract_sm_28[21:21]),.Q(N524));
  AO22X1 U316(.IN1(N506),.IN2(n299),.IN3(N495),.IN4(s_fract_sm_28[20:20]),.Q(N512));
  AO22X1 U317(.IN1(N505),.IN2(n299),.IN3(N494),.IN4(s_fract_sm_28[20:20]),.Q(N511));
  AO22X1 U318(.IN1(N504),.IN2(n299),.IN3(N493),.IN4(s_fract_sm_28[20:20]),.Q(N510));
  AO22X1 U319(.IN1(N503),.IN2(n299),.IN3(N492),.IN4(s_fract_sm_28[20:20]),.Q(N509));
  AO22X1 U320(.IN1(N502),.IN2(n299),.IN3(N491),.IN4(s_fract_sm_28[20:20]),.Q(N508));
  AO22X1 U321(.IN1(N501),.IN2(n299),.IN3(N490),.IN4(s_fract_sm_28[20:20]),.Q(N507));
  AO22X1 U323(.IN1(N489),.IN2(n298),.IN3(N478),.IN4(s_fract_sm_28[19:19]),.Q(N495));
  AO22X1 U324(.IN1(N488),.IN2(n298),.IN3(N477),.IN4(s_fract_sm_28[19:19]),.Q(N494));
  AO22X1 U325(.IN1(N487),.IN2(n298),.IN3(N476),.IN4(s_fract_sm_28[19:19]),.Q(N493));
  AO22X1 U326(.IN1(N486),.IN2(n298),.IN3(N475),.IN4(s_fract_sm_28[19:19]),.Q(N492));
  AO22X1 U327(.IN1(N485),.IN2(n298),.IN3(N474),.IN4(s_fract_sm_28[19:19]),.Q(N491));
  AO22X1 U328(.IN1(N484),.IN2(n298),.IN3(N473),.IN4(s_fract_sm_28[19:19]),.Q(N490));
  AO22X1 U330(.IN1(N472),.IN2(n297),.IN3(N461),.IN4(s_fract_sm_28[18:18]),.Q(N478));
  AO22X1 U331(.IN1(N471),.IN2(n297),.IN3(N460),.IN4(s_fract_sm_28[18:18]),.Q(N477));
  AO22X1 U332(.IN1(N470),.IN2(n297),.IN3(N459),.IN4(s_fract_sm_28[18:18]),.Q(N476));
  AO22X1 U333(.IN1(N469),.IN2(n297),.IN3(N458),.IN4(s_fract_sm_28[18:18]),.Q(N475));
  AO22X1 U334(.IN1(N468),.IN2(n297),.IN3(N457),.IN4(s_fract_sm_28[18:18]),.Q(N474));
  AO22X1 U335(.IN1(N467),.IN2(n297),.IN3(N456),.IN4(s_fract_sm_28[18:18]),.Q(N473));
  AO22X1 U337(.IN1(N455),.IN2(n296),.IN3(N444),.IN4(s_fract_sm_28[17:17]),.Q(N461));
  AO22X1 U338(.IN1(N454),.IN2(n296),.IN3(N443),.IN4(s_fract_sm_28[17:17]),.Q(N460));
  AO22X1 U339(.IN1(N453),.IN2(n296),.IN3(N442),.IN4(s_fract_sm_28[17:17]),.Q(N459));
  AO22X1 U340(.IN1(N452),.IN2(n296),.IN3(N441),.IN4(s_fract_sm_28[17:17]),.Q(N458));
  AO22X1 U341(.IN1(N451),.IN2(n296),.IN3(N440),.IN4(s_fract_sm_28[17:17]),.Q(N457));
  AO22X1 U342(.IN1(N450),.IN2(n296),.IN3(N439),.IN4(s_fract_sm_28[17:17]),.Q(N456));
  AO22X1 U344(.IN1(N438),.IN2(n295),.IN3(N427),.IN4(s_fract_sm_28[16:16]),.Q(N444));
  AO22X1 U345(.IN1(N437),.IN2(n295),.IN3(N426),.IN4(s_fract_sm_28[16:16]),.Q(N443));
  AO22X1 U346(.IN1(N436),.IN2(n295),.IN3(N425),.IN4(s_fract_sm_28[16:16]),.Q(N442));
  AO22X1 U347(.IN1(N435),.IN2(n295),.IN3(N424),.IN4(s_fract_sm_28[16:16]),.Q(N441));
  AO22X1 U348(.IN1(N434),.IN2(n295),.IN3(N423),.IN4(s_fract_sm_28[16:16]),.Q(N440));
  AO22X1 U349(.IN1(N433),.IN2(n295),.IN3(N422),.IN4(s_fract_sm_28[16:16]),.Q(N439));
  AO22X1 U350(.IN1(opb_i[13:13]),.IN2(n37),.IN3(opa_i[13:13]),.IN4(n18),.Q(s_fract_sm_28[16:16]));
  AO22X1 U351(.IN1(N421),.IN2(n294),.IN3(s_fract_sm_28[15:15]),.IN4(N410),.Q(N427));
  AO22X1 U352(.IN1(N420),.IN2(n294),.IN3(N409),.IN4(s_fract_sm_28[15:15]),.Q(N426));
  AO22X1 U353(.IN1(N419),.IN2(n294),.IN3(N408),.IN4(s_fract_sm_28[15:15]),.Q(N425));
  AO22X1 U354(.IN1(N418),.IN2(n294),.IN3(N407),.IN4(s_fract_sm_28[15:15]),.Q(N424));
  AO22X1 U355(.IN1(N417),.IN2(n294),.IN3(N406),.IN4(s_fract_sm_28[15:15]),.Q(N423));
  AO22X1 U356(.IN1(N416),.IN2(n294),.IN3(N405),.IN4(s_fract_sm_28[15:15]),.Q(N422));
  AO22X1 U357(.IN1(opb_i[12:12]),.IN2(n36),.IN3(opa_i[12:12]),.IN4(n18),.Q(s_fract_sm_28[15:15]));
  AO22X1 U358(.IN1(N404),.IN2(n293),.IN3(N393),.IN4(s_fract_sm_28[14:14]),.Q(N410));
  AO22X1 U359(.IN1(N403),.IN2(n293),.IN3(N392),.IN4(s_fract_sm_28[14:14]),.Q(N409));
  AO22X1 U360(.IN1(N402),.IN2(n293),.IN3(N391),.IN4(s_fract_sm_28[14:14]),.Q(N408));
  AO22X1 U361(.IN1(N401),.IN2(n293),.IN3(N390),.IN4(s_fract_sm_28[14:14]),.Q(N407));
  AO22X1 U362(.IN1(N400),.IN2(n293),.IN3(N389),.IN4(s_fract_sm_28[14:14]),.Q(N406));
  AO22X1 U363(.IN1(N399),.IN2(n293),.IN3(N388),.IN4(s_fract_sm_28[14:14]),.Q(N405));
  AO22X1 U364(.IN1(opb_i[11:11]),.IN2(n36),.IN3(opa_i[11:11]),.IN4(n19),.Q(s_fract_sm_28[14:14]));
  AO22X1 U365(.IN1(N387),.IN2(n292),.IN3(N376),.IN4(s_fract_sm_28[13:13]),.Q(N393));
  AO22X1 U366(.IN1(N386),.IN2(n292),.IN3(N375),.IN4(s_fract_sm_28[13:13]),.Q(N392));
  AO22X1 U367(.IN1(N385),.IN2(n292),.IN3(N374),.IN4(s_fract_sm_28[13:13]),.Q(N391));
  AO22X1 U368(.IN1(N384),.IN2(n292),.IN3(N373),.IN4(s_fract_sm_28[13:13]),.Q(N390));
  AO22X1 U369(.IN1(N383),.IN2(n292),.IN3(N372),.IN4(s_fract_sm_28[13:13]),.Q(N389));
  AO22X1 U370(.IN1(N382),.IN2(n292),.IN3(N371),.IN4(s_fract_sm_28[13:13]),.Q(N388));
  AO22X1 U371(.IN1(opb_i[10:10]),.IN2(n36),.IN3(opa_i[10:10]),.IN4(n19),.Q(s_fract_sm_28[13:13]));
  AO22X1 U372(.IN1(N370),.IN2(n291),.IN3(N359),.IN4(s_fract_sm_28[12:12]),.Q(N376));
  AO22X1 U373(.IN1(N369),.IN2(n291),.IN3(N358),.IN4(s_fract_sm_28[12:12]),.Q(N375));
  AO22X1 U374(.IN1(N368),.IN2(n291),.IN3(N357),.IN4(s_fract_sm_28[12:12]),.Q(N374));
  AO22X1 U375(.IN1(N367),.IN2(n291),.IN3(N356),.IN4(s_fract_sm_28[12:12]),.Q(N373));
  AO22X1 U376(.IN1(N366),.IN2(n291),.IN3(N355),.IN4(s_fract_sm_28[12:12]),.Q(N372));
  AO22X1 U377(.IN1(N365),.IN2(n291),.IN3(N354),.IN4(s_fract_sm_28[12:12]),.Q(N371));
  AO22X1 U378(.IN1(opb_i[9:9]),.IN2(n36),.IN3(opa_i[9:9]),.IN4(n19),.Q(s_fract_sm_28[12:12]));
  AO22X1 U379(.IN1(N353),.IN2(n290),.IN3(N342),.IN4(s_fract_sm_28[11:11]),.Q(N359));
  AO22X1 U380(.IN1(N352),.IN2(n290),.IN3(N341),.IN4(s_fract_sm_28[11:11]),.Q(N358));
  AO22X1 U381(.IN1(N351),.IN2(n290),.IN3(N340),.IN4(s_fract_sm_28[11:11]),.Q(N357));
  AO22X1 U382(.IN1(N350),.IN2(n290),.IN3(N339),.IN4(s_fract_sm_28[11:11]),.Q(N356));
  AO22X1 U383(.IN1(N349),.IN2(n290),.IN3(N338),.IN4(s_fract_sm_28[11:11]),.Q(N355));
  AO22X1 U384(.IN1(N348),.IN2(n290),.IN3(N337),.IN4(s_fract_sm_28[11:11]),.Q(N354));
  AO22X1 U385(.IN1(opb_i[8:8]),.IN2(n36),.IN3(opa_i[8:8]),.IN4(n19),.Q(s_fract_sm_28[11:11]));
  AO22X1 U386(.IN1(N336),.IN2(n289),.IN3(N325),.IN4(s_fract_sm_28[10:10]),.Q(N342));
  AO22X1 U387(.IN1(N335),.IN2(n289),.IN3(N324),.IN4(s_fract_sm_28[10:10]),.Q(N341));
  AO22X1 U388(.IN1(N334),.IN2(n289),.IN3(N323),.IN4(s_fract_sm_28[10:10]),.Q(N340));
  AO22X1 U389(.IN1(N333),.IN2(n289),.IN3(N322),.IN4(s_fract_sm_28[10:10]),.Q(N339));
  AO22X1 U390(.IN1(N332),.IN2(n289),.IN3(N321),.IN4(s_fract_sm_28[10:10]),.Q(N338));
  AO22X1 U391(.IN1(N331),.IN2(n289),.IN3(N320),.IN4(s_fract_sm_28[10:10]),.Q(N337));
  AO22X1 U392(.IN1(opb_i[7:7]),.IN2(n36),.IN3(opa_i[7:7]),.IN4(n19),.Q(s_fract_sm_28[10:10]));
  AO22X1 U393(.IN1(N319),.IN2(n288),.IN3(s_fract_sm_28[9:9]),.IN4(N308),.Q(N325));
  AO22X1 U394(.IN1(N318),.IN2(n288),.IN3(N307),.IN4(s_fract_sm_28[9:9]),.Q(N324));
  AO22X1 U395(.IN1(N317),.IN2(n288),.IN3(N306),.IN4(s_fract_sm_28[9:9]),.Q(N323));
  AO22X1 U396(.IN1(N316),.IN2(n288),.IN3(N305),.IN4(s_fract_sm_28[9:9]),.Q(N322));
  AO22X1 U397(.IN1(N315),.IN2(n288),.IN3(N304),.IN4(s_fract_sm_28[9:9]),.Q(N321));
  AO22X1 U398(.IN1(N314),.IN2(n288),.IN3(N303),.IN4(s_fract_sm_28[9:9]),.Q(N320));
  AO22X1 U399(.IN1(opb_i[6:6]),.IN2(n35),.IN3(opa_i[6:6]),.IN4(n19),.Q(s_fract_sm_28[9:9]));
  AO22X1 U400(.IN1(N302),.IN2(n287),.IN3(n6),.IN4(s_fract_sm_28[8:8]),.Q(N308));
  AO22X1 U401(.IN1(N301),.IN2(n287),.IN3(N290),.IN4(s_fract_sm_28[8:8]),.Q(N307));
  AO22X1 U402(.IN1(N300),.IN2(n287),.IN3(N289),.IN4(s_fract_sm_28[8:8]),.Q(N306));
  AO22X1 U403(.IN1(N299),.IN2(n287),.IN3(N288),.IN4(s_fract_sm_28[8:8]),.Q(N305));
  AO22X1 U404(.IN1(N298),.IN2(n287),.IN3(N287),.IN4(s_fract_sm_28[8:8]),.Q(N304));
  AO22X1 U405(.IN1(N297),.IN2(n287),.IN3(N286),.IN4(s_fract_sm_28[8:8]),.Q(N303));
  AO22X1 U408(.IN1(N284),.IN2(n286),.IN3(n11),.IN4(s_fract_sm_28[7:7]),.Q(N290));
  AO22X1 U409(.IN1(N283),.IN2(n286),.IN3(N272),.IN4(s_fract_sm_28[7:7]),.Q(N289));
  AO22X1 U410(.IN1(N282),.IN2(n286),.IN3(N271),.IN4(s_fract_sm_28[7:7]),.Q(N288));
  AO22X1 U411(.IN1(N281),.IN2(n286),.IN3(N270),.IN4(s_fract_sm_28[7:7]),.Q(N287));
  AO22X1 U412(.IN1(N280),.IN2(n286),.IN3(N269),.IN4(s_fract_sm_28[7:7]),.Q(N286));
  AO22X1 U413(.IN1(opb_i[4:4]),.IN2(n35),.IN3(opa_i[4:4]),.IN4(n19),.Q(s_fract_sm_28[7:7]));
  AO22X1 U416(.IN1(N266),.IN2(n285),.IN3(n8),.IN4(s_fract_sm_28[6:6]),.Q(N272));
  AO22X1 U417(.IN1(N265),.IN2(n285),.IN3(N254),.IN4(s_fract_sm_28[6:6]),.Q(N271));
  AO22X1 U418(.IN1(N264),.IN2(n285),.IN3(N253),.IN4(s_fract_sm_28[6:6]),.Q(N270));
  AO22X1 U419(.IN1(N263),.IN2(n285),.IN3(N252),.IN4(s_fract_sm_28[6:6]),.Q(N269));
  AO22X1 U420(.IN1(opb_i[3:3]),.IN2(n35),.IN3(opa_i[3:3]),.IN4(n19),.Q(s_fract_sm_28[6:6]));
  AO22X1 U424(.IN1(N248),.IN2(n284),.IN3(N238),.IN4(s_fract_sm_28[5:5]),.Q(N254));
  AO22X1 U425(.IN1(N247),.IN2(n284),.IN3(n16),.IN4(s_fract_sm_28[5:5]),.Q(N253));
  AO22X1 U426(.IN1(N246),.IN2(n284),.IN3(N236),.IN4(s_fract_sm_28[5:5]),.Q(N252));
  AO22X1 U427(.IN1(opb_i[2:2]),.IN2(n35),.IN3(opa_i[2:2]),.IN4(n19),.Q(s_fract_sm_28[5:5]));
  AO22X1 U432(.IN1(N231),.IN2(n283),.IN3(s_fract_sm_28[4:4]),.IN4(s_fract_sm_28[3:3]),.Q(N236));
  AO22X1 U433(.IN1(opb_i[1:1]),.IN2(n35),.IN3(opa_i[1:1]),.IN4(n19),.Q(s_fract_sm_28[4:4]));
  AO221X1 U436(.IN1(N186),.IN2(n240),.IN3(N170),.IN4(n241),.IN5(n242),.Q(N194));
  AO22X1 U437(.IN1(N146),.IN2(n243),.IN3(N162),.IN4(n244),.Q(n242));
  AO221X1 U438(.IN1(N185),.IN2(n240),.IN3(N169),.IN4(n241),.IN5(n245),.Q(N193));
  AO22X1 U439(.IN1(N145),.IN2(n243),.IN3(N161),.IN4(n244),.Q(n245));
  AO221X1 U440(.IN1(N184),.IN2(n240),.IN3(N168),.IN4(n241),.IN5(n246),.Q(N192));
  AO22X1 U441(.IN1(N144),.IN2(n243),.IN3(N160),.IN4(n244),.Q(n246));
  AO221X1 U442(.IN1(N183),.IN2(n240),.IN3(N167),.IN4(n241),.IN5(n247),.Q(N191));
  AO22X1 U443(.IN1(N143),.IN2(n243),.IN3(N159),.IN4(n244),.Q(n247));
  AO221X1 U444(.IN1(N182),.IN2(n240),.IN3(N166),.IN4(n241),.IN5(n248),.Q(N190));
  AO22X1 U445(.IN1(N142),.IN2(n243),.IN3(N158),.IN4(n244),.Q(n248));
  AO221X1 U446(.IN1(N181),.IN2(n240),.IN3(N165),.IN4(n241),.IN5(n249),.Q(N189));
  AO22X1 U447(.IN1(N141),.IN2(n243),.IN3(N157),.IN4(n244),.Q(n249));
  AO221X1 U448(.IN1(N180),.IN2(n240),.IN3(N164),.IN4(n241),.IN5(n250),.Q(N188));
  AO22X1 U449(.IN1(N140),.IN2(n243),.IN3(N156),.IN4(n244),.Q(n250));
  AO221X1 U450(.IN1(N179),.IN2(n240),.IN3(N163),.IN4(n241),.IN5(n251),.Q(N187));
  AO22X1 U451(.IN1(N139),.IN2(n243),.IN3(N155),.IN4(n244),.Q(n251));
  XOR2X1 U452(.IN1(n237),.IN2(n239),.Q(n252));
  NAND4X0 U453(.IN1(n48),.IN2(n307),.IN3(n253),.IN4(n254),.QN(n239));
  NOR4X0 U454(.IN1(opa_i[30:30]),.IN2(n49),.IN3(opa_i[28:28]),.IN4(opa_i[27:27]),.QN(n254));
  NAND4X0 U455(.IN1(n308),.IN2(n68),.IN3(n255),.IN4(n256),.QN(n237));
  NOR4X0 U456(.IN1(opb_i[30:30]),.IN2(opb_i[29:29]),.IN3(opb_i[28:28]),.IN4(opb_i[27:27]),.QN(n256));
  AO22X1 U457(.IN1(opa_i[30:30]),.IN2(n35),.IN3(opb_i[30:30]),.IN4(n19),.Q(N131));
  AO22X1 U458(.IN1(n49),.IN2(n35),.IN3(opb_i[29:29]),.IN4(n19),.Q(N130));
  AO22X1 U459(.IN1(opa_i[28:28]),.IN2(n35),.IN3(opb_i[28:28]),.IN4(n19),.Q(N129));
  AO22X1 U460(.IN1(opa_i[27:27]),.IN2(n35),.IN3(opb_i[27:27]),.IN4(n19),.Q(N128));
  AO22X1 U461(.IN1(opa_i[26:26]),.IN2(n34),.IN3(opb_i[26:26]),.IN4(n19),.Q(N127));
  AO22X1 U462(.IN1(opa_i[25:25]),.IN2(n34),.IN3(opb_i[25:25]),.IN4(n19),.Q(N126));
  AO22X1 U463(.IN1(opa_i[24:24]),.IN2(n34),.IN3(opb_i[24:24]),.IN4(n19),.Q(N125));
  AO22X1 U464(.IN1(n47),.IN2(n38),.IN3(opb_i[23:23]),.IN4(n31),.Q(N124));
  pre_norm_addsub_DW01_sub_0_inj sub_1_root_sub_148(.A({opa_i[30:30],n49,opa_i[28:24],n47}),.B(opb_i[30:23]),.CI(1'b1),.DIFF({N186,N185,N184,N183,N182,N181,N180,N179}));
  pre_norm_addsub_DW01_sub_1_inj sub_147(.A({opa_i[30:30],n49,opa_i[28:24],n47}),.B(opb_i[30:23]),.CI(1'b0),.DIFF({N170,N169,N168,N167,N166,N165,N164,N163}));
  pre_norm_addsub_DW01_sub_2_inj sub_1_root_sub_146(.A(opb_i[30:23]),.B({opa_i[30:30],n49,opa_i[28:24],n47}),.CI(1'b1),.DIFF({N162,N161,N160,N159,N158,N157,N156,N155}));
  pre_norm_addsub_DW01_sub_3_inj sub_145(.A(opb_i[30:23]),.B({opa_i[30:30],n49,opa_i[28:24],n47}),.CI(1'b0),.DIFF({N146,N145,N144,N143,N142,N141,N140,N139}));
  HADDX1 desc78(.A0(N610),.B0(N609),.C1(\add_105_I28_L14036_C161/carry[2] ),.SO(N620));
  HADDX1 desc79(.A0(N611),.B0(\add_105_I28_L14036_C161/carry[2] ),.C1(\add_105_I28_L14036_C161/carry[3] ),.SO(N621));
  HADDX1 desc80(.A0(N612),.B0(\add_105_I28_L14036_C161/carry[3] ),.C1(\add_105_I28_L14036_C161/carry[4] ),.SO(N622));
  HADDX1 desc81(.A0(N613),.B0(\add_105_I28_L14036_C161/carry[4] ),.C1(\add_105_I28_L14036_C161/carry[5] ),.SO(N623));
  HADDX1 desc82(.A0(N593),.B0(N592),.C1(\add_105_I27_L14036_C161/carry[2] ),.SO(N604));
  HADDX1 desc83(.A0(N594),.B0(\add_105_I27_L14036_C161/carry[2] ),.C1(\add_105_I27_L14036_C161/carry[3] ),.SO(N605));
  HADDX1 desc84(.A0(N595),.B0(\add_105_I27_L14036_C161/carry[3] ),.C1(\add_105_I27_L14036_C161/carry[4] ),.SO(N606));
  HADDX1 desc85(.A0(N596),.B0(\add_105_I27_L14036_C161/carry[4] ),.C1(\add_105_I27_L14036_C161/carry[5] ),.SO(N607));
  HADDX1 desc86(.A0(N576),.B0(N575),.C1(\add_105_I26_L14036_C161/carry[2] ),.SO(N587));
  HADDX1 desc87(.A0(N577),.B0(\add_105_I26_L14036_C161/carry[2] ),.C1(\add_105_I26_L14036_C161/carry[3] ),.SO(N588));
  HADDX1 desc88(.A0(N578),.B0(\add_105_I26_L14036_C161/carry[3] ),.C1(\add_105_I26_L14036_C161/carry[4] ),.SO(N589));
  HADDX1 desc89(.A0(N579),.B0(\add_105_I26_L14036_C161/carry[4] ),.C1(\add_105_I26_L14036_C161/carry[5] ),.SO(N590));
  HADDX1 desc90(.A0(N559),.B0(N558),.C1(\add_105_I25_L14036_C161/carry[2] ),.SO(N570));
  HADDX1 desc91(.A0(N560),.B0(\add_105_I25_L14036_C161/carry[2] ),.C1(\add_105_I25_L14036_C161/carry[3] ),.SO(N571));
  HADDX1 desc92(.A0(N561),.B0(\add_105_I25_L14036_C161/carry[3] ),.C1(\add_105_I25_L14036_C161/carry[4] ),.SO(N572));
  HADDX1 desc93(.A0(N562),.B0(\add_105_I25_L14036_C161/carry[4] ),.C1(\add_105_I25_L14036_C161/carry[5] ),.SO(N573));
  HADDX1 desc94(.A0(N542),.B0(N541),.C1(\add_105_I24_L14036_C161/carry[2] ),.SO(N553));
  HADDX1 desc95(.A0(N543),.B0(\add_105_I24_L14036_C161/carry[2] ),.C1(\add_105_I24_L14036_C161/carry[3] ),.SO(N554));
  HADDX1 desc96(.A0(N544),.B0(\add_105_I24_L14036_C161/carry[3] ),.C1(\add_105_I24_L14036_C161/carry[4] ),.SO(N555));
  HADDX1 desc97(.A0(N545),.B0(\add_105_I24_L14036_C161/carry[4] ),.C1(\add_105_I24_L14036_C161/carry[5] ),.SO(N556));
  HADDX1 desc98(.A0(N525),.B0(N524),.C1(\add_105_I23_L14036_C161/carry[2] ),.SO(N536));
  HADDX1 desc99(.A0(N526),.B0(\add_105_I23_L14036_C161/carry[2] ),.C1(\add_105_I23_L14036_C161/carry[3] ),.SO(N537));
  HADDX1 desc100(.A0(N527),.B0(\add_105_I23_L14036_C161/carry[3] ),.C1(\add_105_I23_L14036_C161/carry[4] ),.SO(N538));
  HADDX1 desc101(.A0(N528),.B0(\add_105_I23_L14036_C161/carry[4] ),.C1(\add_105_I23_L14036_C161/carry[5] ),.SO(N539));
  HADDX1 desc102(.A0(N508),.B0(N507),.C1(\add_105_I22_L14036_C161/carry[2] ),.SO(N519));
  HADDX1 desc103(.A0(N509),.B0(\add_105_I22_L14036_C161/carry[2] ),.C1(\add_105_I22_L14036_C161/carry[3] ),.SO(N520));
  HADDX1 desc104(.A0(N510),.B0(\add_105_I22_L14036_C161/carry[3] ),.C1(\add_105_I22_L14036_C161/carry[4] ),.SO(N521));
  HADDX1 desc105(.A0(N511),.B0(\add_105_I22_L14036_C161/carry[4] ),.C1(\add_105_I22_L14036_C161/carry[5] ),.SO(N522));
  HADDX1 desc106(.A0(N491),.B0(N490),.C1(\add_105_I21_L14036_C161/carry[2] ),.SO(N502));
  HADDX1 desc107(.A0(N492),.B0(\add_105_I21_L14036_C161/carry[2] ),.C1(\add_105_I21_L14036_C161/carry[3] ),.SO(N503));
  HADDX1 desc108(.A0(N493),.B0(\add_105_I21_L14036_C161/carry[3] ),.C1(\add_105_I21_L14036_C161/carry[4] ),.SO(N504));
  HADDX1 desc109(.A0(N494),.B0(\add_105_I21_L14036_C161/carry[4] ),.C1(\add_105_I21_L14036_C161/carry[5] ),.SO(N505));
  HADDX1 desc110(.A0(N474),.B0(N473),.C1(\add_105_I20_L14036_C161/carry[2] ),.SO(N485));
  HADDX1 desc111(.A0(N475),.B0(\add_105_I20_L14036_C161/carry[2] ),.C1(\add_105_I20_L14036_C161/carry[3] ),.SO(N486));
  HADDX1 desc112(.A0(N476),.B0(\add_105_I20_L14036_C161/carry[3] ),.C1(\add_105_I20_L14036_C161/carry[4] ),.SO(N487));
  HADDX1 desc113(.A0(N477),.B0(\add_105_I20_L14036_C161/carry[4] ),.C1(\add_105_I20_L14036_C161/carry[5] ),.SO(N488));
  HADDX1 desc114(.A0(N457),.B0(N456),.C1(\add_105_I19_L14036_C161/carry[2] ),.SO(N468));
  HADDX1 desc115(.A0(N458),.B0(\add_105_I19_L14036_C161/carry[2] ),.C1(\add_105_I19_L14036_C161/carry[3] ),.SO(N469));
  HADDX1 desc116(.A0(N459),.B0(\add_105_I19_L14036_C161/carry[3] ),.C1(\add_105_I19_L14036_C161/carry[4] ),.SO(N470));
  HADDX1 desc117(.A0(N460),.B0(\add_105_I19_L14036_C161/carry[4] ),.C1(\add_105_I19_L14036_C161/carry[5] ),.SO(N471));
  HADDX1 desc118(.A0(N440),.B0(N439),.C1(\add_105_I18_L14036_C161/carry[2] ),.SO(N451));
  HADDX1 desc119(.A0(N441),.B0(\add_105_I18_L14036_C161/carry[2] ),.C1(\add_105_I18_L14036_C161/carry[3] ),.SO(N452));
  HADDX1 desc120(.A0(N442),.B0(\add_105_I18_L14036_C161/carry[3] ),.C1(\add_105_I18_L14036_C161/carry[4] ),.SO(N453));
  HADDX1 desc121(.A0(N443),.B0(\add_105_I18_L14036_C161/carry[4] ),.C1(\add_105_I18_L14036_C161/carry[5] ),.SO(N454));
  HADDX1 desc122(.A0(N423),.B0(N422),.C1(\add_105_I17_L14036_C161/carry[2] ),.SO(N434));
  HADDX1 desc123(.A0(N424),.B0(\add_105_I17_L14036_C161/carry[2] ),.C1(\add_105_I17_L14036_C161/carry[3] ),.SO(N435));
  HADDX1 desc124(.A0(N425),.B0(\add_105_I17_L14036_C161/carry[3] ),.C1(\add_105_I17_L14036_C161/carry[4] ),.SO(N436));
  HADDX1 desc125(.A0(N426),.B0(\add_105_I17_L14036_C161/carry[4] ),.C1(\add_105_I17_L14036_C161/carry[5] ),.SO(N437));
  HADDX1 desc126(.A0(N406),.B0(N405),.C1(\add_105_I16_L14036_C161/carry[2] ),.SO(N417));
  HADDX1 desc127(.A0(N407),.B0(\add_105_I16_L14036_C161/carry[2] ),.C1(\add_105_I16_L14036_C161/carry[3] ),.SO(N418));
  HADDX1 desc128(.A0(N408),.B0(\add_105_I16_L14036_C161/carry[3] ),.C1(\add_105_I16_L14036_C161/carry[4] ),.SO(N419));
  HADDX1 desc129(.A0(N409),.B0(\add_105_I16_L14036_C161/carry[4] ),.C1(\add_105_I16_L14036_C161/carry[5] ),.SO(N420));
  HADDX1 desc130(.A0(N389),.B0(N388),.C1(\add_105_I15_L14036_C161/carry[2] ),.SO(N400));
  HADDX1 desc131(.A0(N390),.B0(\add_105_I15_L14036_C161/carry[2] ),.C1(\add_105_I15_L14036_C161/carry[3] ),.SO(N401));
  HADDX1 desc132(.A0(N391),.B0(\add_105_I15_L14036_C161/carry[3] ),.C1(\add_105_I15_L14036_C161/carry[4] ),.SO(N402));
  HADDX1 desc133(.A0(N392),.B0(\add_105_I15_L14036_C161/carry[4] ),.C1(\add_105_I15_L14036_C161/carry[5] ),.SO(N403));
  HADDX1 desc134(.A0(N372),.B0(N371),.C1(\add_105_I14_L14036_C161/carry[2] ),.SO(N383));
  HADDX1 desc135(.A0(N373),.B0(\add_105_I14_L14036_C161/carry[2] ),.C1(\add_105_I14_L14036_C161/carry[3] ),.SO(N384));
  HADDX1 desc136(.A0(N374),.B0(\add_105_I14_L14036_C161/carry[3] ),.C1(\add_105_I14_L14036_C161/carry[4] ),.SO(N385));
  HADDX1 desc137(.A0(N375),.B0(\add_105_I14_L14036_C161/carry[4] ),.C1(\add_105_I14_L14036_C161/carry[5] ),.SO(N386));
  HADDX1 desc138(.A0(N355),.B0(N354),.C1(\add_105_I13_L14036_C161/carry[2] ),.SO(N366));
  HADDX1 desc139(.A0(N356),.B0(\add_105_I13_L14036_C161/carry[2] ),.C1(\add_105_I13_L14036_C161/carry[3] ),.SO(N367));
  HADDX1 desc140(.A0(N357),.B0(\add_105_I13_L14036_C161/carry[3] ),.C1(\add_105_I13_L14036_C161/carry[4] ),.SO(N368));
  HADDX1 desc141(.A0(N358),.B0(\add_105_I13_L14036_C161/carry[4] ),.C1(\add_105_I13_L14036_C161/carry[5] ),.SO(N369));
  HADDX1 desc142(.A0(N338),.B0(N337),.C1(\add_105_I12_L14036_C161/carry[2] ),.SO(N349));
  HADDX1 desc143(.A0(N339),.B0(\add_105_I12_L14036_C161/carry[2] ),.C1(\add_105_I12_L14036_C161/carry[3] ),.SO(N350));
  HADDX1 desc144(.A0(N340),.B0(\add_105_I12_L14036_C161/carry[3] ),.C1(\add_105_I12_L14036_C161/carry[4] ),.SO(N351));
  HADDX1 desc145(.A0(N341),.B0(\add_105_I12_L14036_C161/carry[4] ),.C1(\add_105_I12_L14036_C161/carry[5] ),.SO(N352));
  HADDX1 desc146(.A0(N321),.B0(N320),.C1(\add_105_I11_L14036_C161/carry[2] ),.SO(N332));
  HADDX1 desc147(.A0(N322),.B0(\add_105_I11_L14036_C161/carry[2] ),.C1(\add_105_I11_L14036_C161/carry[3] ),.SO(N333));
  HADDX1 desc148(.A0(N323),.B0(\add_105_I11_L14036_C161/carry[3] ),.C1(\add_105_I11_L14036_C161/carry[4] ),.SO(N334));
  HADDX1 desc149(.A0(N324),.B0(\add_105_I11_L14036_C161/carry[4] ),.C1(\add_105_I11_L14036_C161/carry[5] ),.SO(N335));
  HADDX1 desc150(.A0(N304),.B0(N303),.C1(\add_105_I10_L14036_C161/carry[2] ),.SO(N315));
  HADDX1 desc151(.A0(N305),.B0(\add_105_I10_L14036_C161/carry[2] ),.C1(\add_105_I10_L14036_C161/carry[3] ),.SO(N316));
  HADDX1 desc152(.A0(N306),.B0(\add_105_I10_L14036_C161/carry[3] ),.C1(\add_105_I10_L14036_C161/carry[4] ),.SO(N317));
  HADDX1 desc153(.A0(N307),.B0(\add_105_I10_L14036_C161/carry[4] ),.C1(\add_105_I10_L14036_C161/carry[5] ),.SO(N318));
  HADDX1 desc154(.A0(N287),.B0(N286),.C1(\add_105_I9_L14036_C161/carry[2] ),.SO(N298));
  HADDX1 desc155(.A0(N288),.B0(\add_105_I9_L14036_C161/carry[2] ),.C1(\add_105_I9_L14036_C161/carry[3] ),.SO(N299));
  HADDX1 desc156(.A0(N289),.B0(\add_105_I9_L14036_C161/carry[3] ),.C1(\add_105_I9_L14036_C161/carry[4] ),.SO(N300));
  HADDX1 desc157(.A0(N290),.B0(\add_105_I9_L14036_C161/carry[4] ),.C1(\add_105_I9_L14036_C161/carry[5] ),.SO(N301));
  HADDX1 desc158(.A0(N270),.B0(N269),.C1(\add_105_I8_L14036_C161/carry[2] ),.SO(N281));
  HADDX1 desc159(.A0(N271),.B0(\add_105_I8_L14036_C161/carry[2] ),.C1(\add_105_I8_L14036_C161/carry[3] ),.SO(N282));
  HADDX1 desc160(.A0(N272),.B0(\add_105_I8_L14036_C161/carry[3] ),.C1(\add_105_I8_L14036_C161/carry[4] ),.SO(N283));
  HADDX1 desc161(.A0(n11),.B0(\add_105_I8_L14036_C161/carry[4] ),.C1(N285),.SO(N284));
  HADDX1 desc162(.A0(N253),.B0(N252),.C1(\add_105_I7_L14036_C161/carry[2] ),.SO(N264));
  HADDX1 desc163(.A0(N254),.B0(\add_105_I7_L14036_C161/carry[2] ),.C1(\add_105_I7_L14036_C161/carry[3] ),.SO(N265));
  HADDX1 desc164(.A0(n8),.B0(\add_105_I7_L14036_C161/carry[3] ),.C1(N267),.SO(N266));
  HADDX1 desc165(.A0(n16),.B0(N236),.C1(\add_105_I6_L14036_C161/carry[2] ),.SO(N247));
  HADDX1 desc166(.A0(N238),.B0(\add_105_I6_L14036_C161/carry[2] ),.C1(N249),.SO(N248));
  NAND2X0 U9(.IN1(N308),.IN2(n150),.QN(n116));
  NBUFFX2 U10(.INP(n428),.Z(n26));
  AND2X1 U11(.IN1(n309),.IN2(n310),.Q(n1));
  NAND2X0 U12(.IN1(n219),.IN2(n293),.QN(n176));
  NAND2X0 U13(.IN1(n133),.IN2(n295),.QN(n224));
  NAND2X0 U14(.IN1(n236),.IN2(n286),.QN(n185));
  NAND2X0 U15(.IN1(n186),.IN2(n288),.QN(n216));
  NAND2X0 U16(.IN1(n184),.IN2(n284),.QN(n210));
  NAND2X0 U17(.IN1(n217),.IN2(n290),.QN(n220));
  NBUFFX4 U18(.INP(n30),.Z(n19));
  NOR2X0 U19(.IN1(n234),.IN2(n144),.QN(n145));
  INVX0 U20(.INP(n220),.ZN(n282));
  INVX0 U21(.INP(N609),.ZN(N619));
  NBUFFX2 U22(.INP(n30),.Z(n18));
  INVX0 U23(.INP(n176),.ZN(n281));
  NOR2X0 U24(.IN1(n18),.IN2(n306),.QN(n240));
  INVX0 U25(.INP(n185),.ZN(n279));
  INVX0 U26(.INP(n34),.ZN(n30));
  NOR2X0 U27(.IN1(n238),.IN2(n18),.QN(s_fractb_28_o[0:0]));
  AND2X1 U28(.IN1(N285),.IN2(n286),.Q(n6));
  NOR2X0 U29(.IN1(n33),.IN2(n238),.QN(s_fracta_28_o[0:0]));
  AND4X1 U30(.IN1(n151),.IN2(n1),.IN3(n153),.IN4(n154),.Q(n7));
  NOR2X0 U31(.IN1(n139),.IN2(n140),.QN(n137));
  NOR2X0 U32(.IN1(n173),.IN2(n174),.QN(n172));
  NOR2X0 U33(.IN1(n160),.IN2(n161),.QN(n159));
  AND2X1 U34(.IN1(N249),.IN2(n284),.Q(n8));
  AND2X1 U35(.IN1(N267),.IN2(n285),.Q(n11));
  AND4X1 U36(.IN1(n116),.IN2(n117),.IN3(n118),.IN4(n119),.Q(n12));
  AND4X1 U37(.IN1(n164),.IN2(n165),.IN3(n166),.IN4(n167),.Q(n13));
  NAND2X0 U38(.IN1(n169),.IN2(n170),.QN(n168));
  NAND2X0 U39(.IN1(n156),.IN2(n157),.QN(n155));
  NAND2X0 U40(.IN1(n128),.IN2(n129),.QN(n126));
  NAND2X0 U41(.IN1(n127),.IN2(N356),.QN(n177));
  NOR2X0 U44(.IN1(n205),.IN2(n206),.QN(n204));
  NOR2X0 U45(.IN1(n191),.IN2(n192),.QN(n190));
  INVX0 U46(.INP(N592),.ZN(N603));
  NOR2X0 U47(.IN1(n234),.IN2(s_fract_sm_28[26:26]),.QN(n144));
  NAND2X1 U48(.IN1(n227),.IN2(n299),.QN(n138));
  NAND2X0 U49(.IN1(n124),.IN2(N405),.QN(n212));
  NAND2X0 U50(.IN1(n282),.IN2(n291),.QN(n218));
  NAND2X1 U51(.IN1(n225),.IN2(n297),.QN(n226));
  NAND2X1 U52(.IN1(n233),.IN2(n304),.QN(n234));
  NAND2X1 U53(.IN1(n231),.IN2(n302),.QN(n232));
  NOR2X0 U54(.IN1(n229),.IN2(n230),.QN(n228));
  INVX0 U55(.INP(N493),.ZN(n103));
  INVX0 U56(.INP(N495),.ZN(n91));
  INVX0 U57(.INP(N510),.ZN(n102));
  INVX0 U58(.INP(N511),.ZN(n96));
  INVX0 U59(.INP(N512),.ZN(n90));
  NOR2X0 U60(.IN1(n232),.IN2(n233),.QN(n142));
  NOR2X0 U61(.IN1(n148),.IN2(n231),.QN(n147));
  INVX0 U62(.INP(N425),.ZN(n107));
  INVX0 U63(.INP(N442),.ZN(n106));
  INVX0 U64(.INP(N427),.ZN(n95));
  INVX0 U65(.INP(N444),.ZN(n94));
  INVX0 U66(.INP(N426),.ZN(n101));
  INVX0 U67(.INP(N443),.ZN(n100));
  INVX0 U68(.INP(N494),.ZN(n97));
  INVX0 U69(.INP(N491),.ZN(n273));
  INVX0 U70(.INP(N492),.ZN(n267));
  INVX0 U71(.INP(N476),.ZN(n104));
  INVX0 U72(.INP(N477),.ZN(n98));
  INVX0 U73(.INP(N474),.ZN(n274));
  INVX0 U74(.INP(N475),.ZN(n268));
  INVX0 U75(.INP(N478),.ZN(n92));
  INVX0 U76(.INP(N459),.ZN(n105));
  INVX0 U77(.INP(N460),.ZN(n99));
  INVX0 U78(.INP(N457),.ZN(n275));
  INVX0 U79(.INP(N508),.ZN(n272));
  INVX0 U80(.INP(N509),.ZN(n266));
  INVX0 U81(.INP(N461),.ZN(n93));
  NAND2X0 U82(.IN1(n227),.IN2(n138),.QN(n136));
  NAND2X1 U83(.IN1(n225),.IN2(n226),.QN(n131));
  NAND2X0 U84(.IN1(n124),.IN2(N406),.QN(n197));
  INVX0 U85(.INP(N423),.ZN(n277));
  INVX0 U86(.INP(N424),.ZN(n271));
  INVX0 U87(.INP(N440),.ZN(n276));
  INVX0 U88(.INP(N441),.ZN(n270));
  INVX0 U89(.INP(N458),.ZN(n269));
  INVX0 U90(.INP(s_fract_sm_28[26:26]),.ZN(n305));
  NOR2X0 U91(.IN1(n218),.IN2(n219),.QN(n123));
  NAND2X1 U92(.IN1(n133),.IN2(n224),.QN(n134));
  NAND2X0 U93(.IN1(N290),.IN2(n125),.QN(n310));
  NAND2X0 U94(.IN1(N358),.IN2(n127),.QN(n309));
  NOR2X0 U95(.IN1(n252),.IN2(n18),.QN(n241));
  NOR2X0 U96(.IN1(n306),.IN2(n33),.QN(n244));
  NOR2X0 U97(.IN1(n252),.IN2(n33),.QN(n243));
  NOR2X0 U98(.IN1(n216),.IN2(n217),.QN(n122));
  NAND2X0 U99(.IN1(n334),.IN2(n22),.QN(n354));
  NOR2X0 U100(.IN1(n185),.IN2(n186),.QN(n150));
  INVX0 U101(.INP(n252),.ZN(n306));
  NOR2X0 U102(.IN1(n210),.IN2(n236),.QN(n149));
  NAND2X0 U103(.IN1(s_fract_sm_28[26:26]),.IN2(n24),.QN(n325));
  NAND2X0 U104(.IN1(n349),.IN2(n20),.QN(n369));
  INVX0 U105(.INP(n184),.ZN(n278));
  INVX0 U106(.INP(n186),.ZN(n280));
  INVX0 U107(.INP(n381),.ZN(n265));
  INVX0 U108(.INP(n340),.ZN(n113));
  INVX0 U109(.INP(n360),.ZN(n114));
  INVX0 U110(.INP(n337),.ZN(n112));
  INVX0 U111(.INP(n338),.ZN(n264));
  INVX0 U112(.INP(n350),.ZN(n111));
  INVX0 U113(.INP(n385),.ZN(n115));
  INVX0 U114(.INP(s_fract_sm_28[5:5]),.ZN(n284));
  NBUFFX2 U115(.INP(N109),.Z(n34));
  OA21X1 U116(.IN1(n14),.IN2(n144),.IN3(n15),.Q(n238));
  AND4X1 U117(.IN1(n88),.IN2(n87),.IN3(n86),.IN4(n85),.Q(n14));
  OR2X1 U118(.IN1(n26),.IN2(n321),.Q(n15));
  INVX0 U119(.INP(N236),.ZN(N246));
  INVX0 U120(.INP(N252),.ZN(N263));
  INVX0 U121(.INP(N303),.ZN(N314));
  INVX0 U122(.INP(N286),.ZN(N297));
  INVX0 U123(.INP(s_fract_sm_28[4:4]),.ZN(n283));
  NAND2X0 U124(.IN1(s_fract_sm_28[3:3]),.IN2(s_fract_sm_28[4:4]),.QN(N238));
  INVX0 U125(.INP(s_fract_sm_28[3:3]),.ZN(N231));
  AND2X1 U126(.IN1(s_fract_sm_28[3:3]),.IN2(s_fract_sm_28[4:4]),.Q(n16));
  INVX0 U127(.INP(N269),.ZN(N280));
  INVX0 U128(.INP(N320),.ZN(N331));
  INVX0 U129(.INP(n56),.ZN(n74));
  INVX0 U130(.INP(n78),.ZN(n89));
  INVX0 U131(.INP(s_fract_sm_28[7:7]),.ZN(n286));
  NBUFFX2 U132(.INP(N109),.Z(n35));
  INVX0 U133(.INP(s_fract_sm_28[6:6]),.ZN(n285));
  INVX0 U134(.INP(N490),.ZN(N501));
  INVX0 U135(.INP(N473),.ZN(N484));
  INVX0 U136(.INP(N456),.ZN(N467));
  INVX0 U137(.INP(N405),.ZN(N416));
  INVX0 U138(.INP(s_fract_sm_28[8:8]),.ZN(n287));
  INVX0 U139(.INP(N541),.ZN(N552));
  INVX0 U140(.INP(N507),.ZN(N518));
  INVX0 U141(.INP(N575),.ZN(N586));
  INVX0 U142(.INP(N524),.ZN(N535));
  INVX0 U152(.INP(N371),.ZN(N382));
  INVX0 U153(.INP(N337),.ZN(N348));
  AOI221X1 U162(.IN1(n125),.IN2(N287),.IN3(n149),.IN4(N270),.IN5(n194),.QN(n17));
  INVX0 U164(.INP(N439),.ZN(N450));
  INVX0 U188(.INP(N422),.ZN(N433));
  INVX0 U272(.INP(N558),.ZN(N569));
  INVX0 U287(.INP(N388),.ZN(N399));
  INVX0 U294(.INP(N354),.ZN(N365));
  NOR2X0 U301(.IN1(n176),.IN2(s_fract_sm_28[15:15]),.QN(n133));
  INVX0 U308(.INP(s_fract_sm_28[11:11]),.ZN(n290));
  INVX0 U315(.INP(s_fract_sm_28[9:9]),.ZN(n288));
  INVX0 U322(.INP(s_fract_sm_28[12:12]),.ZN(n291));
  NOR2X0 U329(.IN1(n185),.IN2(s_fract_sm_28[8:8]),.QN(n186));
  NOR2X0 U336(.IN1(n148),.IN2(s_fract_sm_28[22:22]),.QN(n231));
  INVX0 U343(.INP(s_fract_sm_28[10:10]),.ZN(n289));
  NOR2X0 U406(.IN1(n210),.IN2(s_fract_sm_28[6:6]),.QN(n236));
  NOR2X0 U407(.IN1(n218),.IN2(s_fract_sm_28[13:13]),.QN(n219));
  NOR2X0 U414(.IN1(n216),.IN2(s_fract_sm_28[10:10]),.QN(n217));
  NOR2X0 U415(.IN1(s_fract_sm_28[3:3]),.IN2(s_fract_sm_28[4:4]),.QN(n184));
  NOR2X0 U421(.IN1(n224),.IN2(s_fract_sm_28[17:17]),.QN(n225));
  NOR2X0 U422(.IN1(n226),.IN2(s_fract_sm_28[19:19]),.QN(n227));
  NBUFFX2 U423(.INP(N109),.Z(n36));
  NOR2X0 U428(.IN1(n232),.IN2(s_fract_sm_28[24:24]),.QN(n233));
  INVX0 U429(.INP(s_fract_sm_28[14:14]),.ZN(n293));
  INVX0 U430(.INP(s_fract_sm_28[13:13]),.ZN(n292));
  INVX0 U431(.INP(s_fract_sm_28[15:15]),.ZN(n294));
  INVX0 U434(.INP(s_fract_sm_28[16:16]),.ZN(n295));
  INVX0 U435(.INP(s_fract_sm_28[18:18]),.ZN(n297));
  NBUFFX2 U466(.INP(N109),.Z(n37));
  INVX0 U467(.INP(s_fract_sm_28[17:17]),.ZN(n296));
  INVX0 U468(.INP(s_fract_sm_28[19:19]),.ZN(n298));
  INVX0 U469(.INP(s_fract_sm_28[20:20]),.ZN(n299));
  INVX0 U470(.INP(s_fract_sm_28[22:22]),.ZN(n301));
  INVX0 U471(.INP(s_fract_sm_28[21:21]),.ZN(n300));
  INVX0 U472(.INP(n357),.ZN(n108));
  NAND2X1 U473(.IN1(n355),.IN2(n2),.QN(n372));
  NAND2X1 U474(.IN1(n371),.IN2(n2),.QN(n425));
  NAND2X0 U475(.IN1(n357),.IN2(n2),.QN(n388));
  INVX0 U476(.INP(s_fract_sm_28[25:25]),.ZN(n304));
  INVX0 U477(.INP(s_fract_sm_28[23:23]),.ZN(n302));
  NOR2X0 U478(.IN1(n26),.IN2(n380),.QN(s_fract_shr_28[2:2]));
  NOR2X0 U479(.IN1(n26),.IN2(n365),.QN(s_fract_shr_28[1:1]));
  INVX0 U480(.INP(s_fract_sm_28[24:24]),.ZN(n303));
  NOR2X0 U481(.IN1(n26),.IN2(n327),.QN(s_fract_shr_28[10:10]));
  NOR2X0 U482(.IN1(n26),.IN2(n427),.QN(s_fract_shr_28[9:9]));
  NOR2X0 U483(.IN1(n26),.IN2(n390),.QN(s_fract_shr_28[3:3]));
  NOR2X0 U484(.IN1(n26),.IN2(n397),.QN(s_fract_shr_28[4:4]));
  NOR2X0 U485(.IN1(n26),.IN2(n410),.QN(s_fract_shr_28[6:6]));
  NOR2X0 U486(.IN1(n26),.IN2(n417),.QN(s_fract_shr_28[7:7]));
  NOR2X0 U487(.IN1(n26),.IN2(n422),.QN(s_fract_shr_28[8:8]));
  NOR2X0 U488(.IN1(n26),.IN2(n403),.QN(s_fract_shr_28[5:5]));
  INVX0 U489(.INP(n371),.ZN(n110));
  INVX0 U490(.INP(n355),.ZN(n109));
  INVX0 U491(.INP(n312),.ZN(n258));
  INVX0 U492(.INP(n311),.ZN(n152));
  INVX0 U493(.INP(n319),.ZN(n263));
  INVX0 U494(.INP(n315),.ZN(n259));
  INVX0 U495(.INP(n316),.ZN(n260));
  INVX0 U496(.INP(n318),.ZN(n262));
  INVX0 U497(.INP(n317),.ZN(n261));
  NBUFFX2 U498(.INP(N109),.Z(n33));
  NBUFFX2 U499(.INP(N109),.Z(n44));
  NBUFFX2 U500(.INP(N109),.Z(n43));
  NBUFFX2 U501(.INP(N109),.Z(n45));
  NBUFFX2 U502(.INP(N109),.Z(n38));
  NBUFFX2 U503(.INP(N109),.Z(n46));
  NBUFFX2 U504(.INP(n3),.Z(n24));
  NBUFFX2 U505(.INP(n5),.Z(n20));
  NBUFFX2 U506(.INP(n3),.Z(n25));
  NBUFFX2 U507(.INP(n5),.Z(n21));
  NBUFFX2 U508(.INP(n4),.Z(n23));
  NBUFFX2 U509(.INP(n428),.Z(n27));
  AO22X1 U510(.IN1(opb_i[0:0]),.IN2(n35),.IN3(opa_i[0:0]),.IN4(n19),.Q(s_fract_sm_28[3:3]));
  AO22X1 U511(.IN1(opb_i[5:5]),.IN2(n36),.IN3(opa_i[5:5]),.IN4(n19),.Q(s_fract_sm_28[8:8]));
  INVX0 U512(.INP(opa_i[28:28]),.ZN(n73));
  INVX0 U513(.INP(opa_i[25:25]),.ZN(n72));
  INVX0 U514(.INP(opb_i[26:26]),.ZN(n69));
  INVX0 U515(.INP(opb_i[24:24]),.ZN(n68));
  INVX0 U516(.INP(opb_i[27:27]),.ZN(n70));
  INVX0 U517(.INP(opb_i[30:30]),.ZN(n71));
  AO22X1 U518(.IN1(opb_i[14:14]),.IN2(n36),.IN3(opa_i[14:14]),.IN4(n19),.Q(s_fract_sm_28[17:17]));
  AO22X1 U519(.IN1(opb_i[16:16]),.IN2(n36),.IN3(opa_i[16:16]),.IN4(n19),.Q(s_fract_sm_28[19:19]));
  AO22X1 U520(.IN1(opb_i[15:15]),.IN2(n36),.IN3(opa_i[15:15]),.IN4(n19),.Q(s_fract_sm_28[18:18]));
  INVX0 U521(.INP(opa_i[24:24]),.ZN(n307));
  NOR2X0 U522(.IN1(opa_i[26:26]),.IN2(opa_i[25:25]),.QN(n253));
  AO22X1 U523(.IN1(opb_i[19:19]),.IN2(n37),.IN3(opa_i[19:19]),.IN4(n19),.Q(s_fract_sm_28[22:22]));
  AO22X1 U524(.IN1(opb_i[18:18]),.IN2(n37),.IN3(opa_i[18:18]),.IN4(n19),.Q(s_fract_sm_28[21:21]));
  AO22X1 U525(.IN1(opb_i[17:17]),.IN2(n37),.IN3(opa_i[17:17]),.IN4(n19),.Q(s_fract_sm_28[20:20]));
  INVX0 U526(.INP(opb_i[23:23]),.ZN(n308));
  NOR2X0 U527(.IN1(opb_i[26:26]),.IN2(opb_i[25:25]),.QN(n255));
  AO22X1 U528(.IN1(opb_i[22:22]),.IN2(n37),.IN3(opa_i[22:22]),.IN4(n31),.Q(s_fract_sm_28[25:25]));
  AO22X1 U529(.IN1(opb_i[21:21]),.IN2(n37),.IN3(opa_i[21:21]),.IN4(n19),.Q(s_fract_sm_28[24:24]));
  AO22X1 U530(.IN1(opb_i[20:20]),.IN2(n37),.IN3(opa_i[20:20]),.IN4(n19),.Q(s_fract_sm_28[23:23]));
  NOR2X0 U531(.IN1(n354),.IN2(s_exp_diff[2:2]),.QN(n371));
  NOR2X0 U532(.IN1(n345),.IN2(s_exp_diff[2:2]),.QN(n355));
  NAND2X0 U533(.IN1(s_fract_sm_28[3:3]),.IN2(s_exp_diff[0:0]),.QN(n374));
  NAND2X1 U534(.IN1(s_exp_diff[1:1]),.IN2(n383),.QN(n361));
  NBUFFX2 U535(.INP(s_exp_diff[4:4]),.Z(n29));
  NBUFFX2 U536(.INP(s_exp_diff[4:4]),.Z(n28));
  NBUFFX4 U537(.INP(n4),.Z(n22));
  NAND2X1 U538(.IN1(n67),.IN2(n66),.QN(N109));
  INVX0 U539(.INP(n34),.ZN(n31));
  INVX0 U540(.INP(n34),.ZN(n32));
  INVX0 U541(.INP(n48),.ZN(n47));
  INVX0 U542(.INP(opa_i[23:23]),.ZN(n48));
  INVX0 U543(.INP(n50),.ZN(n49));
  INVX0 U544(.INP(opa_i[29:29]),.ZN(n50));
  XOR2X1 U545(.IN1(\add_105_I9_L14036_C161/carry[5] ),.IN2(n6),.Q(N302));
  XOR2X1 U546(.IN1(\add_105_I10_L14036_C161/carry[5] ),.IN2(N308),.Q(N319));
  XOR2X1 U547(.IN1(\add_105_I11_L14036_C161/carry[5] ),.IN2(N325),.Q(N336));
  XOR2X1 U548(.IN1(\add_105_I12_L14036_C161/carry[5] ),.IN2(N342),.Q(N353));
  XOR2X1 U549(.IN1(\add_105_I13_L14036_C161/carry[5] ),.IN2(N359),.Q(N370));
  XOR2X1 U550(.IN1(\add_105_I14_L14036_C161/carry[5] ),.IN2(N376),.Q(N387));
  XOR2X1 U551(.IN1(\add_105_I15_L14036_C161/carry[5] ),.IN2(N393),.Q(N404));
  XOR2X1 U552(.IN1(\add_105_I16_L14036_C161/carry[5] ),.IN2(N410),.Q(N421));
  XOR2X1 U553(.IN1(\add_105_I17_L14036_C161/carry[5] ),.IN2(N427),.Q(N438));
  XOR2X1 U554(.IN1(\add_105_I18_L14036_C161/carry[5] ),.IN2(N444),.Q(N455));
  XOR2X1 U555(.IN1(\add_105_I19_L14036_C161/carry[5] ),.IN2(N461),.Q(N472));
  XOR2X1 U556(.IN1(\add_105_I20_L14036_C161/carry[5] ),.IN2(N478),.Q(N489));
  XOR2X1 U557(.IN1(\add_105_I21_L14036_C161/carry[5] ),.IN2(N495),.Q(N506));
  XOR2X1 U558(.IN1(\add_105_I22_L14036_C161/carry[5] ),.IN2(N512),.Q(N523));
  XOR2X1 U559(.IN1(\add_105_I23_L14036_C161/carry[5] ),.IN2(N529),.Q(N540));
  XOR2X1 U560(.IN1(\add_105_I24_L14036_C161/carry[5] ),.IN2(N546),.Q(N557));
  XOR2X1 U561(.IN1(\add_105_I25_L14036_C161/carry[5] ),.IN2(N563),.Q(N574));
  XOR2X1 U562(.IN1(\add_105_I26_L14036_C161/carry[5] ),.IN2(N580),.Q(N591));
  XOR2X1 U563(.IN1(\add_105_I27_L14036_C161/carry[5] ),.IN2(N597),.Q(N608));
  XOR2X1 U564(.IN1(\add_105_I28_L14036_C161/carry[5] ),.IN2(N614),.Q(N624));
  NAND2X0 U565(.IN1(opb_i[28:28]),.IN2(n73),.QN(n61));
  NAND3X0 U566(.IN1(n61),.IN2(n70),.IN3(opa_i[27:27]),.QN(n51));
  OA21X1 U567(.IN1(opb_i[28:28]),.IN2(n73),.IN3(n51),.Q(n55));
  NOR2X0 U568(.IN1(n71),.IN2(opa_i[30:30]),.QN(n53));
  NOR2X0 U569(.IN1(opb_i[29:29]),.IN2(n53),.QN(n52));
  AOI22X1 U570(.IN1(opa_i[30:30]),.IN2(n71),.IN3(n52),.IN4(n49),.QN(n54));
  AO21X1 U571(.IN1(opb_i[29:29]),.IN2(n50),.IN3(n53),.Q(n56));
  AO22X1 U572(.IN1(n55),.IN2(n54),.IN3(n54),.IN4(n56),.Q(n67));
  NOR2X0 U573(.IN1(opa_i[24:24]),.IN2(n68),.QN(n57));
  NOR2X0 U574(.IN1(opb_i[23:23]),.IN2(n57),.QN(n59));
  NOR2X0 U575(.IN1(n69),.IN2(opa_i[26:26]),.QN(n60));
  NOR2X0 U576(.IN1(opb_i[25:25]),.IN2(n60),.QN(n58));
  AO22X1 U577(.IN1(opa_i[26:26]),.IN2(n69),.IN3(n58),.IN4(opa_i[25:25]),.Q(n62));
  AO221X1 U578(.IN1(opa_i[24:24]),.IN2(n68),.IN3(n59),.IN4(n47),.IN5(n62),.Q(n65));
  AOI21X1 U579(.IN1(n72),.IN2(opb_i[25:25]),.IN3(n60),.QN(n63));
  OA221X1 U580(.IN1(n63),.IN2(n62),.IN3(opa_i[27:27]),.IN4(n70),.IN5(n61),.Q(n64));
  NAND3X0 U581(.IN1(n74),.IN2(n65),.IN3(n64),.QN(n66));
  NOR2X0 U582(.IN1(s_exp_diff[1:1]),.IN2(n17),.QN(n75));
  NOR2X0 U583(.IN1(s_rzeros[0:0]),.IN2(n75),.QN(n77));
  NOR2X0 U584(.IN1(n13),.IN2(s_exp_diff[3:3]),.QN(n79));
  NOR2X0 U585(.IN1(s_rzeros[2:2]),.IN2(n79),.QN(n76));
  AO22X1 U586(.IN1(s_exp_diff[3:3]),.IN2(n13),.IN3(n76),.IN4(s_exp_diff[2:2]),.Q(n78));
  AO221X1 U587(.IN1(s_exp_diff[1:1]),.IN2(n17),.IN3(n77),.IN4(s_exp_diff[0:0]),.IN5(n78),.Q(n83));
  AO21X1 U588(.IN1(s_rzeros[2:2]),.IN2(n5),.IN3(n79),.Q(n80));
  NAND2X0 U589(.IN1(n89),.IN2(n80),.QN(n82));
  OR2X1 U590(.IN1(n12),.IN2(s_exp_diff[5:5]),.Q(n84));
  OR2X1 U591(.IN1(n7),.IN2(n29),.Q(n81));
  NAND4X0 U592(.IN1(n83),.IN2(n82),.IN3(n84),.IN4(n81),.QN(n88));
  NAND3X0 U593(.IN1(n84),.IN2(n7),.IN3(n29),.QN(n87));
  NOR2X0 U594(.IN1(s_exp_diff[7:7]),.IN2(s_exp_diff[6:6]),.QN(n86));
  NAND2X0 U595(.IN1(s_exp_diff[5:5]),.IN2(n12),.QN(n85));
  OR3X1 U596(.IN1(s_exp_diff[7:7]),.IN2(s_exp_diff[6:6]),.IN3(s_exp_diff[5:5]),.Q(n428));
  MUX21X1 U597(.IN1(n294),.IN2(n293),.S(n25),.Q(n322));
  MUX21X1 U598(.IN1(n292),.IN2(n291),.S(n25),.Q(n324));
  MUX21X1 U599(.IN1(n322),.IN2(n324),.S(n22),.Q(n331));
  MUX21X1 U600(.IN1(n290),.IN2(n289),.S(n25),.Q(n323));
  MUX21X1 U601(.IN1(n288),.IN2(n287),.S(n25),.Q(n373));
  MUX21X1 U602(.IN1(n323),.IN2(n373),.S(n23),.Q(n392));
  MUX21X1 U603(.IN1(n331),.IN2(n392),.S(n21),.Q(n418));
  MUX21X1 U604(.IN1(s_fract_sm_28[7:7]),.IN2(s_fract_sm_28[6:6]),.S(n25),.Q(n311));
  MUX21X1 U605(.IN1(s_fract_sm_28[5:5]),.IN2(s_fract_sm_28[4:4]),.S(n25),.Q(n312));
  MUX21X1 U606(.IN1(n152),.IN2(n258),.S(n23),.Q(n391));
  OR2X1 U607(.IN1(n374),.IN2(n23),.Q(n313));
  MUX21X1 U608(.IN1(n391),.IN2(n313),.S(n21),.Q(n314));
  MUX21X1 U609(.IN1(n418),.IN2(n314),.S(n2),.Q(n320));
  MUX21X1 U610(.IN1(s_fract_sm_28[25:25]),.IN2(s_fract_sm_28[24:24]),.S(n25),.Q(n315));
  MUX21X1 U611(.IN1(n325),.IN2(n259),.S(n23),.Q(n330));
  OR2X1 U612(.IN1(n330),.IN2(s_exp_diff[2:2]),.Q(n370));
  MUX21X1 U613(.IN1(s_fract_sm_28[23:23]),.IN2(s_fract_sm_28[22:22]),.S(n25),.Q(n316));
  MUX21X1 U614(.IN1(s_fract_sm_28[21:21]),.IN2(s_fract_sm_28[20:20]),.S(n25),.Q(n317));
  MUX21X1 U615(.IN1(n260),.IN2(n261),.S(n23),.Q(n329));
  MUX21X1 U616(.IN1(s_fract_sm_28[19:19]),.IN2(s_fract_sm_28[18:18]),.S(n25),.Q(n318));
  MUX21X1 U617(.IN1(s_fract_sm_28[17:17]),.IN2(s_fract_sm_28[16:16]),.S(n25),.Q(n319));
  MUX21X1 U618(.IN1(n262),.IN2(n263),.S(n23),.Q(n332));
  MUX21X1 U619(.IN1(n329),.IN2(n332),.S(n21),.Q(n419));
  MUX21X1 U620(.IN1(n370),.IN2(n419),.S(n2),.Q(n353));
  MUX21X1 U621(.IN1(n320),.IN2(n353),.S(n28),.Q(n321));
  MUX21X1 U622(.IN1(n259),.IN2(n260),.S(n23),.Q(n344));
  MUX21X1 U623(.IN1(n261),.IN2(n262),.S(n23),.Q(n347));
  MUX21X1 U624(.IN1(n344),.IN2(n347),.S(n21),.Q(n356));
  MUX21X1 U625(.IN1(n263),.IN2(n322),.S(n22),.Q(n346));
  MUX21X1 U626(.IN1(n324),.IN2(n323),.S(n22),.Q(n405));
  MUX21X1 U627(.IN1(n346),.IN2(n405),.S(n21),.Q(n377));
  MUX21X1 U628(.IN1(n356),.IN2(n377),.S(n2),.Q(n326));
  OR2X1 U629(.IN1(n325),.IN2(s_exp_diff[1:1]),.Q(n345));
  MUX21X1 U630(.IN1(n326),.IN2(n372),.S(n28),.Q(n327));
  MUX21X1 U631(.IN1(s_fract_sm_28[26:26]),.IN2(s_fract_sm_28[25:25]),.S(n25),.Q(n334));
  MUX21X1 U632(.IN1(s_fract_sm_28[24:24]),.IN2(s_fract_sm_28[23:23]),.S(n24),.Q(n336));
  MUX21X1 U633(.IN1(n334),.IN2(n336),.S(n22),.Q(n349));
  MUX21X1 U634(.IN1(s_fract_sm_28[22:22]),.IN2(s_fract_sm_28[21:21]),.S(n24),.Q(n335));
  MUX21X1 U635(.IN1(s_fract_sm_28[20:20]),.IN2(s_fract_sm_28[19:19]),.S(n24),.Q(n339));
  MUX21X1 U636(.IN1(n335),.IN2(n339),.S(n22),.Q(n350));
  MUX21X1 U637(.IN1(n349),.IN2(n350),.S(n21),.Q(n357));
  MUX21X1 U638(.IN1(s_fract_sm_28[18:18]),.IN2(s_fract_sm_28[17:17]),.S(n24),.Q(n338));
  MUX21X1 U639(.IN1(n295),.IN2(n294),.S(n24),.Q(n342));
  MUX21X1 U640(.IN1(n264),.IN2(n342),.S(n22),.Q(n351));
  MUX21X1 U641(.IN1(n293),.IN2(n292),.S(n24),.Q(n341));
  MUX21X1 U642(.IN1(n291),.IN2(n290),.S(n24),.Q(n358));
  MUX21X1 U643(.IN1(n341),.IN2(n358),.S(n22),.Q(n412));
  MUX21X1 U644(.IN1(n351),.IN2(n412),.S(n21),.Q(n387));
  MUX21X1 U645(.IN1(n108),.IN2(n387),.S(n2),.Q(n328));
  NOR3X0 U646(.IN1(n27),.IN2(n28),.IN3(n328),.QN(s_fract_shr_28[11:11]));
  MUX21X1 U647(.IN1(n330),.IN2(n329),.S(n21),.Q(n366));
  MUX21X1 U648(.IN1(n332),.IN2(n331),.S(n21),.Q(n394));
  MUX21X1 U649(.IN1(n366),.IN2(n394),.S(n2),.Q(n333));
  NOR3X0 U650(.IN1(n27),.IN2(n29),.IN3(n333),.QN(s_fract_shr_28[12:12]));
  MUX21X1 U651(.IN1(n336),.IN2(n335),.S(n22),.Q(n337));
  MUX21X1 U652(.IN1(n354),.IN2(n112),.S(n21),.Q(n367));
  MUX21X1 U653(.IN1(n339),.IN2(n338),.S(n22),.Q(n340));
  MUX21X1 U654(.IN1(n342),.IN2(n341),.S(n22),.Q(n359));
  MUX21X1 U655(.IN1(n113),.IN2(n359),.S(n21),.Q(n400));
  MUX21X1 U656(.IN1(n367),.IN2(n400),.S(n2),.Q(n343));
  NOR3X0 U657(.IN1(n27),.IN2(n29),.IN3(n343),.QN(s_fract_shr_28[13:13]));
  MUX21X1 U658(.IN1(n345),.IN2(n344),.S(n21),.Q(n368));
  MUX21X1 U659(.IN1(n347),.IN2(n346),.S(n20),.Q(n407));
  MUX21X1 U660(.IN1(n368),.IN2(n407),.S(n2),.Q(n348));
  NOR3X0 U661(.IN1(n348),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[14:14]));
  MUX21X1 U662(.IN1(n111),.IN2(n351),.S(n20),.Q(n414));
  MUX21X1 U663(.IN1(n369),.IN2(n414),.S(n2),.Q(n352));
  NOR3X0 U664(.IN1(n352),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[15:15]));
  NOR3X0 U665(.IN1(n27),.IN2(n29),.IN3(n353),.QN(s_fract_shr_28[16:16]));
  MUX21X1 U666(.IN1(n112),.IN2(n113),.S(n20),.Q(n424));
  MUX21X1 U667(.IN1(n110),.IN2(n424),.S(n2),.Q(n363));
  NOR3X0 U668(.IN1(n363),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[17:17]));
  MUX21X1 U669(.IN1(n109),.IN2(n356),.S(n2),.Q(n378));
  NOR3X0 U670(.IN1(n378),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[18:18]));
  NOR3X0 U671(.IN1(n388),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[19:19]));
  MUX21X1 U672(.IN1(n289),.IN2(n288),.S(n24),.Q(n382));
  MUX21X1 U673(.IN1(n358),.IN2(n382),.S(n22),.Q(n398));
  MUX21X1 U674(.IN1(n359),.IN2(n398),.S(n20),.Q(n423));
  MUX21X1 U675(.IN1(s_fract_sm_28[8:8]),.IN2(s_fract_sm_28[7:7]),.S(n24),.Q(n381));
  MUX21X1 U676(.IN1(s_fract_sm_28[6:6]),.IN2(s_fract_sm_28[5:5]),.S(n24),.Q(n384));
  MUX21X1 U677(.IN1(n381),.IN2(n384),.S(n22),.Q(n360));
  MUX21X1 U678(.IN1(s_fract_sm_28[4:4]),.IN2(s_fract_sm_28[3:3]),.S(n24),.Q(n383));
  MUX21X1 U679(.IN1(n114),.IN2(n361),.S(n20),.Q(n362));
  MUX21X1 U680(.IN1(n423),.IN2(n362),.S(n2),.Q(n364));
  MUX21X1 U681(.IN1(n364),.IN2(n363),.S(n28),.Q(n365));
  OR2X1 U682(.IN1(n366),.IN2(s_exp_diff[3:3]),.Q(n395));
  NOR3X0 U683(.IN1(n395),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[20:20]));
  OR2X1 U684(.IN1(n367),.IN2(s_exp_diff[3:3]),.Q(n401));
  NOR3X0 U685(.IN1(n401),.IN2(n29),.IN3(n27),.QN(s_fract_shr_28[21:21]));
  OR2X1 U686(.IN1(n368),.IN2(s_exp_diff[3:3]),.Q(n408));
  NOR3X0 U687(.IN1(n27),.IN2(n29),.IN3(n408),.QN(s_fract_shr_28[22:22]));
  OR2X1 U688(.IN1(n369),.IN2(s_exp_diff[3:3]),.Q(n415));
  NOR3X0 U689(.IN1(n27),.IN2(n29),.IN3(n415),.QN(s_fract_shr_28[23:23]));
  OR2X1 U690(.IN1(n370),.IN2(s_exp_diff[3:3]),.Q(n420));
  NOR3X0 U691(.IN1(n27),.IN2(n29),.IN3(n420),.QN(s_fract_shr_28[24:24]));
  NOR3X0 U692(.IN1(n425),.IN2(n29),.IN3(n26),.QN(s_fract_shr_28[25:25]));
  NOR3X0 U693(.IN1(n372),.IN2(n28),.IN3(n26),.QN(s_fract_shr_28[26:26]));
  MUX21X1 U694(.IN1(n373),.IN2(n152),.S(n22),.Q(n404));
  MUX21X1 U695(.IN1(n258),.IN2(n374),.S(n22),.Q(n375));
  MUX21X1 U696(.IN1(n404),.IN2(n375),.S(n20),.Q(n376));
  MUX21X1 U697(.IN1(n377),.IN2(n376),.S(n2),.Q(n379));
  MUX21X1 U698(.IN1(n379),.IN2(n378),.S(n28),.Q(n380));
  MUX21X1 U699(.IN1(n382),.IN2(n265),.S(n22),.Q(n411));
  MUX21X1 U700(.IN1(n384),.IN2(n383),.S(n22),.Q(n385));
  MUX21X1 U701(.IN1(n411),.IN2(n115),.S(n20),.Q(n386));
  MUX21X1 U702(.IN1(n387),.IN2(n386),.S(n2),.Q(n389));
  MUX21X1 U703(.IN1(n389),.IN2(n388),.S(n28),.Q(n390));
  MUX21X1 U704(.IN1(n392),.IN2(n391),.S(n20),.Q(n393));
  MUX21X1 U705(.IN1(n394),.IN2(n393),.S(n2),.Q(n396));
  MUX21X1 U706(.IN1(n396),.IN2(n395),.S(n28),.Q(n397));
  MUX21X1 U707(.IN1(n398),.IN2(n114),.S(n20),.Q(n399));
  MUX21X1 U708(.IN1(n400),.IN2(n399),.S(n2),.Q(n402));
  MUX21X1 U709(.IN1(n402),.IN2(n401),.S(n28),.Q(n403));
  MUX21X1 U710(.IN1(n405),.IN2(n404),.S(n20),.Q(n406));
  MUX21X1 U711(.IN1(n407),.IN2(n406),.S(n2),.Q(n409));
  MUX21X1 U712(.IN1(n409),.IN2(n408),.S(n28),.Q(n410));
  MUX21X1 U713(.IN1(n412),.IN2(n411),.S(n20),.Q(n413));
  MUX21X1 U714(.IN1(n414),.IN2(n413),.S(n2),.Q(n416));
  MUX21X1 U715(.IN1(n416),.IN2(n415),.S(n28),.Q(n417));
  MUX21X1 U716(.IN1(n419),.IN2(n418),.S(n2),.Q(n421));
  MUX21X1 U717(.IN1(n421),.IN2(n420),.S(n28),.Q(n422));
  MUX21X1 U718(.IN1(n424),.IN2(n423),.S(n2),.Q(n426));
  MUX21X1 U719(.IN1(n426),.IN2(n425),.S(n28),.Q(n427));
assign fracta_28_o[27:27]=1'b0;
assign fractb_28_o[27:27]=1'b0;
endmodule
module addsub_28_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [27:0] A ;
input [27:0] B ;
output [27:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire [28:0] carry ;
// instances
  FADDX1 U2_26(.A(A[26:26]),.B(n27),.CI(carry[26:26]),.CO(carry[27:27]),.S(DIFF[26:26]));
  FADDX1 U2_25(.A(A[25:25]),.B(n26),.CI(carry[25:25]),.CO(carry[26:26]),.S(DIFF[25:25]));
  FADDX1 U2_24(.A(A[24:24]),.B(n25),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n24),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n23),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n22),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n21),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n20),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n19),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n18),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n17),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n16),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n15),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n14),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n13),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n12),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n11),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n10),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n9),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n8),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n7),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n6),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n5),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n4),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n3),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n2),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_27(.IN1(A[27:27]),.IN2(n28),.IN3(carry[27:27]),.Q(DIFF[27:27]));
  INVX0 U1(.INP(B[24:24]),.ZN(n25));
  INVX0 U2(.INP(B[10:10]),.ZN(n11));
  INVX0 U3(.INP(B[14:14]),.ZN(n15));
  INVX0 U4(.INP(B[18:18]),.ZN(n19));
  INVX0 U5(.INP(B[6:6]),.ZN(n7));
  INVX0 U6(.INP(B[16:16]),.ZN(n17));
  INVX0 U7(.INP(B[20:20]),.ZN(n21));
  INVX0 U8(.INP(B[22:22]),.ZN(n23));
  INVX0 U9(.INP(B[11:11]),.ZN(n12));
  INVX0 U10(.INP(B[12:12]),.ZN(n13));
  INVX0 U11(.INP(B[15:15]),.ZN(n16));
  INVX0 U12(.INP(B[17:17]),.ZN(n18));
  INVX0 U13(.INP(B[19:19]),.ZN(n20));
  INVX0 U14(.INP(B[21:21]),.ZN(n22));
  INVX0 U15(.INP(B[8:8]),.ZN(n9));
  INVX0 U16(.INP(B[23:23]),.ZN(n24));
  INVX0 U17(.INP(B[25:25]),.ZN(n26));
  INVX0 U18(.INP(B[7:7]),.ZN(n8));
  INVX0 U19(.INP(B[26:26]),.ZN(n27));
  INVX0 U20(.INP(B[3:3]),.ZN(n4));
  INVX0 U21(.INP(B[4:4]),.ZN(n5));
  INVX0 U22(.INP(B[9:9]),.ZN(n10));
  INVX0 U23(.INP(B[13:13]),.ZN(n14));
  INVX0 U24(.INP(B[5:5]),.ZN(n6));
  INVX0 U25(.INP(B[2:2]),.ZN(n3));
  INVX0 U26(.INP(B[1:1]),.ZN(n2));
  NAND2X1 U27(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U28(.INP(A[0:0]),.ZN(n1));
  INVX0 U29(.INP(B[27:27]),.ZN(n28));
  XOR2X1 U30(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module addsub_28_DW01_sub_1_inj (A,B,CI,DIFF,CO);
input [27:0] A ;
input [27:0] B ;
output [27:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire [28:0] carry ;
// instances
  FADDX1 U2_26(.A(A[26:26]),.B(n27),.CI(carry[26:26]),.CO(carry[27:27]),.S(DIFF[26:26]));
  FADDX1 U2_25(.A(A[25:25]),.B(n26),.CI(carry[25:25]),.CO(carry[26:26]),.S(DIFF[25:25]));
  FADDX1 U2_24(.A(A[24:24]),.B(n25),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n24),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n23),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n22),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n21),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n20),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n19),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n18),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n17),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n16),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n15),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n14),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n13),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n12),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n11),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n10),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n9),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n8),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n7),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n6),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n5),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n4),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n3),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n2),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_27(.IN1(A[27:27]),.IN2(n28),.IN3(carry[27:27]),.Q(DIFF[27:27]));
  INVX0 U1(.INP(B[16:16]),.ZN(n17));
  INVX0 U2(.INP(B[20:20]),.ZN(n21));
  INVX0 U3(.INP(B[18:18]),.ZN(n19));
  INVX0 U4(.INP(B[22:22]),.ZN(n23));
  INVX0 U5(.INP(B[12:12]),.ZN(n13));
  INVX0 U6(.INP(B[8:8]),.ZN(n9));
  INVX0 U7(.INP(B[10:10]),.ZN(n11));
  INVX0 U8(.INP(B[14:14]),.ZN(n15));
  INVX0 U9(.INP(B[6:6]),.ZN(n7));
  INVX0 U10(.INP(B[2:2]),.ZN(n3));
  INVX0 U11(.INP(B[26:26]),.ZN(n27));
  INVX0 U12(.INP(B[25:25]),.ZN(n26));
  INVX0 U13(.INP(B[4:4]),.ZN(n5));
  INVX0 U14(.INP(B[17:17]),.ZN(n18));
  INVX0 U15(.INP(B[21:21]),.ZN(n22));
  INVX0 U16(.INP(B[24:24]),.ZN(n25));
  INVX0 U17(.INP(B[19:19]),.ZN(n20));
  INVX0 U18(.INP(B[23:23]),.ZN(n24));
  INVX0 U19(.INP(B[3:3]),.ZN(n4));
  INVX0 U20(.INP(B[11:11]),.ZN(n12));
  INVX0 U21(.INP(B[15:15]),.ZN(n16));
  INVX0 U22(.INP(B[7:7]),.ZN(n8));
  INVX0 U23(.INP(B[1:1]),.ZN(n2));
  NAND2X1 U24(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U25(.INP(A[0:0]),.ZN(n1));
  INVX0 U26(.INP(B[9:9]),.ZN(n10));
  INVX0 U27(.INP(B[13:13]),.ZN(n14));
  INVX0 U28(.INP(B[5:5]),.ZN(n6));
  INVX0 U29(.INP(B[27:27]),.ZN(n28));
  XOR2X1 U30(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module addsub_28_DW01_add_0_inj (A,B,CI,SUM,CO);
input [27:0] A ;
input [27:0] B ;
output [27:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire [27:1] carry ;
// instances
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(carry[26:26]),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_25(.A(A[25:25]),.B(B[25:25]),.CI(carry[25:25]),.CO(carry[26:26]),.S(SUM[25:25]));
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(carry[24:24]),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(carry[13:13]),.CO(carry[14:14]),.S(SUM[13:13]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(carry[12:12]),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_11(.A(A[11:11]),.B(B[11:11]),.CI(carry[11:11]),.CO(carry[12:12]),.S(SUM[11:11]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(carry[10:10]),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_9(.A(A[9:9]),.B(B[9:9]),.CI(carry[9:9]),.CO(carry[10:10]),.S(SUM[9:9]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(carry[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  XOR3X1 U1_27(.IN1(A[27:27]),.IN2(B[27:27]),.IN3(carry[27:27]),.Q(SUM[27:27]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  XOR2X1 U2(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module addsub_28_DW_cmp_0_inj (A,B,TC,GE_LT,GE_GT_EQ,GE_LT_GT_LE,EQ_NE);
input [27:0] A ;
input [27:0] B ;
input TC ;
input GE_LT ;
input GE_GT_EQ ;
output GE_LT_GT_LE ;
output EQ_NE ;
wire n1111 ;
wire n1112 ;
wire n1113 ;
wire n1114 ;
wire n1115 ;
wire n1116 ;
wire n1117 ;
wire n1118 ;
wire n1119 ;
wire n1120 ;
wire n1121 ;
wire n1122 ;
wire n1123 ;
wire n1124 ;
wire n1125 ;
wire n1126 ;
wire n1127 ;
wire n1128 ;
wire n1129 ;
wire n1130 ;
wire n1131 ;
wire n1132 ;
wire n1133 ;
wire n1134 ;
wire n1135 ;
wire n1136 ;
wire n1137 ;
wire n1138 ;
wire n1139 ;
wire n1140 ;
wire n1141 ;
wire n1142 ;
wire n1143 ;
wire n1144 ;
wire n1145 ;
wire n1146 ;
wire n1147 ;
wire n1148 ;
wire n1149 ;
wire n1150 ;
wire n1151 ;
wire n1152 ;
wire n1153 ;
wire n1154 ;
wire n1155 ;
wire n1156 ;
wire n1157 ;
wire n1158 ;
wire n1159 ;
wire n1160 ;
wire n1161 ;
wire n1162 ;
wire n1163 ;
wire n1164 ;
wire n1165 ;
wire n1166 ;
wire n1167 ;
wire n1168 ;
wire n1169 ;
wire n1170 ;
wire n1171 ;
wire n1172 ;
wire n1173 ;
wire n1174 ;
wire n1175 ;
wire n1176 ;
wire n1177 ;
wire n1178 ;
wire n1179 ;
wire n1180 ;
wire n1181 ;
wire n1182 ;
wire n1183 ;
wire n1184 ;
wire n1185 ;
wire n1186 ;
wire n1187 ;
wire n1188 ;
wire n1189 ;
wire n1190 ;
wire n1191 ;
wire n1192 ;
wire n1193 ;
wire n1194 ;
wire n1195 ;
wire n1196 ;
wire n1197 ;
wire n1198 ;
wire n1199 ;
wire n1200 ;
wire n1201 ;
wire n1202 ;
wire n1203 ;
wire n1204 ;
wire n1205 ;
wire n1206 ;
wire n1207 ;
wire n1208 ;
wire n1209 ;
wire n1210 ;
wire n1211 ;
wire n1212 ;
wire n1213 ;
wire n1214 ;
wire n1215 ;
wire n1216 ;
wire n1217 ;
wire n1218 ;
// instances
  INVX0 U566(.INP(n1152),.ZN(n1136));
  INVX0 U567(.INP(n1183),.ZN(n1116));
  INVX0 U568(.INP(n1200),.ZN(n1142));
  INVX0 U569(.INP(n1157),.ZN(n1131));
  INVX0 U570(.INP(n1209),.ZN(n1138));
  INVX0 U571(.INP(B[20:20]),.ZN(n1137));
  INVX0 U572(.INP(n1163),.ZN(n1121));
  INVX0 U573(.INP(n1162),.ZN(n1124));
  INVX0 U574(.INP(B[14:14]),.ZN(n1128));
  INVX0 U575(.INP(B[6:6]),.ZN(n1117));
  INVX0 U576(.INP(A[1:1]),.ZN(n1111));
  INVX0 U577(.INP(A[12:12]),.ZN(n1125));
  INVX0 U578(.INP(A[8:8]),.ZN(n1119));
  INVX0 U579(.INP(A[24:24]),.ZN(n1143));
  INVX0 U580(.INP(A[25:25]),.ZN(n1144));
  INVX0 U581(.INP(A[26:26]),.ZN(n1145));
  INVX0 U582(.INP(A[4:4]),.ZN(n1114));
  INVX0 U583(.INP(A[21:21]),.ZN(n1139));
  INVX0 U584(.INP(A[17:17]),.ZN(n1132));
  INVX0 U585(.INP(A[3:3]),.ZN(n1113));
  INVX0 U586(.INP(A[23:23]),.ZN(n1141));
  INVX0 U587(.INP(A[19:19]),.ZN(n1135));
  INVX0 U588(.INP(A[11:11]),.ZN(n1123));
  INVX0 U589(.INP(A[7:7]),.ZN(n1118));
  INVX0 U590(.INP(A[15:15]),.ZN(n1129));
  INVX0 U591(.INP(B[2:2]),.ZN(n1112));
  INVX0 U592(.INP(B[9:9]),.ZN(n1120));
  INVX0 U593(.INP(B[13:13]),.ZN(n1126));
  INVX0 U594(.INP(B[5:5]),.ZN(n1115));
  INVX0 U595(.INP(n1151),.ZN(n1133));
  INVX0 U596(.INP(B[18:18]),.ZN(n1134));
  INVX0 U597(.INP(B[10:10]),.ZN(n1122));
  INVX0 U598(.INP(B[22:22]),.ZN(n1140));
  INVX0 U599(.INP(B[16:16]),.ZN(n1130));
  INVX0 U600(.INP(n1172),.ZN(n1127));
  INVX0 U601(.INP(A[27:27]),.ZN(n1146));
  AO21X1 U602(.IN1(n1147),.IN2(n1148),.IN3(n1149),.Q(GE_LT_GT_LE));
  NOR4X0 U603(.IN1(n1150),.IN2(n1151),.IN3(n1152),.IN4(n1153),.QN(n1149));
  NAND4X0 U604(.IN1(n1154),.IN2(n1155),.IN3(n1131),.IN4(n1156),.QN(n1150));
  NAND2X0 U605(.IN1(A[16:16]),.IN2(n1130),.QN(n1156));
  NAND2X0 U606(.IN1(n1158),.IN2(n1159),.QN(n1155));
  NAND4X0 U607(.IN1(n1121),.IN2(n1124),.IN3(n1160),.IN4(n1161),.QN(n1159));
  OR2X1 U608(.IN1(n1119),.IN2(B[8:8]),.Q(n1161));
  NAND3X0 U609(.IN1(n1164),.IN2(n1165),.IN3(n1158),.QN(n1154));
  AND2X1 U610(.IN1(n1166),.IN2(n1167),.Q(n1158));
  AO221X1 U611(.IN1(n1168),.IN2(n1163),.IN3(n1169),.IN4(n1168),.IN5(n1162),.Q(n1167));
  NAND3X0 U612(.IN1(n1170),.IN2(n1171),.IN3(n1127),.QN(n1162));
  OR2X1 U613(.IN1(n1125),.IN2(B[12:12]),.Q(n1171));
  OA21X1 U614(.IN1(A[9:9]),.IN2(n1120),.IN3(n1173),.Q(n1169));
  NAND3X0 U615(.IN1(n1160),.IN2(n1119),.IN3(B[8:8]),.QN(n1173));
  NAND2X0 U616(.IN1(A[9:9]),.IN2(n1120),.QN(n1160));
  AO21X1 U617(.IN1(A[10:10]),.IN2(n1122),.IN3(n1174),.Q(n1163));
  AOI22X1 U618(.IN1(B[11:11]),.IN2(n1123),.IN3(n1175),.IN4(B[10:10]),.QN(n1168));
  NOR2X0 U619(.IN1(A[10:10]),.IN2(n1174),.QN(n1175));
  NOR2X0 U620(.IN1(n1123),.IN2(B[11:11]),.QN(n1174));
  AO22X1 U621(.IN1(n1176),.IN2(n1177),.IN3(n1177),.IN4(n1172),.Q(n1166));
  AO21X1 U622(.IN1(A[14:14]),.IN2(n1128),.IN3(n1178),.Q(n1172));
  AOI22X1 U623(.IN1(B[15:15]),.IN2(n1129),.IN3(n1179),.IN4(B[14:14]),.QN(n1177));
  NOR2X0 U624(.IN1(A[14:14]),.IN2(n1178),.QN(n1179));
  NOR2X0 U625(.IN1(n1129),.IN2(B[15:15]),.QN(n1178));
  OA21X1 U626(.IN1(A[13:13]),.IN2(n1126),.IN3(n1180),.Q(n1176));
  NAND3X0 U627(.IN1(n1170),.IN2(n1125),.IN3(B[12:12]),.QN(n1180));
  NAND2X0 U628(.IN1(A[13:13]),.IN2(n1126),.QN(n1170));
  AO22X1 U629(.IN1(n1181),.IN2(n1182),.IN3(n1182),.IN4(n1183),.Q(n1165));
  AOI22X1 U630(.IN1(B[7:7]),.IN2(n1118),.IN3(n1184),.IN4(B[6:6]),.QN(n1182));
  NOR2X0 U631(.IN1(A[6:6]),.IN2(n1185),.QN(n1184));
  OA21X1 U632(.IN1(A[5:5]),.IN2(n1115),.IN3(n1186),.Q(n1181));
  NAND3X0 U633(.IN1(n1187),.IN2(n1114),.IN3(B[4:4]),.QN(n1186));
  NAND3X0 U634(.IN1(n1116),.IN2(n1188),.IN3(n1189),.QN(n1164));
  OA221X1 U635(.IN1(n1190),.IN2(n1191),.IN3(B[4:4]),.IN4(n1114),.IN5(n1187),.Q(n1189));
  NAND2X0 U636(.IN1(A[5:5]),.IN2(n1115),.QN(n1187));
  AOI21X1 U637(.IN1(n1112),.IN2(A[2:2]),.IN3(n1192),.QN(n1190));
  AO221X1 U638(.IN1(B[1:1]),.IN2(n1111),.IN3(n1193),.IN4(B[0:0]),.IN5(n1191),.Q(n1188));
  AO22X1 U639(.IN1(B[3:3]),.IN2(n1113),.IN3(n1194),.IN4(B[2:2]),.Q(n1191));
  NOR2X0 U640(.IN1(A[2:2]),.IN2(n1192),.QN(n1194));
  NOR2X0 U641(.IN1(n1113),.IN2(B[3:3]),.QN(n1192));
  NOR2X0 U642(.IN1(A[0:0]),.IN2(n1195),.QN(n1193));
  NOR2X0 U643(.IN1(B[1:1]),.IN2(n1111),.QN(n1195));
  AO21X1 U644(.IN1(A[6:6]),.IN2(n1117),.IN3(n1185),.Q(n1183));
  NOR2X0 U645(.IN1(n1118),.IN2(B[7:7]),.QN(n1185));
  NAND2X0 U646(.IN1(n1142),.IN2(n1153),.QN(n1148));
  OR4X1 U647(.IN1(n1196),.IN2(n1197),.IN3(n1198),.IN4(n1199),.Q(n1153));
  NOR2X0 U648(.IN1(n1143),.IN2(B[24:24]),.QN(n1199));
  AO221X1 U649(.IN1(n1201),.IN2(n1202),.IN3(n1203),.IN4(n1136),.IN5(n1200),.Q(n1147));
  AO22X1 U650(.IN1(B[27:27]),.IN2(n1146),.IN3(n1204),.IN4(n1205),.Q(n1200));
  AO222X1 U651(.IN1(n1206),.IN2(B[24:24]),.IN3(B[25:25]),.IN4(n1144),.IN5(B[26:26]),.IN6(n1145),.Q(n1205));
  NOR2X0 U652(.IN1(A[24:24]),.IN2(n1198),.QN(n1206));
  NOR2X0 U653(.IN1(n1144),.IN2(B[25:25]),.QN(n1198));
  NOR2X0 U654(.IN1(n1197),.IN2(n1196),.QN(n1204));
  NOR2X0 U655(.IN1(n1146),.IN2(B[27:27]),.QN(n1196));
  NOR2X0 U656(.IN1(n1145),.IN2(B[26:26]),.QN(n1197));
  NAND3X0 U657(.IN1(n1138),.IN2(n1207),.IN3(n1208),.QN(n1152));
  NAND2X0 U658(.IN1(A[20:20]),.IN2(n1137),.QN(n1207));
  OA21X1 U659(.IN1(n1133),.IN2(n1210),.IN3(n1211),.Q(n1203));
  AO221X1 U660(.IN1(B[17:17]),.IN2(n1132),.IN3(n1212),.IN4(B[16:16]),.IN5(n1210),.Q(n1211));
  NOR2X0 U661(.IN1(A[16:16]),.IN2(n1157),.QN(n1212));
  NOR2X0 U662(.IN1(n1132),.IN2(B[17:17]),.QN(n1157));
  AO22X1 U663(.IN1(B[19:19]),.IN2(n1135),.IN3(n1213),.IN4(B[18:18]),.Q(n1210));
  NOR2X0 U664(.IN1(A[18:18]),.IN2(n1214),.QN(n1213));
  AO21X1 U665(.IN1(A[18:18]),.IN2(n1134),.IN3(n1214),.Q(n1151));
  NOR2X0 U666(.IN1(n1135),.IN2(B[19:19]),.QN(n1214));
  OR2X1 U667(.IN1(n1215),.IN2(n1208),.Q(n1202));
  AOI21X1 U668(.IN1(A[22:22]),.IN2(n1140),.IN3(n1216),.QN(n1208));
  AO221X1 U669(.IN1(B[21:21]),.IN2(n1139),.IN3(n1217),.IN4(B[20:20]),.IN5(n1215),.Q(n1201));
  AO22X1 U670(.IN1(B[23:23]),.IN2(n1141),.IN3(n1218),.IN4(B[22:22]),.Q(n1215));
  NOR2X0 U671(.IN1(A[22:22]),.IN2(n1216),.QN(n1218));
  NOR2X0 U672(.IN1(n1141),.IN2(B[23:23]),.QN(n1216));
  NOR2X0 U673(.IN1(A[20:20]),.IN2(n1209),.QN(n1217));
  NOR2X0 U674(.IN1(n1139),.IN2(B[21:21]),.QN(n1209));
endmodule
module addsub_28_inj (clk_i,fpu_op_i,fracta_i,fractb_i,signa_i,signb_i,fract_o,sign_o);
input [27:0] fracta_i ;
input [27:0] fractb_i ;
output [27:0] fract_o ;
input clk_i ;
input fpu_op_i ;
input signa_i ;
input signb_i ;
output sign_o ;
wire s_sign_o ;
wire N6 ;
wire N39 ;
wire N40 ;
wire N41 ;
wire N42 ;
wire N43 ;
wire N44 ;
wire N45 ;
wire N46 ;
wire N47 ;
wire N48 ;
wire N49 ;
wire N50 ;
wire N51 ;
wire N52 ;
wire N53 ;
wire N54 ;
wire N55 ;
wire N56 ;
wire N57 ;
wire N58 ;
wire N59 ;
wire N60 ;
wire N61 ;
wire N62 ;
wire N63 ;
wire N64 ;
wire N65 ;
wire N66 ;
wire N68 ;
wire N69 ;
wire N70 ;
wire N71 ;
wire N72 ;
wire N73 ;
wire N74 ;
wire N75 ;
wire N76 ;
wire N77 ;
wire N78 ;
wire N79 ;
wire N80 ;
wire N81 ;
wire N82 ;
wire N83 ;
wire N84 ;
wire N85 ;
wire N86 ;
wire N87 ;
wire N88 ;
wire N89 ;
wire N90 ;
wire N91 ;
wire N92 ;
wire N93 ;
wire N94 ;
wire N95 ;
wire N96 ;
wire N97 ;
wire N98 ;
wire N99 ;
wire N100 ;
wire N101 ;
wire N102 ;
wire N103 ;
wire N104 ;
wire N105 ;
wire N106 ;
wire N107 ;
wire N108 ;
wire N109 ;
wire N110 ;
wire N111 ;
wire N112 ;
wire N113 ;
wire N114 ;
wire N115 ;
wire N116 ;
wire N117 ;
wire N118 ;
wire N119 ;
wire N120 ;
wire N121 ;
wire N122 ;
wire N123 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n29 ;
wire n30 ;
wire [27:0] s_fract_o ;
// instances
  DFFX1 desc167(.D(s_fract_o[27:27]),.CLK(clk_i),.Q(fract_o[27:27]));
  DFFX1 desc168(.D(s_fract_o[26:26]),.CLK(clk_i),.Q(fract_o[26:26]));
  DFFX1 desc169(.D(s_fract_o[25:25]),.CLK(clk_i),.Q(fract_o[25:25]));
  DFFX1 desc170(.D(s_fract_o[24:24]),.CLK(clk_i),.Q(fract_o[24:24]));
  DFFX1 desc171(.D(s_fract_o[23:23]),.CLK(clk_i),.Q(fract_o[23:23]));
  DFFX1 desc172(.D(s_fract_o[22:22]),.CLK(clk_i),.Q(fract_o[22:22]));
  DFFX1 desc173(.D(s_fract_o[21:21]),.CLK(clk_i),.Q(fract_o[21:21]));
  DFFX1 desc174(.D(s_fract_o[20:20]),.CLK(clk_i),.Q(fract_o[20:20]));
  DFFX1 desc175(.D(s_fract_o[19:19]),.CLK(clk_i),.Q(fract_o[19:19]));
  DFFX1 desc176(.D(s_fract_o[18:18]),.CLK(clk_i),.Q(fract_o[18:18]));
  DFFX1 desc177(.D(s_fract_o[17:17]),.CLK(clk_i),.Q(fract_o[17:17]));
  DFFX1 desc178(.D(s_fract_o[16:16]),.CLK(clk_i),.Q(fract_o[16:16]));
  DFFX1 desc179(.D(s_fract_o[15:15]),.CLK(clk_i),.Q(fract_o[15:15]));
  DFFX1 desc180(.D(s_fract_o[14:14]),.CLK(clk_i),.Q(fract_o[14:14]));
  DFFX1 desc181(.D(s_fract_o[13:13]),.CLK(clk_i),.Q(fract_o[13:13]));
  DFFX1 desc182(.D(s_fract_o[12:12]),.CLK(clk_i),.Q(fract_o[12:12]));
  DFFX1 desc183(.D(s_fract_o[11:11]),.CLK(clk_i),.Q(fract_o[11:11]));
  DFFX1 desc184(.D(s_fract_o[10:10]),.CLK(clk_i),.Q(fract_o[10:10]));
  DFFX1 desc185(.D(s_fract_o[9:9]),.CLK(clk_i),.Q(fract_o[9:9]));
  DFFX1 desc186(.D(s_fract_o[8:8]),.CLK(clk_i),.Q(fract_o[8:8]));
  DFFX1 desc187(.D(s_fract_o[7:7]),.CLK(clk_i),.Q(fract_o[7:7]));
  DFFX1 desc188(.D(s_fract_o[6:6]),.CLK(clk_i),.Q(fract_o[6:6]));
  DFFX1 desc189(.D(s_fract_o[5:5]),.CLK(clk_i),.Q(fract_o[5:5]));
  DFFX1 desc190(.D(s_fract_o[4:4]),.CLK(clk_i),.Q(fract_o[4:4]));
  DFFX1 desc191(.D(s_fract_o[3:3]),.CLK(clk_i),.Q(fract_o[3:3]));
  DFFX1 desc192(.D(s_fract_o[2:2]),.CLK(clk_i),.Q(fract_o[2:2]));
  DFFX1 desc193(.D(s_fract_o[1:1]),.CLK(clk_i),.Q(fract_o[1:1]));
  DFFX1 desc194(.D(s_fract_o[0:0]),.CLK(clk_i),.Q(fract_o[0:0]));
  DFFX1 sign_o_reg(.D(s_sign_o),.CLK(clk_i),.Q(sign_o));
  OA22X1 U16(.IN1(N6),.IN2(n16),.IN3(n29),.IN4(n13),.Q(n15));
  XOR2X1 U17(.IN1(fpu_op_i),.IN2(n30),.Q(n16));
  NOR4X0 U18(.IN1(n17),.IN2(n18),.IN3(n19),.IN4(n20),.QN(n14));
  OR4X1 U19(.IN1(s_fract_o[2:2]),.IN2(s_fract_o[3:3]),.IN3(s_fract_o[4:4]),.IN4(s_fract_o[5:5]),.Q(n20));
  OR4X1 U20(.IN1(s_fract_o[6:6]),.IN2(s_fract_o[7:7]),.IN3(s_fract_o[8:8]),.IN4(s_fract_o[9:9]),.Q(n19));
  OR4X1 U21(.IN1(s_fract_o[22:22]),.IN2(s_fract_o[23:23]),.IN3(s_fract_o[21:21]),.IN4(n21),.Q(n18));
  OR4X1 U22(.IN1(s_fract_o[27:27]),.IN2(s_fract_o[26:26]),.IN3(s_fract_o[25:25]),.IN4(s_fract_o[24:24]),.Q(n21));
  NOR4X0 U23(.IN1(n24),.IN2(s_fract_o[15:15]),.IN3(s_fract_o[17:17]),.IN4(s_fract_o[16:16]),.QN(n23));
  OR4X1 U24(.IN1(s_fract_o[18:18]),.IN2(s_fract_o[19:19]),.IN3(s_fract_o[1:1]),.IN4(s_fract_o[20:20]),.Q(n24));
  NOR4X0 U25(.IN1(n25),.IN2(n26),.IN3(s_fract_o[10:10]),.IN4(s_fract_o[0:0]),.QN(n22));
  OR4X1 U26(.IN1(s_fract_o[11:11]),.IN2(s_fract_o[12:12]),.IN3(s_fract_o[13:13]),.IN4(s_fract_o[14:14]),.Q(n25));
  AO222X1 U27(.IN1(N77),.IN2(n10),.IN3(N105),.IN4(n7),.IN5(N48),.IN6(n6),.Q(s_fract_o[9:9]));
  AO222X1 U28(.IN1(N76),.IN2(n10),.IN3(N104),.IN4(n7),.IN5(N47),.IN6(n6),.Q(s_fract_o[8:8]));
  AO222X1 U29(.IN1(N75),.IN2(n10),.IN3(N103),.IN4(n7),.IN5(N46),.IN6(n6),.Q(s_fract_o[7:7]));
  AO222X1 U30(.IN1(N74),.IN2(n10),.IN3(N102),.IN4(n7),.IN5(N45),.IN6(n6),.Q(s_fract_o[6:6]));
  AO222X1 U31(.IN1(N73),.IN2(n10),.IN3(N101),.IN4(n7),.IN5(N44),.IN6(n6),.Q(s_fract_o[5:5]));
  AO222X1 U32(.IN1(N72),.IN2(n10),.IN3(N100),.IN4(n7),.IN5(N43),.IN6(n6),.Q(s_fract_o[4:4]));
  AO222X1 U33(.IN1(N71),.IN2(n10),.IN3(N99),.IN4(n7),.IN5(N42),.IN6(n6),.Q(s_fract_o[3:3]));
  AO222X1 U34(.IN1(N70),.IN2(n10),.IN3(N98),.IN4(n7),.IN5(N41),.IN6(n6),.Q(s_fract_o[2:2]));
  AO222X1 U35(.IN1(N95),.IN2(n10),.IN3(N123),.IN4(n7),.IN5(N66),.IN6(n6),.Q(s_fract_o[27:27]));
  AO222X1 U36(.IN1(N94),.IN2(n10),.IN3(N122),.IN4(n7),.IN5(N65),.IN6(n6),.Q(s_fract_o[26:26]));
  AO222X1 U37(.IN1(N93),.IN2(n10),.IN3(N121),.IN4(n7),.IN5(N64),.IN6(n6),.Q(s_fract_o[25:25]));
  AO222X1 U38(.IN1(N92),.IN2(n10),.IN3(N120),.IN4(n7),.IN5(N63),.IN6(n6),.Q(s_fract_o[24:24]));
  AO222X1 U39(.IN1(N91),.IN2(n11),.IN3(N119),.IN4(n8),.IN5(N62),.IN6(n6),.Q(s_fract_o[23:23]));
  AO222X1 U40(.IN1(N90),.IN2(n11),.IN3(N118),.IN4(n8),.IN5(N61),.IN6(n6),.Q(s_fract_o[22:22]));
  AO222X1 U41(.IN1(N89),.IN2(n11),.IN3(N117),.IN4(n8),.IN5(N60),.IN6(n6),.Q(s_fract_o[21:21]));
  AO222X1 U42(.IN1(N88),.IN2(n11),.IN3(N116),.IN4(n8),.IN5(N59),.IN6(n6),.Q(s_fract_o[20:20]));
  AO222X1 U43(.IN1(N69),.IN2(n11),.IN3(N97),.IN4(n8),.IN5(N40),.IN6(n6),.Q(s_fract_o[1:1]));
  AO222X1 U44(.IN1(N87),.IN2(n11),.IN3(N115),.IN4(n8),.IN5(N58),.IN6(n6),.Q(s_fract_o[19:19]));
  AO222X1 U45(.IN1(N86),.IN2(n11),.IN3(N114),.IN4(n8),.IN5(N57),.IN6(n6),.Q(s_fract_o[18:18]));
  AO222X1 U46(.IN1(N85),.IN2(n11),.IN3(N113),.IN4(n8),.IN5(N56),.IN6(n6),.Q(s_fract_o[17:17]));
  AO222X1 U47(.IN1(N84),.IN2(n11),.IN3(N112),.IN4(n8),.IN5(N55),.IN6(n6),.Q(s_fract_o[16:16]));
  AO222X1 U48(.IN1(N83),.IN2(n11),.IN3(N111),.IN4(n8),.IN5(N54),.IN6(n6),.Q(s_fract_o[15:15]));
  AO222X1 U49(.IN1(N82),.IN2(n11),.IN3(N110),.IN4(n8),.IN5(N53),.IN6(n6),.Q(s_fract_o[14:14]));
  AO222X1 U50(.IN1(N81),.IN2(n11),.IN3(N109),.IN4(n8),.IN5(N52),.IN6(n6),.Q(s_fract_o[13:13]));
  AO222X1 U51(.IN1(N80),.IN2(n12),.IN3(N108),.IN4(n9),.IN5(N51),.IN6(n6),.Q(s_fract_o[12:12]));
  AO222X1 U52(.IN1(N79),.IN2(n12),.IN3(N107),.IN4(n9),.IN5(N50),.IN6(n6),.Q(s_fract_o[11:11]));
  AO222X1 U53(.IN1(N78),.IN2(n12),.IN3(N106),.IN4(n9),.IN5(N49),.IN6(n6),.Q(s_fract_o[10:10]));
  AO222X1 U54(.IN1(N68),.IN2(n12),.IN3(N96),.IN4(n9),.IN5(N39),.IN6(n6),.Q(s_fract_o[0:0]));
  addsub_28_DW01_sub_0_inj sub_119(.A(fractb_i),.B(fracta_i),.CI(1'b0),.DIFF({N123,N122,N121,N120,N119,N118,N117,N116,N115,N114,N113,N112,N111,N110,N109,N108,N107,N106,N105,N104,N103,N102,N101,N100,N99,N98,N97,N96}));
  addsub_28_DW01_sub_1_inj sub_117(.A(fracta_i),.B(fractb_i),.CI(1'b0),.DIFF({N95,N94,N93,N92,N91,N90,N89,N88,N87,N86,N85,N84,N83,N82,N81,N80,N79,N78,N77,N76,N75,N74,N73,N72,N71,N70,N69,N68}));
  addsub_28_DW01_add_0_inj add_114(.A(fracta_i),.B(fractb_i),.CI(1'b0),.SUM({N66,N65,N64,N63,N62,N61,N60,N59,N58,N57,N56,N55,N54,N53,N52,N51,N50,N49,N48,N47,N46,N45,N44,N43,N42,N41,N40,N39}));
  addsub_28_DW_cmp_0_inj lt_gt_100(.A(fractb_i),.B(fracta_i),.TC(1'b0),.GE_LT(1'b1),.GE_GT_EQ(1'b0),.GE_LT_GT_LE(N6));
  XNOR3X1 U3(.IN1(n30),.IN2(n29),.IN3(fpu_op_i),.Q(n6));
  NBUFFX2 U4(.INP(n28),.Z(n8));
  NBUFFX2 U5(.INP(n28),.Z(n7));
  NBUFFX2 U11(.INP(n27),.Z(n11));
  NBUFFX2 U12(.INP(n27),.Z(n10));
  NBUFFX2 U13(.INP(n28),.Z(n9));
  NBUFFX2 U14(.INP(n27),.Z(n12));
  INVX0 U15(.INP(N6),.ZN(n13));
  NAND2X0 U55(.IN1(n22),.IN2(n23),.QN(n17));
  NOR2X0 U56(.IN1(n29),.IN2(n30),.QN(n26));
  NOR2X0 U57(.IN1(n13),.IN2(n6),.QN(n27));
  NOR2X0 U58(.IN1(n6),.IN2(N6),.QN(n28));
  NOR2X0 U59(.IN1(n14),.IN2(n15),.QN(s_sign_o));
  INVX0 U60(.INP(signb_i),.ZN(n30));
  INVX0 U61(.INP(signa_i),.ZN(n29));
endmodule
module post_norm_addsub_DW01_inc_0_inj (A,SUM);
input [8:0] A ;
output [8:0] SUM ;
wire [8:2] carry ;
// instances
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[8:8]),.IN2(A[8:8]),.Q(SUM[8:8]));
endmodule
module post_norm_addsub_DW01_add_0_inj (A,B,CI,SUM,CO);
input [27:0] A ;
input [27:0] B ;
output [27:0] SUM ;
input CI ;
output CO ;
wire \A[0]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
// instances
  XNOR2X1 U1(.IN1(A[27:27]),.IN2(n24),.Q(SUM[27:27]));
  NAND2X0 U2(.IN1(A[26:26]),.IN2(n22),.QN(n24));
  AND2X1 U3(.IN1(A[3:3]),.IN2(B[3:3]),.Q(n1));
  AND2X1 U4(.IN1(A[4:4]),.IN2(n1),.Q(n2));
  AND2X1 U5(.IN1(A[5:5]),.IN2(n2),.Q(n3));
  AND2X1 U6(.IN1(A[6:6]),.IN2(n3),.Q(n4));
  AND2X1 U7(.IN1(A[7:7]),.IN2(n4),.Q(n5));
  AND2X1 U8(.IN1(A[8:8]),.IN2(n5),.Q(n6));
  AND2X1 U9(.IN1(A[9:9]),.IN2(n6),.Q(n7));
  AND2X1 U10(.IN1(A[10:10]),.IN2(n7),.Q(n8));
  AND2X1 U11(.IN1(A[11:11]),.IN2(n8),.Q(n9));
  AND2X1 U12(.IN1(A[12:12]),.IN2(n9),.Q(n10));
  AND2X1 U13(.IN1(A[13:13]),.IN2(n10),.Q(n11));
  AND2X1 U14(.IN1(A[14:14]),.IN2(n11),.Q(n12));
  AND2X1 U15(.IN1(A[15:15]),.IN2(n12),.Q(n13));
  AND2X1 U16(.IN1(A[16:16]),.IN2(n13),.Q(n14));
  AND2X1 U17(.IN1(A[17:17]),.IN2(n14),.Q(n15));
  AND2X1 U18(.IN1(A[18:18]),.IN2(n15),.Q(n16));
  AND2X1 U19(.IN1(A[19:19]),.IN2(n16),.Q(n17));
  AND2X1 U20(.IN1(A[20:20]),.IN2(n17),.Q(n18));
  AND2X1 U21(.IN1(A[21:21]),.IN2(n18),.Q(n19));
  AND2X1 U22(.IN1(A[23:23]),.IN2(n23),.Q(n20));
  AND2X1 U23(.IN1(A[24:24]),.IN2(n20),.Q(n21));
  AND2X1 U24(.IN1(A[25:25]),.IN2(n21),.Q(n22));
  AND2X1 U25(.IN1(A[22:22]),.IN2(n19),.Q(n23));
  XOR2X1 U26(.IN1(A[26:26]),.IN2(n22),.Q(SUM[26:26]));
  XOR2X1 U27(.IN1(A[25:25]),.IN2(n21),.Q(SUM[25:25]));
  XOR2X1 U28(.IN1(A[24:24]),.IN2(n20),.Q(SUM[24:24]));
  XOR2X1 U29(.IN1(A[23:23]),.IN2(n23),.Q(SUM[23:23]));
  XOR2X1 U30(.IN1(A[22:22]),.IN2(n19),.Q(SUM[22:22]));
  XOR2X1 U31(.IN1(A[21:21]),.IN2(n18),.Q(SUM[21:21]));
  XOR2X1 U32(.IN1(A[20:20]),.IN2(n17),.Q(SUM[20:20]));
  XOR2X1 U33(.IN1(A[19:19]),.IN2(n16),.Q(SUM[19:19]));
  XOR2X1 U34(.IN1(A[18:18]),.IN2(n15),.Q(SUM[18:18]));
  XOR2X1 U35(.IN1(A[17:17]),.IN2(n14),.Q(SUM[17:17]));
  XOR2X1 U36(.IN1(A[16:16]),.IN2(n13),.Q(SUM[16:16]));
  XOR2X1 U37(.IN1(A[15:15]),.IN2(n12),.Q(SUM[15:15]));
  XOR2X1 U38(.IN1(A[14:14]),.IN2(n11),.Q(SUM[14:14]));
  XOR2X1 U39(.IN1(A[13:13]),.IN2(n10),.Q(SUM[13:13]));
  XOR2X1 U40(.IN1(A[12:12]),.IN2(n9),.Q(SUM[12:12]));
  XOR2X1 U41(.IN1(A[11:11]),.IN2(n8),.Q(SUM[11:11]));
  XOR2X1 U42(.IN1(A[10:10]),.IN2(n7),.Q(SUM[10:10]));
  XOR2X1 U43(.IN1(A[9:9]),.IN2(n6),.Q(SUM[9:9]));
  XOR2X1 U44(.IN1(A[8:8]),.IN2(n5),.Q(SUM[8:8]));
  XOR2X1 U45(.IN1(A[7:7]),.IN2(n4),.Q(SUM[7:7]));
  XOR2X1 U46(.IN1(A[6:6]),.IN2(n3),.Q(SUM[6:6]));
  XOR2X1 U47(.IN1(A[5:5]),.IN2(n2),.Q(SUM[5:5]));
  XOR2X1 U48(.IN1(A[4:4]),.IN2(n1),.Q(SUM[4:4]));
  XOR2X1 U49(.IN1(A[3:3]),.IN2(B[3:3]),.Q(SUM[3:3]));
assign SUM[2:2]=A[2:2];
assign SUM[1:1]=A[1:1];
assign SUM[0:0]=\A[0] ;
assign \A[0] =A[0:0];
endmodule
module post_norm_addsub_inj (clk_i,opa_i,opb_i,fract_28_i,exp_i,sign_i,fpu_op_i,rmode_i,output_o,ine_o);
input [31:0] opa_i ;
input [31:0] opb_i ;
input [27:0] fract_28_i ;
input [7:0] exp_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input clk_i ;
input sign_i ;
input fpu_op_i ;
output ine_o ;
wire N160 ;
wire N162 ;
wire N169 ;
wire N170 ;
wire N171 ;
wire N172 ;
wire N174 ;
wire N175 ;
wire N176 ;
wire N177 ;
wire N184 ;
wire N185 ;
wire N186 ;
wire N187 ;
wire N188 ;
wire N190 ;
wire N191 ;
wire N192 ;
wire N193 ;
wire N194 ;
wire N201 ;
wire N202 ;
wire N203 ;
wire N204 ;
wire N205 ;
wire N206 ;
wire N207 ;
wire N208 ;
wire N209 ;
wire N210 ;
wire N211 ;
wire N218 ;
wire N219 ;
wire N220 ;
wire N221 ;
wire N222 ;
wire N223 ;
wire N224 ;
wire N225 ;
wire N226 ;
wire N227 ;
wire N228 ;
wire N229 ;
wire N235 ;
wire N236 ;
wire N237 ;
wire N238 ;
wire N239 ;
wire N240 ;
wire N241 ;
wire N242 ;
wire N243 ;
wire N244 ;
wire N245 ;
wire N246 ;
wire N252 ;
wire N253 ;
wire N254 ;
wire N255 ;
wire N256 ;
wire N257 ;
wire N258 ;
wire N259 ;
wire N260 ;
wire N261 ;
wire N262 ;
wire N263 ;
wire N269 ;
wire N270 ;
wire N271 ;
wire N272 ;
wire N273 ;
wire N274 ;
wire N275 ;
wire N276 ;
wire N277 ;
wire N278 ;
wire N279 ;
wire N280 ;
wire N286 ;
wire N287 ;
wire N288 ;
wire N289 ;
wire N290 ;
wire N291 ;
wire N292 ;
wire N293 ;
wire N294 ;
wire N295 ;
wire N296 ;
wire N297 ;
wire N303 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N308 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N313 ;
wire N314 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N324 ;
wire N325 ;
wire N326 ;
wire N327 ;
wire N328 ;
wire N329 ;
wire N330 ;
wire N331 ;
wire N337 ;
wire N338 ;
wire N339 ;
wire N340 ;
wire N341 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N345 ;
wire N346 ;
wire N347 ;
wire N348 ;
wire N354 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N361 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N365 ;
wire N371 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N377 ;
wire N378 ;
wire N379 ;
wire N380 ;
wire N381 ;
wire N382 ;
wire N388 ;
wire N389 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N394 ;
wire N395 ;
wire N396 ;
wire N397 ;
wire N398 ;
wire N399 ;
wire N405 ;
wire N406 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N411 ;
wire N412 ;
wire N413 ;
wire N414 ;
wire N415 ;
wire N416 ;
wire N422 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N433 ;
wire N439 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N450 ;
wire N456 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N462 ;
wire N463 ;
wire N464 ;
wire N465 ;
wire N466 ;
wire N467 ;
wire N473 ;
wire N474 ;
wire N475 ;
wire N476 ;
wire N477 ;
wire N478 ;
wire N479 ;
wire N480 ;
wire N481 ;
wire N482 ;
wire N483 ;
wire N484 ;
wire N490 ;
wire N491 ;
wire N492 ;
wire N493 ;
wire N494 ;
wire N495 ;
wire N496 ;
wire N497 ;
wire N498 ;
wire N499 ;
wire N500 ;
wire N501 ;
wire N507 ;
wire N508 ;
wire N509 ;
wire N510 ;
wire N511 ;
wire N512 ;
wire N513 ;
wire N514 ;
wire N515 ;
wire N516 ;
wire N517 ;
wire N518 ;
wire N524 ;
wire N525 ;
wire N526 ;
wire N527 ;
wire N528 ;
wire N529 ;
wire N530 ;
wire N531 ;
wire N532 ;
wire N533 ;
wire N534 ;
wire N535 ;
wire N541 ;
wire N542 ;
wire N543 ;
wire N544 ;
wire N545 ;
wire N546 ;
wire \s_shr1[0]  ;
wire N920 ;
wire N921 ;
wire N922 ;
wire N923 ;
wire N924 ;
wire N925 ;
wire N950 ;
wire N951 ;
wire N952 ;
wire N953 ;
wire N954 ;
wire N955 ;
wire N957 ;
wire N958 ;
wire N959 ;
wire N960 ;
wire N961 ;
wire N962 ;
wire N963 ;
wire N971 ;
wire N972 ;
wire N973 ;
wire N974 ;
wire N975 ;
wire N976 ;
wire N977 ;
wire N978 ;
wire N979 ;
wire N980 ;
wire N981 ;
wire N982 ;
wire N983 ;
wire N984 ;
wire N985 ;
wire N986 ;
wire N987 ;
wire N988 ;
wire N989 ;
wire N990 ;
wire N991 ;
wire N992 ;
wire N993 ;
wire N994 ;
wire N995 ;
wire N996 ;
wire N997 ;
wire N998 ;
wire N999 ;
wire N1000 ;
wire N1001 ;
wire N1002 ;
wire N1003 ;
wire N1004 ;
wire N1005 ;
wire N1006 ;
wire N1007 ;
wire N1008 ;
wire N1009 ;
wire N1010 ;
wire N1011 ;
wire N1012 ;
wire N1013 ;
wire N1014 ;
wire N1015 ;
wire N1016 ;
wire N1017 ;
wire N1018 ;
wire N1019 ;
wire N1020 ;
wire N1021 ;
wire N1022 ;
wire N1023 ;
wire N1024 ;
wire N1025 ;
wire N1026 ;
wire N1027 ;
wire N1028 ;
wire N1029 ;
wire N1030 ;
wire N1031 ;
wire N1032 ;
wire N1033 ;
wire N1034 ;
wire N1035 ;
wire N1036 ;
wire N1037 ;
wire N1038 ;
wire N1039 ;
wire N1040 ;
wire N1041 ;
wire N1042 ;
wire N1043 ;
wire N1044 ;
wire N1045 ;
wire N1046 ;
wire N1047 ;
wire N1048 ;
wire N1049 ;
wire N1050 ;
wire N1051 ;
wire N1052 ;
wire N1053 ;
wire N1054 ;
wire s_roundup ;
wire N1092 ;
wire N1093 ;
wire N1094 ;
wire N1095 ;
wire N1096 ;
wire N1097 ;
wire N1098 ;
wire N1099 ;
wire N1100 ;
wire N1176 ;
wire n39 ;
wire n40 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire \sub_172_aco/carry[7]  ;
wire \sub_172_aco/carry[6]  ;
wire \sub_172_aco/carry[5]  ;
wire \sub_172_aco/carry[4]  ;
wire \sub_172_aco/carry[3]  ;
wire \sub_172_aco/carry[2]  ;
wire \sub_172_aco/carry[1]  ;
wire \add_90_I27_L14036_C129/carry[5]  ;
wire \add_90_I27_L14036_C129/carry[4]  ;
wire \add_90_I27_L14036_C129/carry[3]  ;
wire \add_90_I27_L14036_C129/carry[2]  ;
wire \add_90_I26_L14036_C129/carry[5]  ;
wire \add_90_I26_L14036_C129/carry[4]  ;
wire \add_90_I26_L14036_C129/carry[3]  ;
wire \add_90_I26_L14036_C129/carry[2]  ;
wire \add_90_I25_L14036_C129/carry[5]  ;
wire \add_90_I25_L14036_C129/carry[4]  ;
wire \add_90_I25_L14036_C129/carry[3]  ;
wire \add_90_I25_L14036_C129/carry[2]  ;
wire \add_90_I24_L14036_C129/carry[5]  ;
wire \add_90_I24_L14036_C129/carry[4]  ;
wire \add_90_I24_L14036_C129/carry[3]  ;
wire \add_90_I24_L14036_C129/carry[2]  ;
wire \add_90_I23_L14036_C129/carry[5]  ;
wire \add_90_I23_L14036_C129/carry[4]  ;
wire \add_90_I23_L14036_C129/carry[3]  ;
wire \add_90_I23_L14036_C129/carry[2]  ;
wire \add_90_I22_L14036_C129/carry[5]  ;
wire \add_90_I22_L14036_C129/carry[4]  ;
wire \add_90_I22_L14036_C129/carry[3]  ;
wire \add_90_I22_L14036_C129/carry[2]  ;
wire \add_90_I21_L14036_C129/carry[5]  ;
wire \add_90_I21_L14036_C129/carry[4]  ;
wire \add_90_I21_L14036_C129/carry[3]  ;
wire \add_90_I21_L14036_C129/carry[2]  ;
wire \add_90_I20_L14036_C129/carry[5]  ;
wire \add_90_I20_L14036_C129/carry[4]  ;
wire \add_90_I20_L14036_C129/carry[3]  ;
wire \add_90_I20_L14036_C129/carry[2]  ;
wire \add_90_I19_L14036_C129/carry[5]  ;
wire \add_90_I19_L14036_C129/carry[4]  ;
wire \add_90_I19_L14036_C129/carry[3]  ;
wire \add_90_I19_L14036_C129/carry[2]  ;
wire \add_90_I18_L14036_C129/carry[5]  ;
wire \add_90_I18_L14036_C129/carry[4]  ;
wire \add_90_I18_L14036_C129/carry[3]  ;
wire \add_90_I18_L14036_C129/carry[2]  ;
wire \add_90_I17_L14036_C129/carry[5]  ;
wire \add_90_I17_L14036_C129/carry[4]  ;
wire \add_90_I17_L14036_C129/carry[3]  ;
wire \add_90_I17_L14036_C129/carry[2]  ;
wire \add_90_I16_L14036_C129/carry[5]  ;
wire \add_90_I16_L14036_C129/carry[4]  ;
wire \add_90_I16_L14036_C129/carry[3]  ;
wire \add_90_I16_L14036_C129/carry[2]  ;
wire \add_90_I15_L14036_C129/carry[5]  ;
wire \add_90_I15_L14036_C129/carry[4]  ;
wire \add_90_I15_L14036_C129/carry[3]  ;
wire \add_90_I15_L14036_C129/carry[2]  ;
wire \add_90_I14_L14036_C129/carry[5]  ;
wire \add_90_I14_L14036_C129/carry[4]  ;
wire \add_90_I14_L14036_C129/carry[3]  ;
wire \add_90_I14_L14036_C129/carry[2]  ;
wire \add_90_I13_L14036_C129/carry[5]  ;
wire \add_90_I13_L14036_C129/carry[4]  ;
wire \add_90_I13_L14036_C129/carry[3]  ;
wire \add_90_I13_L14036_C129/carry[2]  ;
wire \add_90_I12_L14036_C129/carry[5]  ;
wire \add_90_I12_L14036_C129/carry[4]  ;
wire \add_90_I12_L14036_C129/carry[3]  ;
wire \add_90_I12_L14036_C129/carry[2]  ;
wire \add_90_I11_L14036_C129/carry[5]  ;
wire \add_90_I11_L14036_C129/carry[4]  ;
wire \add_90_I11_L14036_C129/carry[3]  ;
wire \add_90_I11_L14036_C129/carry[2]  ;
wire \add_90_I10_L14036_C129/carry[5]  ;
wire \add_90_I10_L14036_C129/carry[4]  ;
wire \add_90_I10_L14036_C129/carry[3]  ;
wire \add_90_I10_L14036_C129/carry[2]  ;
wire \add_90_I9_L14036_C129/carry[5]  ;
wire \add_90_I9_L14036_C129/carry[4]  ;
wire \add_90_I9_L14036_C129/carry[3]  ;
wire \add_90_I9_L14036_C129/carry[2]  ;
wire \add_90_I8_L14036_C129/carry[5]  ;
wire \add_90_I8_L14036_C129/carry[4]  ;
wire \add_90_I8_L14036_C129/carry[3]  ;
wire \add_90_I8_L14036_C129/carry[2]  ;
wire \add_90_I7_L14036_C129/carry[4]  ;
wire \add_90_I7_L14036_C129/carry[3]  ;
wire \add_90_I7_L14036_C129/carry[2]  ;
wire \add_90_I6_L14036_C129/carry[2]  ;
wire \add_90_I6_L14036_C129/carry[3]  ;
wire \add_90_I5_L14036_C129/carry[2]  ;
wire \add_90_I5_L14036_C129/A[1]  ;
wire \sub_0_root_add_0_root_sub_132/carry[8]  ;
wire \sub_0_root_add_0_root_sub_132/carry[7]  ;
wire \sub_0_root_add_0_root_sub_132/carry[6]  ;
wire \sub_0_root_add_0_root_sub_132/carry[5]  ;
wire \sub_0_root_add_0_root_sub_132/carry[4]  ;
wire \sub_0_root_add_0_root_sub_132/carry[3]  ;
wire \sub_0_root_add_0_root_sub_132/carry[2]  ;
wire \sub_0_root_add_0_root_sub_132/carry[1]  ;
wire \sub_0_root_add_0_root_sub_132/B[2]  ;
wire \sub_0_root_add_0_root_sub_132/B[5]  ;
wire \sub_0_root_add_0_root_sub_132/A[0]  ;
wire \sub_0_root_add_0_root_sub_132/A[1]  ;
wire \sub_0_root_add_0_root_sub_132/A[2]  ;
wire \sub_0_root_add_0_root_sub_132/A[3]  ;
wire \sub_0_root_add_0_root_sub_132/A[4]  ;
wire \sub_0_root_add_0_root_sub_132/A[5]  ;
wire \sub_0_root_add_0_root_sub_132/A[6]  ;
wire \sub_0_root_add_0_root_sub_132/A[7]  ;
wire \sub_0_root_add_0_root_sub_132/A[8]  ;
wire \add_1_root_add_0_root_sub_132/carry[7]  ;
wire \add_1_root_add_0_root_sub_132/carry[6]  ;
wire \add_1_root_add_0_root_sub_132/carry[5]  ;
wire \add_1_root_add_0_root_sub_132/carry[4]  ;
wire \add_1_root_add_0_root_sub_132/carry[3]  ;
wire \add_1_root_add_0_root_sub_132/carry[2]  ;
wire \add_1_root_add_0_root_sub_132/carry[1]  ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n126 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n381 ;
wire n382 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n404 ;
wire n405 ;
wire n406 ;
wire n407 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n416 ;
wire n417 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire n429 ;
wire n430 ;
wire n431 ;
wire n432 ;
wire n433 ;
wire n434 ;
wire n435 ;
wire n436 ;
wire n437 ;
wire n438 ;
wire n439 ;
wire n440 ;
wire n441 ;
wire n442 ;
wire n443 ;
wire n444 ;
wire n445 ;
wire n446 ;
wire n447 ;
wire n448 ;
wire n449 ;
wire n450 ;
wire n451 ;
wire [31:0] s_output_o ;
wire [5:0] s_zeros ;
wire [9:0] s_exp10 ;
wire [5:0] s_shl1 ;
wire [8:0] s_expo9_1 ;
wire [27:0] s_fracto28_1 ;
wire [8:0] s_expo9_2 ;
wire [27:0] s_fracto28_rnd ;
// instances
  DFFX1 desc195(.D(s_output_o[31:31]),.CLK(clk_i),.Q(output_o[31:31]));
  DFFX1 desc196(.D(N963),.CLK(clk_i),.Q(s_expo9_1[7:7]));
  DFFX1 desc197(.D(N962),.CLK(clk_i),.Q(s_expo9_1[6:6]));
  DFFX1 desc198(.D(N961),.CLK(clk_i),.Q(s_expo9_1[5:5]));
  DFFX1 desc199(.D(N960),.CLK(clk_i),.Q(s_expo9_1[4:4]));
  DFFX1 desc200(.D(N959),.CLK(clk_i),.Q(s_expo9_1[3:3]));
  DFFX1 desc201(.D(N958),.CLK(clk_i),.Q(s_expo9_1[2:2]));
  DFFX1 desc202(.D(N957),.CLK(clk_i),.Q(s_expo9_1[1:1]));
  DFFSSRX1 desc203(.D(s_exp10[0:0]),.RSTB(1'b1),.SETB(n155),.CLK(clk_i),.Q(s_expo9_1[0:0]));
  DFFSSRX1 desc204(.D(fract_28_i[27:27]),.RSTB(n155),.SETB(1'b1),.CLK(clk_i),.Q(\s_shr1[0] ),.QN(n10));
  DFFX1 desc205(.D(N955),.CLK(clk_i),.Q(s_shl1[5:5]));
  DFFX1 desc206(.D(N954),.CLK(clk_i),.Q(s_shl1[4:4]));
  DFFX1 desc207(.D(N953),.CLK(clk_i),.Q(n2),.QN(n6));
  DFFX1 desc208(.D(N952),.CLK(clk_i),.Q(n3),.QN(n9));
  DFFX1 desc209(.D(N951),.CLK(clk_i),.Q(n5),.QN(n7));
  DFFX1 desc210(.D(N950),.CLK(clk_i),.Q(n4),.QN(n8));
  DFFX1 desc211(.D(N1054),.CLK(clk_i),.Q(s_fracto28_1[27:27]));
  DFFX1 desc212(.D(N1053),.CLK(clk_i),.Q(s_fracto28_1[26:26]));
  DFFX1 desc213(.D(N1052),.CLK(clk_i),.Q(s_fracto28_1[25:25]));
  DFFX1 desc214(.D(N1051),.CLK(clk_i),.Q(s_fracto28_1[24:24]));
  DFFX1 desc215(.D(N1050),.CLK(clk_i),.Q(s_fracto28_1[23:23]));
  DFFX1 desc216(.D(N1049),.CLK(clk_i),.Q(s_fracto28_1[22:22]));
  DFFX1 desc217(.D(N1048),.CLK(clk_i),.Q(s_fracto28_1[21:21]));
  DFFX1 desc218(.D(N1047),.CLK(clk_i),.Q(s_fracto28_1[20:20]));
  DFFX1 desc219(.D(N1046),.CLK(clk_i),.Q(s_fracto28_1[19:19]));
  DFFX1 desc220(.D(N1045),.CLK(clk_i),.Q(s_fracto28_1[18:18]));
  DFFX1 desc221(.D(N1044),.CLK(clk_i),.Q(s_fracto28_1[17:17]));
  DFFX1 desc222(.D(N1043),.CLK(clk_i),.Q(s_fracto28_1[16:16]));
  DFFX1 desc223(.D(N1042),.CLK(clk_i),.Q(s_fracto28_1[15:15]));
  DFFX1 desc224(.D(N1041),.CLK(clk_i),.Q(s_fracto28_1[14:14]));
  DFFX1 desc225(.D(N1040),.CLK(clk_i),.Q(s_fracto28_1[13:13]));
  DFFX1 desc226(.D(N1039),.CLK(clk_i),.Q(s_fracto28_1[12:12]));
  DFFX1 desc227(.D(N1038),.CLK(clk_i),.Q(s_fracto28_1[11:11]));
  DFFX1 desc228(.D(N1037),.CLK(clk_i),.Q(s_fracto28_1[10:10]));
  DFFX1 desc229(.D(N1036),.CLK(clk_i),.Q(s_fracto28_1[9:9]));
  DFFX1 desc230(.D(N1035),.CLK(clk_i),.Q(s_fracto28_1[8:8]));
  DFFX1 desc231(.D(N1034),.CLK(clk_i),.Q(s_fracto28_1[7:7]));
  DFFX1 desc232(.D(N1033),.CLK(clk_i),.Q(s_fracto28_1[6:6]));
  DFFX1 desc233(.D(N1032),.CLK(clk_i),.Q(s_fracto28_1[5:5]));
  DFFX1 desc234(.D(N1031),.CLK(clk_i),.Q(s_fracto28_1[4:4]));
  DFFX1 desc235(.D(N1030),.CLK(clk_i),.Q(s_fracto28_1[3:3]),.QN(n39));
  DFFX1 desc236(.D(N1029),.CLK(clk_i),.Q(s_fracto28_1[2:2]),.QN(n40));
  DFFX1 desc237(.D(N1028),.CLK(clk_i),.Q(s_fracto28_1[1:1]));
  DFFX1 desc238(.D(N1027),.CLK(clk_i),.Q(s_fracto28_1[0:0]));
  DFFX1 ine_o_reg(.D(N1176),.CLK(clk_i),.Q(ine_o));
  DFFX1 desc239(.D(s_output_o[9:9]),.CLK(clk_i),.Q(output_o[9:9]));
  DFFX1 desc240(.D(s_output_o[8:8]),.CLK(clk_i),.Q(output_o[8:8]));
  DFFX1 desc241(.D(s_output_o[7:7]),.CLK(clk_i),.Q(output_o[7:7]));
  DFFX1 desc242(.D(s_output_o[6:6]),.CLK(clk_i),.Q(output_o[6:6]));
  DFFX1 desc243(.D(s_output_o[5:5]),.CLK(clk_i),.Q(output_o[5:5]));
  DFFX1 desc244(.D(s_output_o[4:4]),.CLK(clk_i),.Q(output_o[4:4]));
  DFFX1 desc245(.D(s_output_o[3:3]),.CLK(clk_i),.Q(output_o[3:3]));
  DFFX1 desc246(.D(s_output_o[2:2]),.CLK(clk_i),.Q(output_o[2:2]));
  DFFX1 desc247(.D(s_output_o[21:21]),.CLK(clk_i),.Q(output_o[21:21]));
  DFFX1 desc248(.D(s_output_o[20:20]),.CLK(clk_i),.Q(output_o[20:20]));
  DFFX1 desc249(.D(s_output_o[1:1]),.CLK(clk_i),.Q(output_o[1:1]));
  DFFX1 desc250(.D(s_output_o[19:19]),.CLK(clk_i),.Q(output_o[19:19]));
  DFFX1 desc251(.D(s_output_o[18:18]),.CLK(clk_i),.Q(output_o[18:18]));
  DFFX1 desc252(.D(s_output_o[17:17]),.CLK(clk_i),.Q(output_o[17:17]));
  DFFX1 desc253(.D(s_output_o[16:16]),.CLK(clk_i),.Q(output_o[16:16]));
  DFFX1 desc254(.D(s_output_o[15:15]),.CLK(clk_i),.Q(output_o[15:15]));
  DFFX1 desc255(.D(s_output_o[14:14]),.CLK(clk_i),.Q(output_o[14:14]));
  DFFX1 desc256(.D(s_output_o[13:13]),.CLK(clk_i),.Q(output_o[13:13]));
  DFFX1 desc257(.D(s_output_o[12:12]),.CLK(clk_i),.Q(output_o[12:12]));
  DFFX1 desc258(.D(s_output_o[11:11]),.CLK(clk_i),.Q(output_o[11:11]));
  DFFX1 desc259(.D(s_output_o[10:10]),.CLK(clk_i),.Q(output_o[10:10]));
  DFFX1 desc260(.D(s_output_o[0:0]),.CLK(clk_i),.Q(output_o[0:0]));
  DFFX1 desc261(.D(s_output_o[22:22]),.CLK(clk_i),.Q(output_o[22:22]));
  DFFX1 desc262(.D(s_output_o[30:30]),.CLK(clk_i),.Q(output_o[30:30]));
  DFFX1 desc263(.D(s_output_o[29:29]),.CLK(clk_i),.Q(output_o[29:29]));
  DFFX1 desc264(.D(s_output_o[28:28]),.CLK(clk_i),.Q(output_o[28:28]));
  DFFX1 desc265(.D(s_output_o[27:27]),.CLK(clk_i),.Q(output_o[27:27]));
  DFFX1 desc266(.D(s_output_o[26:26]),.CLK(clk_i),.Q(output_o[26:26]));
  DFFX1 desc267(.D(s_output_o[25:25]),.CLK(clk_i),.Q(output_o[25:25]));
  DFFX1 desc268(.D(s_output_o[24:24]),.CLK(clk_i),.Q(output_o[24:24]));
  DFFX1 desc269(.D(s_output_o[23:23]),.CLK(clk_i),.Q(output_o[23:23]));
  AO22X1 U143(.IN1(n107),.IN2(n40),.IN3(n108),.IN4(n109),.Q(n106));
  NAND3X0 U144(.IN1(rmode_i[1:1]),.IN2(n110),.IN3(sign_i),.QN(n109));
  OR2X1 U145(.IN1(n110),.IN2(sign_i),.Q(n108));
  NAND4X0 U146(.IN1(s_fracto28_1[2:2]),.IN2(n111),.IN3(n327),.IN4(n326),.QN(n105));
  NOR3X0 U147(.IN1(s_fracto28_1[1:1]),.IN2(s_fracto28_1[0:0]),.IN3(n112),.QN(n107));
  AO22X1 U148(.IN1(s_fracto28_rnd[13:13]),.IN2(n113),.IN3(s_fracto28_rnd[12:12]),.IN4(n114),.Q(s_output_o[9:9]));
  AO22X1 U149(.IN1(n113),.IN2(s_fracto28_rnd[12:12]),.IN3(s_fracto28_rnd[11:11]),.IN4(n21),.Q(s_output_o[8:8]));
  AO22X1 U150(.IN1(s_fracto28_rnd[11:11]),.IN2(n113),.IN3(s_fracto28_rnd[10:10]),.IN4(n114),.Q(s_output_o[7:7]));
  AO22X1 U151(.IN1(s_fracto28_rnd[10:10]),.IN2(n113),.IN3(s_fracto28_rnd[9:9]),.IN4(n21),.Q(s_output_o[6:6]));
  AO22X1 U152(.IN1(s_fracto28_rnd[9:9]),.IN2(n113),.IN3(s_fracto28_rnd[8:8]),.IN4(n114),.Q(s_output_o[5:5]));
  AO22X1 U153(.IN1(s_fracto28_rnd[8:8]),.IN2(n113),.IN3(s_fracto28_rnd[7:7]),.IN4(n21),.Q(s_output_o[4:4]));
  AO22X1 U154(.IN1(s_fracto28_rnd[7:7]),.IN2(n113),.IN3(s_fracto28_rnd[6:6]),.IN4(n114),.Q(s_output_o[3:3]));
  AO22X1 U155(.IN1(sign_i),.IN2(n115),.IN3(n324),.IN4(n116),.Q(s_output_o[31:31]));
  AO22X1 U156(.IN1(opa_i[31:31]),.IN2(n325),.IN3(opb_i[31:31]),.IN4(n117),.Q(n116));
  NAND3X0 U157(.IN1(n325),.IN2(n120),.IN3(n121),.QN(n119));
  AO221X1 U158(.IN1(n122),.IN2(s_expo9_2[7:7]),.IN3(n123),.IN4(N1099),.IN5(n57),.Q(s_output_o[30:30]));
  AO22X1 U159(.IN1(s_fracto28_rnd[6:6]),.IN2(n113),.IN3(s_fracto28_rnd[5:5]),.IN4(n21),.Q(s_output_o[2:2]));
  AO221X1 U160(.IN1(n122),.IN2(s_expo9_2[6:6]),.IN3(n123),.IN4(N1098),.IN5(n57),.Q(s_output_o[29:29]));
  AO221X1 U161(.IN1(n122),.IN2(s_expo9_2[5:5]),.IN3(n123),.IN4(N1097),.IN5(n57),.Q(s_output_o[28:28]));
  AO221X1 U162(.IN1(n122),.IN2(s_expo9_2[4:4]),.IN3(n123),.IN4(N1096),.IN5(n57),.Q(s_output_o[27:27]));
  AO221X1 U163(.IN1(n122),.IN2(s_expo9_2[3:3]),.IN3(n123),.IN4(N1095),.IN5(n57),.Q(s_output_o[26:26]));
  AO221X1 U164(.IN1(n122),.IN2(s_expo9_2[2:2]),.IN3(n123),.IN4(N1094),.IN5(n57),.Q(s_output_o[25:25]));
  AO221X1 U165(.IN1(n122),.IN2(s_expo9_2[1:1]),.IN3(n123),.IN4(N1093),.IN5(n57),.Q(s_output_o[24:24]));
  AO221X1 U166(.IN1(n122),.IN2(s_expo9_2[0:0]),.IN3(n123),.IN4(N1092),.IN5(n57),.Q(s_output_o[23:23]));
  AND2X1 U167(.IN1(s_fracto28_rnd[27:27]),.IN2(n125),.Q(n123));
  AND2X1 U168(.IN1(n125),.IN2(n60),.Q(n122));
  AO22X1 U170(.IN1(s_fracto28_rnd[26:26]),.IN2(s_fracto28_rnd[27:27]),.IN3(s_fracto28_rnd[25:25]),.IN4(n60),.Q(n127));
  AO21X1 U171(.IN1(n121),.IN2(n128),.IN3(n325),.Q(n118));
  NAND4X0 U172(.IN1(n131),.IN2(n132),.IN3(n133),.IN4(n134),.QN(n130));
  NOR4X0 U173(.IN1(n135),.IN2(opa_i[4:4]),.IN3(opa_i[6:6]),.IN4(opa_i[5:5]),.QN(n134));
  OR3X1 U174(.IN1(opa_i[9:9]),.IN2(opa_i[8:8]),.IN3(opa_i[7:7]),.Q(n135));
  NOR4X0 U175(.IN1(n136),.IN2(opa_i[1:1]),.IN3(opa_i[21:21]),.IN4(opa_i[20:20]),.QN(n133));
  OR3X1 U176(.IN1(opa_i[3:3]),.IN2(opa_i[2:2]),.IN3(opa_i[22:22]),.Q(n136));
  NOR4X0 U177(.IN1(n137),.IN2(opa_i[14:14]),.IN3(opa_i[16:16]),.IN4(opa_i[15:15]),.QN(n132));
  OR3X1 U178(.IN1(opa_i[19:19]),.IN2(opa_i[18:18]),.IN3(opa_i[17:17]),.Q(n137));
  NOR4X0 U179(.IN1(n138),.IN2(opa_i[11:11]),.IN3(opa_i[13:13]),.IN4(opa_i[12:12]),.QN(n131));
  OR2X1 U180(.IN1(opa_i[10:10]),.IN2(opa_i[0:0]),.Q(n138));
  AO21X1 U181(.IN1(n129),.IN2(n139),.IN3(n120),.Q(n128));
  NAND4X0 U182(.IN1(n140),.IN2(n141),.IN3(n142),.IN4(n143),.QN(n120));
  NOR4X0 U183(.IN1(n144),.IN2(opb_i[4:4]),.IN3(opb_i[6:6]),.IN4(opb_i[5:5]),.QN(n143));
  OR3X1 U184(.IN1(opb_i[9:9]),.IN2(opb_i[8:8]),.IN3(opb_i[7:7]),.Q(n144));
  NOR4X0 U185(.IN1(n145),.IN2(opb_i[1:1]),.IN3(opb_i[21:21]),.IN4(opb_i[20:20]),.QN(n142));
  OR3X1 U186(.IN1(opb_i[3:3]),.IN2(opb_i[2:2]),.IN3(opb_i[22:22]),.Q(n145));
  NOR4X0 U187(.IN1(n146),.IN2(opb_i[14:14]),.IN3(opb_i[16:16]),.IN4(opb_i[15:15]),.QN(n141));
  OR3X1 U188(.IN1(opb_i[19:19]),.IN2(opb_i[18:18]),.IN3(opb_i[17:17]),.Q(n146));
  NOR4X0 U189(.IN1(n147),.IN2(opb_i[11:11]),.IN3(opb_i[13:13]),.IN4(opb_i[12:12]),.QN(n140));
  OR2X1 U190(.IN1(opb_i[10:10]),.IN2(opb_i[0:0]),.Q(n147));
  XOR3X1 U191(.IN1(opb_i[31:31]),.IN2(opa_i[31:31]),.IN3(fpu_op_i),.Q(n139));
  AO22X1 U192(.IN1(s_fracto28_rnd[25:25]),.IN2(n113),.IN3(s_fracto28_rnd[24:24]),.IN4(n114),.Q(s_output_o[21:21]));
  AO22X1 U193(.IN1(s_fracto28_rnd[24:24]),.IN2(n113),.IN3(s_fracto28_rnd[23:23]),.IN4(n21),.Q(s_output_o[20:20]));
  AO22X1 U194(.IN1(s_fracto28_rnd[5:5]),.IN2(n113),.IN3(s_fracto28_rnd[4:4]),.IN4(n114),.Q(s_output_o[1:1]));
  AO22X1 U195(.IN1(s_fracto28_rnd[23:23]),.IN2(n113),.IN3(s_fracto28_rnd[22:22]),.IN4(n21),.Q(s_output_o[19:19]));
  AO22X1 U196(.IN1(s_fracto28_rnd[22:22]),.IN2(n113),.IN3(s_fracto28_rnd[21:21]),.IN4(n114),.Q(s_output_o[18:18]));
  AO22X1 U197(.IN1(s_fracto28_rnd[21:21]),.IN2(n113),.IN3(s_fracto28_rnd[20:20]),.IN4(n21),.Q(s_output_o[17:17]));
  AO22X1 U198(.IN1(s_fracto28_rnd[20:20]),.IN2(n113),.IN3(s_fracto28_rnd[19:19]),.IN4(n114),.Q(s_output_o[16:16]));
  AO22X1 U199(.IN1(s_fracto28_rnd[19:19]),.IN2(n113),.IN3(s_fracto28_rnd[18:18]),.IN4(n21),.Q(s_output_o[15:15]));
  AO22X1 U200(.IN1(s_fracto28_rnd[18:18]),.IN2(n113),.IN3(s_fracto28_rnd[17:17]),.IN4(n114),.Q(s_output_o[14:14]));
  AO22X1 U201(.IN1(s_fracto28_rnd[17:17]),.IN2(n113),.IN3(s_fracto28_rnd[16:16]),.IN4(n21),.Q(s_output_o[13:13]));
  AO22X1 U202(.IN1(s_fracto28_rnd[16:16]),.IN2(n113),.IN3(s_fracto28_rnd[15:15]),.IN4(n114),.Q(s_output_o[12:12]));
  AO22X1 U203(.IN1(s_fracto28_rnd[15:15]),.IN2(n113),.IN3(s_fracto28_rnd[14:14]),.IN4(n21),.Q(s_output_o[11:11]));
  AO22X1 U204(.IN1(s_fracto28_rnd[14:14]),.IN2(n113),.IN3(s_fracto28_rnd[13:13]),.IN4(n114),.Q(s_output_o[10:10]));
  AO22X1 U205(.IN1(s_fracto28_rnd[4:4]),.IN2(n113),.IN3(s_fracto28_rnd[3:3]),.IN4(n21),.Q(s_output_o[0:0]));
  AND2X1 U208(.IN1(n124),.IN2(n125),.Q(n148));
  NAND4X0 U209(.IN1(n149),.IN2(n150),.IN3(s_zeros[1:1]),.IN4(n151),.QN(n125));
  AND3X1 U210(.IN1(s_zeros[3:3]),.IN2(s_zeros[0:0]),.IN3(s_zeros[4:4]),.Q(n151));
  NOR3X0 U211(.IN1(n121),.IN2(n129),.IN3(n152),.QN(n124));
  AO21X1 U212(.IN1(s_exp10[7:7]),.IN2(n153),.IN3(n154),.Q(N963));
  AO21X1 U213(.IN1(s_exp10[6:6]),.IN2(n153),.IN3(n154),.Q(N962));
  AO21X1 U214(.IN1(s_exp10[5:5]),.IN2(n153),.IN3(n154),.Q(N961));
  AO21X1 U215(.IN1(s_exp10[4:4]),.IN2(n153),.IN3(n154),.Q(N960));
  AO21X1 U216(.IN1(s_exp10[3:3]),.IN2(n153),.IN3(n154),.Q(N959));
  AO21X1 U217(.IN1(s_exp10[2:2]),.IN2(n153),.IN3(n154),.Q(N958));
  AO21X1 U218(.IN1(s_exp10[1:1]),.IN2(n153),.IN3(n154),.Q(N957));
  AND2X1 U219(.IN1(s_exp10[8:8]),.IN2(n153),.Q(n154));
  AO22X1 U220(.IN1(\sub_0_root_add_0_root_sub_132/B[5] ),.IN2(n155),.IN3(N925),.IN4(n156),.Q(N955));
  AO221X1 U221(.IN1(n159),.IN2(N246),.IN3(n160),.IN4(n161),.IN5(n162),.Q(n158));
  AO22X1 U222(.IN1(n163),.IN2(N229),.IN3(n164),.IN4(n12),.Q(n162));
  NAND3X0 U223(.IN1(n165),.IN2(n166),.IN3(n167),.QN(n161));
  AOI222X1 U224(.IN1(n168),.IN2(N297),.IN3(n169),.IN4(N348),.IN5(n170),.IN6(n171),.QN(n167));
  NAND3X0 U225(.IN1(n172),.IN2(n173),.IN3(n174),.QN(n171));
  OA222X1 U226(.IN1(n52),.IN2(n175),.IN3(n49),.IN4(n176),.IN5(n177),.IN6(n178),.Q(n174));
  AO222X1 U227(.IN1(n181),.IN2(N484),.IN3(n16),.IN4(N467),.IN5(n182),.IN6(N501),.Q(n180));
  AO222X1 U228(.IN1(N546),.IN2(n318),.IN3(n183),.IN4(N518),.IN5(n184),.IN6(N535),.Q(n179));
  AOI22X1 U229(.IN1(N365),.IN2(n18),.IN3(N382),.IN4(n185),.QN(n173));
  OA22X1 U230(.IN1(n51),.IN2(n186),.IN3(n50),.IN4(n187),.Q(n172));
  AOI22X1 U231(.IN1(N263),.IN2(n20),.IN3(N280),.IN4(n188),.QN(n166));
  AOI22X1 U232(.IN1(N314),.IN2(n189),.IN3(N331),.IN4(n190),.QN(n165));
  AO22X1 U233(.IN1(n155),.IN2(s_zeros[4:4]),.IN3(N924),.IN4(n156),.Q(N954));
  AND2X1 U234(.IN1(n157),.IN2(n191),.Q(s_zeros[4:4]));
  AO221X1 U235(.IN1(n160),.IN2(n192),.IN3(n193),.IN4(N194),.IN5(n194),.Q(n191));
  AO222X1 U236(.IN1(n163),.IN2(N228),.IN3(n164),.IN4(N211),.IN5(n159),.IN6(N245),.Q(n194));
  NAND3X0 U237(.IN1(n195),.IN2(n196),.IN3(n197),.QN(n192));
  AOI222X1 U238(.IN1(n168),.IN2(N296),.IN3(n169),.IN4(N347),.IN5(n170),.IN6(n198),.QN(n197));
  NAND3X0 U239(.IN1(n199),.IN2(n200),.IN3(n201),.QN(n198));
  OA222X1 U240(.IN1(n56),.IN2(n175),.IN3(n53),.IN4(n176),.IN5(n202),.IN6(n178),.Q(n201));
  AO222X1 U241(.IN1(n181),.IN2(N483),.IN3(n16),.IN4(N466),.IN5(n182),.IN6(N500),.Q(n204));
  AO222X1 U242(.IN1(N545),.IN2(n318),.IN3(n183),.IN4(N517),.IN5(n184),.IN6(N534),.Q(n203));
  AOI22X1 U243(.IN1(N364),.IN2(n18),.IN3(N381),.IN4(n185),.QN(n200));
  OA22X1 U244(.IN1(n55),.IN2(n186),.IN3(n54),.IN4(n187),.Q(n199));
  AOI22X1 U245(.IN1(N262),.IN2(n20),.IN3(N279),.IN4(n188),.QN(n196));
  AOI22X1 U246(.IN1(N313),.IN2(n189),.IN3(N330),.IN4(n190),.QN(n195));
  AO22X1 U247(.IN1(n155),.IN2(s_zeros[3:3]),.IN3(N923),.IN4(n156),.Q(N953));
  AND2X1 U248(.IN1(n157),.IN2(n205),.Q(s_zeros[3:3]));
  AO221X1 U249(.IN1(n160),.IN2(n206),.IN3(n193),.IN4(N193),.IN5(n207),.Q(n205));
  AO222X1 U250(.IN1(n163),.IN2(N227),.IN3(n164),.IN4(N210),.IN5(n159),.IN6(N244),.Q(n207));
  NAND3X0 U251(.IN1(n208),.IN2(n209),.IN3(n210),.QN(n206));
  AOI222X1 U252(.IN1(n168),.IN2(N295),.IN3(n169),.IN4(N346),.IN5(n170),.IN6(n211),.QN(n210));
  NAND3X0 U253(.IN1(n212),.IN2(n213),.IN3(n214),.QN(n211));
  OA222X1 U254(.IN1(n91),.IN2(n175),.IN3(n88),.IN4(n176),.IN5(n215),.IN6(n178),.Q(n214));
  AO222X1 U255(.IN1(n181),.IN2(N482),.IN3(n16),.IN4(N465),.IN5(n182),.IN6(N499),.Q(n217));
  AO222X1 U256(.IN1(N544),.IN2(n318),.IN3(n183),.IN4(N516),.IN5(n184),.IN6(N533),.Q(n216));
  AOI22X1 U257(.IN1(N363),.IN2(n18),.IN3(N380),.IN4(n185),.QN(n213));
  OA22X1 U258(.IN1(n90),.IN2(n186),.IN3(n89),.IN4(n187),.Q(n212));
  AOI22X1 U259(.IN1(N261),.IN2(n20),.IN3(N278),.IN4(n188),.QN(n209));
  AOI22X1 U260(.IN1(N312),.IN2(n189),.IN3(N329),.IN4(n190),.QN(n208));
  AO22X1 U261(.IN1(\sub_0_root_add_0_root_sub_132/B[2] ),.IN2(n155),.IN3(N922),.IN4(n156),.Q(N952));
  AO21X1 U262(.IN1(n218),.IN2(n219),.IN3(n220),.Q(n149));
  AOI222X1 U263(.IN1(N226),.IN2(n163),.IN3(n221),.IN4(n222),.IN5(N209),.IN6(n164),.QN(n219));
  AOI222X1 U264(.IN1(N192),.IN2(n193),.IN3(N243),.IN4(n159),.IN5(n223),.IN6(n160),.QN(n218));
  OR2X1 U265(.IN1(n224),.IN2(n225),.Q(n223));
  AO222X1 U266(.IN1(n170),.IN2(n226),.IN3(n169),.IN4(N345),.IN5(n168),.IN6(N294),.Q(n225));
  NAND3X0 U267(.IN1(n227),.IN2(n228),.IN3(n229),.QN(n226));
  OA222X1 U268(.IN1(n95),.IN2(n175),.IN3(n92),.IN4(n176),.IN5(n230),.IN6(n178),.Q(n229));
  AO222X1 U269(.IN1(n181),.IN2(N481),.IN3(n16),.IN4(N464),.IN5(n182),.IN6(N498),.Q(n232));
  AO222X1 U270(.IN1(N543),.IN2(n318),.IN3(n183),.IN4(N515),.IN5(n184),.IN6(N532),.Q(n231));
  AOI22X1 U271(.IN1(N362),.IN2(n18),.IN3(N379),.IN4(n185),.QN(n228));
  OA22X1 U272(.IN1(n94),.IN2(n186),.IN3(n93),.IN4(n187),.Q(n227));
  AO221X1 U273(.IN1(n189),.IN2(N311),.IN3(n190),.IN4(N328),.IN5(n233),.Q(n224));
  AO22X1 U274(.IN1(n188),.IN2(N277),.IN3(n20),.IN4(N260),.Q(n233));
  AO22X1 U275(.IN1(n155),.IN2(s_zeros[1:1]),.IN3(N921),.IN4(n156),.Q(N951));
  AO22X1 U276(.IN1(n86),.IN2(n234),.IN3(fract_28_i[24:24]),.IN4(n157),.Q(s_zeros[1:1]));
  NAND4X0 U277(.IN1(n235),.IN2(n236),.IN3(n237),.IN4(n238),.QN(n234));
  AOI222X1 U278(.IN1(N242),.IN2(n159),.IN3(N208),.IN4(n164),.IN5(N225),.IN6(n163),.QN(n238));
  AO21X1 U279(.IN1(n239),.IN2(n240),.IN3(n101),.Q(n236));
  AOI221X1 U280(.IN1(N327),.IN2(n190),.IN3(N310),.IN4(n189),.IN5(n241),.QN(n240));
  AO22X1 U281(.IN1(N259),.IN2(n20),.IN3(N276),.IN4(n188),.Q(n241));
  AOI222X1 U282(.IN1(n168),.IN2(N293),.IN3(n169),.IN4(N344),.IN5(n170),.IN6(n242),.QN(n239));
  NAND3X0 U283(.IN1(n243),.IN2(n244),.IN3(n245),.QN(n242));
  OA222X1 U284(.IN1(n99),.IN2(n175),.IN3(n96),.IN4(n176),.IN5(n246),.IN6(n178),.Q(n245));
  AO222X1 U285(.IN1(n181),.IN2(N480),.IN3(n16),.IN4(N463),.IN5(n182),.IN6(N497),.Q(n248));
  AO222X1 U286(.IN1(N542),.IN2(n318),.IN3(n183),.IN4(N514),.IN5(n184),.IN6(N531),.Q(n247));
  AOI22X1 U287(.IN1(N361),.IN2(n18),.IN3(N378),.IN4(n185),.QN(n244));
  OA22X1 U288(.IN1(n98),.IN2(n186),.IN3(n97),.IN4(n187),.Q(n243));
  AO22X1 U289(.IN1(n155),.IN2(s_zeros[0:0]),.IN3(N920),.IN4(n156),.Q(N950));
  AOI21X1 U290(.IN1(n249),.IN2(n250),.IN3(n153),.QN(n156));
  NOR4X0 U291(.IN1(exp_i[7:7]),.IN2(exp_i[6:6]),.IN3(exp_i[5:5]),.IN4(exp_i[4:4]),.QN(n250));
  NOR4X0 U292(.IN1(exp_i[3:3]),.IN2(exp_i[2:2]),.IN3(exp_i[1:1]),.IN4(exp_i[0:0]),.QN(n249));
  AO22X1 U293(.IN1(n86),.IN2(n251),.IN3(n252),.IN4(n253),.Q(s_zeros[0:0]));
  NAND4X0 U294(.IN1(n254),.IN2(n255),.IN3(N169),.IN4(n256),.QN(n251));
  AOI222X1 U295(.IN1(N241),.IN2(n159),.IN3(N207),.IN4(n164),.IN5(N224),.IN6(n163),.QN(n256));
  AND2X1 U296(.IN1(n257),.IN2(n258),.Q(n163));
  AO21X1 U297(.IN1(n260),.IN2(n261),.IN3(n101),.Q(n255));
  AOI221X1 U298(.IN1(N326),.IN2(n190),.IN3(N309),.IN4(n189),.IN5(n262),.QN(n261));
  AO22X1 U299(.IN1(N258),.IN2(n20),.IN3(N275),.IN4(n188),.Q(n262));
  AND2X1 U300(.IN1(n265),.IN2(n266),.Q(n190));
  AOI222X1 U301(.IN1(n168),.IN2(N292),.IN3(n169),.IN4(N343),.IN5(n170),.IN6(n267),.QN(n260));
  NAND3X0 U302(.IN1(n268),.IN2(n269),.IN3(n270),.QN(n267));
  OA222X1 U303(.IN1(N405),.IN2(n175),.IN3(N456),.IN4(n176),.IN5(n271),.IN6(n178),.Q(n270));
  AO222X1 U304(.IN1(n181),.IN2(N479),.IN3(n16),.IN4(N462),.IN5(n182),.IN6(N496),.Q(n273));
  AND2X1 U305(.IN1(n274),.IN2(n275),.Q(n182));
  AO222X1 U306(.IN1(N541),.IN2(n318),.IN3(n183),.IN4(N513),.IN5(n184),.IN6(N530),.Q(n272));
  AND2X1 U307(.IN1(n276),.IN2(n277),.Q(n184));
  NAND3X0 U308(.IN1(n323),.IN2(n322),.IN3(n276),.QN(n277));
  AOI22X1 U309(.IN1(N360),.IN2(n18),.IN3(N377),.IN4(n185),.QN(n269));
  OA22X1 U310(.IN1(N422),.IN2(n186),.IN3(N439),.IN4(n187),.Q(n268));
  OR2X1 U311(.IN1(n280),.IN2(n281),.Q(n186));
  AND2X1 U312(.IN1(n263),.IN2(n264),.Q(n168));
  AND2X1 U313(.IN1(n102),.IN2(n259),.Q(n193));
  AND2X1 U314(.IN1(n282),.IN2(n87),.Q(n157));
  NOR4X0 U315(.IN1(n284),.IN2(n285),.IN3(s_exp10[5:5]),.IN4(s_exp10[4:4]),.QN(n283));
  OR3X1 U316(.IN1(s_exp10[7:7]),.IN2(s_exp10[8:8]),.IN3(s_exp10[6:6]),.Q(n285));
  OR4X1 U317(.IN1(s_exp10[0:0]),.IN2(s_exp10[1:1]),.IN3(s_exp10[2:2]),.IN4(s_exp10[3:3]),.Q(n284));
  AO22X1 U318(.IN1(N529),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N518),.Q(N535));
  AO22X1 U319(.IN1(N528),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N517),.Q(N534));
  AO22X1 U320(.IN1(N527),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N516),.Q(N533));
  AO22X1 U321(.IN1(N526),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N515),.Q(N532));
  AO22X1 U322(.IN1(N525),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N514),.Q(N531));
  AO22X1 U323(.IN1(N524),.IN2(n322),.IN3(fract_28_i[1:1]),.IN4(N513),.Q(N530));
  AO22X1 U324(.IN1(N512),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N501),.Q(N518));
  AO22X1 U325(.IN1(N511),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N500),.Q(N517));
  AO22X1 U326(.IN1(N510),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N499),.Q(N516));
  AO22X1 U327(.IN1(N509),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N498),.Q(N515));
  AO22X1 U328(.IN1(N508),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N497),.Q(N514));
  AO22X1 U329(.IN1(N507),.IN2(n321),.IN3(fract_28_i[2:2]),.IN4(N496),.Q(N513));
  AO22X1 U330(.IN1(N495),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N484),.Q(N501));
  AO22X1 U331(.IN1(N494),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N483),.Q(N500));
  AO22X1 U332(.IN1(N493),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N482),.Q(N499));
  AO22X1 U333(.IN1(N492),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N481),.Q(N498));
  AO22X1 U334(.IN1(N491),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N480),.Q(N497));
  AO22X1 U335(.IN1(N490),.IN2(n320),.IN3(fract_28_i[3:3]),.IN4(N479),.Q(N496));
  AO22X1 U336(.IN1(N478),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N467),.Q(N484));
  AO22X1 U337(.IN1(N477),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N466),.Q(N483));
  AO22X1 U338(.IN1(N476),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N465),.Q(N482));
  AO22X1 U339(.IN1(N475),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N464),.Q(N481));
  AO22X1 U340(.IN1(N474),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N463),.Q(N480));
  AO22X1 U341(.IN1(N473),.IN2(n319),.IN3(fract_28_i[4:4]),.IN4(N462),.Q(N479));
  AO22X1 U342(.IN1(N461),.IN2(n317),.IN3(n16),.IN4(N450),.Q(N467));
  AO22X1 U343(.IN1(N460),.IN2(n317),.IN3(n16),.IN4(N449),.Q(N466));
  AO22X1 U344(.IN1(N459),.IN2(n317),.IN3(n16),.IN4(N448),.Q(N465));
  AO22X1 U345(.IN1(N458),.IN2(n317),.IN3(n16),.IN4(N447),.Q(N464));
  AO22X1 U346(.IN1(N457),.IN2(n317),.IN3(n16),.IN4(N446),.Q(N463));
  AO22X1 U347(.IN1(N456),.IN2(n317),.IN3(n16),.IN4(N445),.Q(N462));
  AO22X1 U348(.IN1(N444),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N433),.Q(N450));
  AO22X1 U349(.IN1(N443),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N432),.Q(N449));
  AO22X1 U350(.IN1(N442),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N431),.Q(N448));
  AO22X1 U351(.IN1(N441),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N430),.Q(N447));
  AO22X1 U352(.IN1(N440),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N429),.Q(N446));
  AO22X1 U353(.IN1(N439),.IN2(n316),.IN3(fract_28_i[6:6]),.IN4(N428),.Q(N445));
  AO22X1 U354(.IN1(N427),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N416),.Q(N433));
  AO22X1 U355(.IN1(N426),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N415),.Q(N432));
  AO22X1 U356(.IN1(N425),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N414),.Q(N431));
  AO22X1 U357(.IN1(N424),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N413),.Q(N430));
  AO22X1 U358(.IN1(N423),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N412),.Q(N429));
  AO22X1 U359(.IN1(N422),.IN2(n315),.IN3(fract_28_i[7:7]),.IN4(N411),.Q(N428));
  AO22X1 U360(.IN1(N410),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N399),.Q(N416));
  AO22X1 U361(.IN1(N409),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N398),.Q(N415));
  AO22X1 U362(.IN1(N408),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N397),.Q(N414));
  AO22X1 U363(.IN1(N407),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N396),.Q(N413));
  AO22X1 U364(.IN1(N406),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N395),.Q(N412));
  AO22X1 U365(.IN1(N405),.IN2(n314),.IN3(fract_28_i[8:8]),.IN4(N394),.Q(N411));
  AO22X1 U366(.IN1(N393),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N382),.Q(N399));
  AO22X1 U367(.IN1(N392),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N381),.Q(N398));
  AO22X1 U368(.IN1(N391),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N380),.Q(N397));
  AO22X1 U369(.IN1(N390),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N379),.Q(N396));
  AO22X1 U370(.IN1(N389),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N378),.Q(N395));
  AO22X1 U371(.IN1(N388),.IN2(n313),.IN3(fract_28_i[9:9]),.IN4(N377),.Q(N394));
  AO22X1 U372(.IN1(N376),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N365),.Q(N382));
  AO22X1 U373(.IN1(N375),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N364),.Q(N381));
  AO22X1 U374(.IN1(N374),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N363),.Q(N380));
  AO22X1 U375(.IN1(N373),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N362),.Q(N379));
  AO22X1 U376(.IN1(N372),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N361),.Q(N378));
  AO22X1 U377(.IN1(N371),.IN2(n312),.IN3(fract_28_i[10:10]),.IN4(N360),.Q(N377));
  AO22X1 U378(.IN1(N359),.IN2(n310),.IN3(n18),.IN4(N348),.Q(N365));
  AO22X1 U379(.IN1(N358),.IN2(n310),.IN3(n18),.IN4(N347),.Q(N364));
  AO22X1 U380(.IN1(N357),.IN2(n310),.IN3(n18),.IN4(N346),.Q(N363));
  AO22X1 U381(.IN1(N356),.IN2(n310),.IN3(n18),.IN4(N345),.Q(N362));
  AO22X1 U382(.IN1(N355),.IN2(n310),.IN3(n18),.IN4(N344),.Q(N361));
  AO22X1 U383(.IN1(N354),.IN2(n310),.IN3(n18),.IN4(N343),.Q(N360));
  AO22X1 U384(.IN1(N342),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N331),.Q(N348));
  AO22X1 U385(.IN1(N341),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N330),.Q(N347));
  AO22X1 U386(.IN1(N340),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N329),.Q(N346));
  AO22X1 U387(.IN1(N339),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N328),.Q(N345));
  AO22X1 U388(.IN1(N338),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N327),.Q(N344));
  AO22X1 U389(.IN1(N337),.IN2(n309),.IN3(fract_28_i[12:12]),.IN4(N326),.Q(N343));
  AO22X1 U390(.IN1(N325),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N314),.Q(N331));
  AO22X1 U391(.IN1(N324),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N313),.Q(N330));
  AO22X1 U392(.IN1(N323),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N312),.Q(N329));
  AO22X1 U393(.IN1(N322),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N311),.Q(N328));
  AO22X1 U394(.IN1(N321),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N310),.Q(N327));
  AO22X1 U395(.IN1(N320),.IN2(n308),.IN3(fract_28_i[13:13]),.IN4(N309),.Q(N326));
  AO22X1 U396(.IN1(N308),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N297),.Q(N314));
  AO22X1 U397(.IN1(N307),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N296),.Q(N313));
  AO22X1 U398(.IN1(N306),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N295),.Q(N312));
  AO22X1 U399(.IN1(N305),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N294),.Q(N311));
  AO22X1 U400(.IN1(N304),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N293),.Q(N310));
  AO22X1 U401(.IN1(N303),.IN2(n307),.IN3(fract_28_i[14:14]),.IN4(N292),.Q(N309));
  AO22X1 U402(.IN1(N291),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N280),.Q(N297));
  AO22X1 U403(.IN1(N290),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N279),.Q(N296));
  AO22X1 U404(.IN1(N289),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N278),.Q(N295));
  AO22X1 U405(.IN1(N288),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N277),.Q(N294));
  AO22X1 U406(.IN1(N287),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N276),.Q(N293));
  AO22X1 U407(.IN1(N286),.IN2(n306),.IN3(fract_28_i[15:15]),.IN4(N275),.Q(N292));
  AO22X1 U408(.IN1(N274),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N263),.Q(N280));
  AO22X1 U409(.IN1(N273),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N262),.Q(N279));
  AO22X1 U410(.IN1(N272),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N261),.Q(N278));
  AO22X1 U411(.IN1(N271),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N260),.Q(N277));
  AO22X1 U412(.IN1(N270),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N259),.Q(N276));
  AO22X1 U413(.IN1(N269),.IN2(n305),.IN3(fract_28_i[16:16]),.IN4(N258),.Q(N275));
  AO22X1 U414(.IN1(N257),.IN2(n304),.IN3(n20),.IN4(N246),.Q(N263));
  AO22X1 U415(.IN1(N256),.IN2(n304),.IN3(n20),.IN4(N245),.Q(N262));
  AO22X1 U416(.IN1(N255),.IN2(n304),.IN3(n20),.IN4(N244),.Q(N261));
  AO22X1 U417(.IN1(N254),.IN2(n304),.IN3(n20),.IN4(N243),.Q(N260));
  AO22X1 U418(.IN1(N253),.IN2(n304),.IN3(n20),.IN4(N242),.Q(N259));
  AO22X1 U419(.IN1(N252),.IN2(n304),.IN3(n20),.IN4(N241),.Q(N258));
  AO22X1 U420(.IN1(N240),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N229),.Q(N246));
  AO22X1 U421(.IN1(N239),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N228),.Q(N245));
  AO22X1 U422(.IN1(N238),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N227),.Q(N244));
  AO22X1 U423(.IN1(N237),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N226),.Q(N243));
  AO22X1 U424(.IN1(N236),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N225),.Q(N242));
  AO22X1 U425(.IN1(N235),.IN2(n303),.IN3(fract_28_i[18:18]),.IN4(N224),.Q(N241));
  AO22X1 U426(.IN1(N223),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(n12),.Q(N229));
  AO22X1 U427(.IN1(N222),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(N211),.Q(N228));
  AO22X1 U428(.IN1(N221),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(N210),.Q(N227));
  AO22X1 U429(.IN1(N220),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(N209),.Q(N226));
  AO22X1 U430(.IN1(N219),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(N208),.Q(N225));
  AO22X1 U431(.IN1(N218),.IN2(n302),.IN3(fract_28_i[19:19]),.IN4(N207),.Q(N224));
  AO22X1 U433(.IN1(N205),.IN2(n126),.IN3(fract_28_i[20:20]),.IN4(N194),.Q(N211));
  AO22X1 U434(.IN1(N204),.IN2(n126),.IN3(fract_28_i[20:20]),.IN4(N193),.Q(N210));
  AO22X1 U435(.IN1(N203),.IN2(n126),.IN3(fract_28_i[20:20]),.IN4(N192),.Q(N209));
  AO22X1 U436(.IN1(N202),.IN2(n126),.IN3(fract_28_i[20:20]),.IN4(N191),.Q(N208));
  AO22X1 U437(.IN1(N201),.IN2(n126),.IN3(fract_28_i[20:20]),.IN4(N190),.Q(N207));
  AO22X1 U440(.IN1(N187),.IN2(n104),.IN3(N177),.IN4(fract_28_i[21:21]),.Q(N193));
  AO22X1 U441(.IN1(N186),.IN2(n104),.IN3(fract_28_i[21:21]),.IN4(N176),.Q(N192));
  AO22X1 U442(.IN1(N185),.IN2(n104),.IN3(fract_28_i[21:21]),.IN4(N175),.Q(N191));
  AO22X1 U443(.IN1(N184),.IN2(n104),.IN3(fract_28_i[21:21]),.IN4(N174),.Q(N190));
  AND2X1 U445(.IN1(N172),.IN2(n103),.Q(N177));
  AO22X1 U446(.IN1(N171),.IN2(n103),.IN3(fract_28_i[22:22]),.IN4(N162),.Q(N176));
  AO22X1 U447(.IN1(N170),.IN2(n103),.IN3(fract_28_i[22:22]),.IN4(\add_90_I5_L14036_C129/A[1] ),.Q(N175));
  AO22X1 U448(.IN1(N169),.IN2(n103),.IN3(fract_28_i[22:22]),.IN4(N160),.Q(N174));
  AND2X1 U450(.IN1(n286),.IN2(n287),.Q(N162));
  XNOR2X1 U451(.IN1(n286),.IN2(n287),.Q(n237));
  AO21X1 U452(.IN1(n253),.IN2(n100),.IN3(n282),.Q(n287));
  XOR2X1 U453(.IN1(n288),.IN2(fract_28_i[23:23]),.Q(N160));
  XNOR2X1 U454(.IN1(n100),.IN2(n253),.Q(n288));
  XOR2X1 U455(.IN1(fract_28_i[25:25]),.IN2(fract_28_i[26:26]),.Q(n253));
  NOR3X0 U456(.IN1(n289),.IN2(n129),.IN3(n121),.QN(N1176));
  NAND4X0 U457(.IN1(opb_i[30:30]),.IN2(opb_i[29:29]),.IN3(opb_i[28:28]),.IN4(opb_i[27:27]),.QN(n291));
  NAND4X0 U458(.IN1(opb_i[26:26]),.IN2(opb_i[25:25]),.IN3(opb_i[24:24]),.IN4(opb_i[23:23]),.QN(n290));
  NAND4X0 U459(.IN1(opa_i[30:30]),.IN2(opa_i[29:29]),.IN3(opa_i[28:28]),.IN4(opa_i[27:27]),.QN(n293));
  NAND4X0 U460(.IN1(opa_i[26:26]),.IN2(opa_i[25:25]),.IN3(opa_i[24:24]),.IN4(opa_i[23:23]),.QN(n292));
  NOR4X0 U461(.IN1(n294),.IN2(s_fracto28_rnd[0:0]),.IN3(s_fracto28_rnd[2:2]),.IN4(s_fracto28_rnd[1:1]),.QN(n289));
  AO221X1 U462(.IN1(\s_shr1[0] ),.IN2(fract_28_i[0:0]),.IN3(s_fracto28_rnd[3:3]),.IN4(s_fracto28_rnd[27:27]),.IN5(n152),.Q(n294));
  NAND4X0 U463(.IN1(s_expo9_2[3:3]),.IN2(s_expo9_2[2:2]),.IN3(n297),.IN4(n298),.QN(n296));
  AND4X1 U464(.IN1(s_expo9_2[4:4]),.IN2(s_expo9_2[5:5]),.IN3(s_expo9_2[6:6]),.IN4(s_expo9_2[7:7]),.Q(n298));
  AND3X1 U465(.IN1(s_expo9_2[1:1]),.IN2(n58),.IN3(s_expo9_2[0:0]),.Q(n297));
  NAND4X0 U466(.IN1(s_fracto28_rnd[27:27]),.IN2(N1099),.IN3(n299),.IN4(n300),.QN(n295));
  NOR4X0 U467(.IN1(n301),.IN2(n59),.IN3(N1100),.IN4(s_expo9_2[0:0]),.QN(n300));
  AND3X1 U468(.IN1(N1097),.IN2(N1096),.IN3(N1098),.Q(n299));
  AO22X1 U469(.IN1(N998),.IN2(\s_shr1[0] ),.IN3(N1026),.IN4(n10),.Q(N1054));
  AO22X1 U470(.IN1(N997),.IN2(\s_shr1[0] ),.IN3(N1025),.IN4(n10),.Q(N1053));
  AO22X1 U471(.IN1(N996),.IN2(\s_shr1[0] ),.IN3(N1024),.IN4(n10),.Q(N1052));
  AO22X1 U472(.IN1(N995),.IN2(\s_shr1[0] ),.IN3(N1023),.IN4(n10),.Q(N1051));
  AO22X1 U473(.IN1(N994),.IN2(\s_shr1[0] ),.IN3(N1022),.IN4(n10),.Q(N1050));
  AO22X1 U474(.IN1(N993),.IN2(\s_shr1[0] ),.IN3(N1021),.IN4(n10),.Q(N1049));
  AO22X1 U475(.IN1(N992),.IN2(\s_shr1[0] ),.IN3(N1020),.IN4(n10),.Q(N1048));
  AO22X1 U476(.IN1(N991),.IN2(\s_shr1[0] ),.IN3(N1019),.IN4(n10),.Q(N1047));
  AO22X1 U477(.IN1(N990),.IN2(\s_shr1[0] ),.IN3(N1018),.IN4(n10),.Q(N1046));
  AO22X1 U478(.IN1(N989),.IN2(\s_shr1[0] ),.IN3(N1017),.IN4(n10),.Q(N1045));
  AO22X1 U479(.IN1(N988),.IN2(\s_shr1[0] ),.IN3(N1016),.IN4(n10),.Q(N1044));
  AO22X1 U480(.IN1(N987),.IN2(\s_shr1[0] ),.IN3(N1015),.IN4(n10),.Q(N1043));
  AO22X1 U481(.IN1(N986),.IN2(\s_shr1[0] ),.IN3(N1014),.IN4(n10),.Q(N1042));
  AO22X1 U482(.IN1(N985),.IN2(\s_shr1[0] ),.IN3(N1013),.IN4(n10),.Q(N1041));
  AO22X1 U483(.IN1(N984),.IN2(\s_shr1[0] ),.IN3(N1012),.IN4(n10),.Q(N1040));
  AO22X1 U484(.IN1(N983),.IN2(\s_shr1[0] ),.IN3(N1011),.IN4(n10),.Q(N1039));
  AO22X1 U485(.IN1(N982),.IN2(\s_shr1[0] ),.IN3(N1010),.IN4(n10),.Q(N1038));
  AO22X1 U486(.IN1(N981),.IN2(\s_shr1[0] ),.IN3(N1009),.IN4(n10),.Q(N1037));
  AO22X1 U487(.IN1(N980),.IN2(\s_shr1[0] ),.IN3(N1008),.IN4(n33),.Q(N1036));
  AO22X1 U488(.IN1(N979),.IN2(\s_shr1[0] ),.IN3(N1007),.IN4(n33),.Q(N1035));
  AO22X1 U489(.IN1(N978),.IN2(\s_shr1[0] ),.IN3(N1006),.IN4(n33),.Q(N1034));
  AO22X1 U490(.IN1(N977),.IN2(n32),.IN3(N1005),.IN4(n33),.Q(N1033));
  AO22X1 U491(.IN1(N976),.IN2(n32),.IN3(N1004),.IN4(n33),.Q(N1032));
  AO22X1 U492(.IN1(N975),.IN2(n32),.IN3(N1003),.IN4(n33),.Q(N1031));
  AO22X1 U493(.IN1(N974),.IN2(n32),.IN3(N1002),.IN4(n33),.Q(N1030));
  AO22X1 U494(.IN1(N973),.IN2(n32),.IN3(N1001),.IN4(n33),.Q(N1029));
  AO22X1 U495(.IN1(N972),.IN2(n32),.IN3(N1000),.IN4(n33),.Q(N1028));
  AO22X1 U496(.IN1(N971),.IN2(\s_shr1[0] ),.IN3(N999),.IN4(n33),.Q(N1027));
  post_norm_addsub_DW01_inc_0_inj add_188(.A({n14,s_expo9_2[7:0]}),.SUM({N1100,N1099,N1098,N1097,N1096,N1095,N1094,N1093,N1092}));
  post_norm_addsub_DW01_add_0_inj add_182_aco(.A(s_fracto28_1),.B({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,s_roundup,1'b0,1'b0,1'b0}),.CI(1'b0),.SUM(s_fracto28_rnd));
  HADDX1 desc270(.A0(N531),.B0(N530),.C1(\add_90_I27_L14036_C129/carry[2] ),.SO(N542));
  HADDX1 desc271(.A0(N532),.B0(\add_90_I27_L14036_C129/carry[2] ),.C1(\add_90_I27_L14036_C129/carry[3] ),.SO(N543));
  HADDX1 desc272(.A0(N533),.B0(\add_90_I27_L14036_C129/carry[3] ),.C1(\add_90_I27_L14036_C129/carry[4] ),.SO(N544));
  HADDX1 desc273(.A0(N534),.B0(\add_90_I27_L14036_C129/carry[4] ),.C1(\add_90_I27_L14036_C129/carry[5] ),.SO(N545));
  HADDX1 desc274(.A0(N514),.B0(N513),.C1(\add_90_I26_L14036_C129/carry[2] ),.SO(N525));
  HADDX1 desc275(.A0(N515),.B0(\add_90_I26_L14036_C129/carry[2] ),.C1(\add_90_I26_L14036_C129/carry[3] ),.SO(N526));
  HADDX1 desc276(.A0(N516),.B0(\add_90_I26_L14036_C129/carry[3] ),.C1(\add_90_I26_L14036_C129/carry[4] ),.SO(N527));
  HADDX1 desc277(.A0(N517),.B0(\add_90_I26_L14036_C129/carry[4] ),.C1(\add_90_I26_L14036_C129/carry[5] ),.SO(N528));
  HADDX1 desc278(.A0(N497),.B0(N496),.C1(\add_90_I25_L14036_C129/carry[2] ),.SO(N508));
  HADDX1 desc279(.A0(N498),.B0(\add_90_I25_L14036_C129/carry[2] ),.C1(\add_90_I25_L14036_C129/carry[3] ),.SO(N509));
  HADDX1 desc280(.A0(N499),.B0(\add_90_I25_L14036_C129/carry[3] ),.C1(\add_90_I25_L14036_C129/carry[4] ),.SO(N510));
  HADDX1 desc281(.A0(N500),.B0(\add_90_I25_L14036_C129/carry[4] ),.C1(\add_90_I25_L14036_C129/carry[5] ),.SO(N511));
  HADDX1 desc282(.A0(N480),.B0(N479),.C1(\add_90_I24_L14036_C129/carry[2] ),.SO(N491));
  HADDX1 desc283(.A0(N481),.B0(\add_90_I24_L14036_C129/carry[2] ),.C1(\add_90_I24_L14036_C129/carry[3] ),.SO(N492));
  HADDX1 desc284(.A0(N482),.B0(\add_90_I24_L14036_C129/carry[3] ),.C1(\add_90_I24_L14036_C129/carry[4] ),.SO(N493));
  HADDX1 desc285(.A0(N483),.B0(\add_90_I24_L14036_C129/carry[4] ),.C1(\add_90_I24_L14036_C129/carry[5] ),.SO(N494));
  HADDX1 desc286(.A0(N463),.B0(N462),.C1(\add_90_I23_L14036_C129/carry[2] ),.SO(N474));
  HADDX1 desc287(.A0(N464),.B0(\add_90_I23_L14036_C129/carry[2] ),.C1(\add_90_I23_L14036_C129/carry[3] ),.SO(N475));
  HADDX1 desc288(.A0(N465),.B0(\add_90_I23_L14036_C129/carry[3] ),.C1(\add_90_I23_L14036_C129/carry[4] ),.SO(N476));
  HADDX1 desc289(.A0(N466),.B0(\add_90_I23_L14036_C129/carry[4] ),.C1(\add_90_I23_L14036_C129/carry[5] ),.SO(N477));
  HADDX1 desc290(.A0(N446),.B0(N445),.C1(\add_90_I22_L14036_C129/carry[2] ),.SO(N457));
  HADDX1 desc291(.A0(N447),.B0(\add_90_I22_L14036_C129/carry[2] ),.C1(\add_90_I22_L14036_C129/carry[3] ),.SO(N458));
  HADDX1 desc292(.A0(N448),.B0(\add_90_I22_L14036_C129/carry[3] ),.C1(\add_90_I22_L14036_C129/carry[4] ),.SO(N459));
  HADDX1 desc293(.A0(N449),.B0(\add_90_I22_L14036_C129/carry[4] ),.C1(\add_90_I22_L14036_C129/carry[5] ),.SO(N460));
  HADDX1 desc294(.A0(N429),.B0(N428),.C1(\add_90_I21_L14036_C129/carry[2] ),.SO(N440));
  HADDX1 desc295(.A0(N430),.B0(\add_90_I21_L14036_C129/carry[2] ),.C1(\add_90_I21_L14036_C129/carry[3] ),.SO(N441));
  HADDX1 desc296(.A0(N431),.B0(\add_90_I21_L14036_C129/carry[3] ),.C1(\add_90_I21_L14036_C129/carry[4] ),.SO(N442));
  HADDX1 desc297(.A0(N432),.B0(\add_90_I21_L14036_C129/carry[4] ),.C1(\add_90_I21_L14036_C129/carry[5] ),.SO(N443));
  HADDX1 desc298(.A0(N412),.B0(N411),.C1(\add_90_I20_L14036_C129/carry[2] ),.SO(N423));
  HADDX1 desc299(.A0(N413),.B0(\add_90_I20_L14036_C129/carry[2] ),.C1(\add_90_I20_L14036_C129/carry[3] ),.SO(N424));
  HADDX1 desc300(.A0(N414),.B0(\add_90_I20_L14036_C129/carry[3] ),.C1(\add_90_I20_L14036_C129/carry[4] ),.SO(N425));
  HADDX1 desc301(.A0(N415),.B0(\add_90_I20_L14036_C129/carry[4] ),.C1(\add_90_I20_L14036_C129/carry[5] ),.SO(N426));
  HADDX1 desc302(.A0(N395),.B0(N394),.C1(\add_90_I19_L14036_C129/carry[2] ),.SO(N406));
  HADDX1 desc303(.A0(N396),.B0(\add_90_I19_L14036_C129/carry[2] ),.C1(\add_90_I19_L14036_C129/carry[3] ),.SO(N407));
  HADDX1 desc304(.A0(N397),.B0(\add_90_I19_L14036_C129/carry[3] ),.C1(\add_90_I19_L14036_C129/carry[4] ),.SO(N408));
  HADDX1 desc305(.A0(N398),.B0(\add_90_I19_L14036_C129/carry[4] ),.C1(\add_90_I19_L14036_C129/carry[5] ),.SO(N409));
  HADDX1 desc306(.A0(N378),.B0(N377),.C1(\add_90_I18_L14036_C129/carry[2] ),.SO(N389));
  HADDX1 desc307(.A0(N379),.B0(\add_90_I18_L14036_C129/carry[2] ),.C1(\add_90_I18_L14036_C129/carry[3] ),.SO(N390));
  HADDX1 desc308(.A0(N380),.B0(\add_90_I18_L14036_C129/carry[3] ),.C1(\add_90_I18_L14036_C129/carry[4] ),.SO(N391));
  HADDX1 desc309(.A0(N381),.B0(\add_90_I18_L14036_C129/carry[4] ),.C1(\add_90_I18_L14036_C129/carry[5] ),.SO(N392));
  HADDX1 desc310(.A0(N361),.B0(N360),.C1(\add_90_I17_L14036_C129/carry[2] ),.SO(N372));
  HADDX1 desc311(.A0(N362),.B0(\add_90_I17_L14036_C129/carry[2] ),.C1(\add_90_I17_L14036_C129/carry[3] ),.SO(N373));
  HADDX1 desc312(.A0(N363),.B0(\add_90_I17_L14036_C129/carry[3] ),.C1(\add_90_I17_L14036_C129/carry[4] ),.SO(N374));
  HADDX1 desc313(.A0(N364),.B0(\add_90_I17_L14036_C129/carry[4] ),.C1(\add_90_I17_L14036_C129/carry[5] ),.SO(N375));
  HADDX1 desc314(.A0(N344),.B0(N343),.C1(\add_90_I16_L14036_C129/carry[2] ),.SO(N355));
  HADDX1 desc315(.A0(N345),.B0(\add_90_I16_L14036_C129/carry[2] ),.C1(\add_90_I16_L14036_C129/carry[3] ),.SO(N356));
  HADDX1 desc316(.A0(N346),.B0(\add_90_I16_L14036_C129/carry[3] ),.C1(\add_90_I16_L14036_C129/carry[4] ),.SO(N357));
  HADDX1 desc317(.A0(N347),.B0(\add_90_I16_L14036_C129/carry[4] ),.C1(\add_90_I16_L14036_C129/carry[5] ),.SO(N358));
  HADDX1 desc318(.A0(N327),.B0(N326),.C1(\add_90_I15_L14036_C129/carry[2] ),.SO(N338));
  HADDX1 desc319(.A0(N328),.B0(\add_90_I15_L14036_C129/carry[2] ),.C1(\add_90_I15_L14036_C129/carry[3] ),.SO(N339));
  HADDX1 desc320(.A0(N329),.B0(\add_90_I15_L14036_C129/carry[3] ),.C1(\add_90_I15_L14036_C129/carry[4] ),.SO(N340));
  HADDX1 desc321(.A0(N330),.B0(\add_90_I15_L14036_C129/carry[4] ),.C1(\add_90_I15_L14036_C129/carry[5] ),.SO(N341));
  HADDX1 desc322(.A0(N310),.B0(N309),.C1(\add_90_I14_L14036_C129/carry[2] ),.SO(N321));
  HADDX1 desc323(.A0(N311),.B0(\add_90_I14_L14036_C129/carry[2] ),.C1(\add_90_I14_L14036_C129/carry[3] ),.SO(N322));
  HADDX1 desc324(.A0(N312),.B0(\add_90_I14_L14036_C129/carry[3] ),.C1(\add_90_I14_L14036_C129/carry[4] ),.SO(N323));
  HADDX1 desc325(.A0(N313),.B0(\add_90_I14_L14036_C129/carry[4] ),.C1(\add_90_I14_L14036_C129/carry[5] ),.SO(N324));
  HADDX1 desc326(.A0(N293),.B0(N292),.C1(\add_90_I13_L14036_C129/carry[2] ),.SO(N304));
  HADDX1 desc327(.A0(N294),.B0(\add_90_I13_L14036_C129/carry[2] ),.C1(\add_90_I13_L14036_C129/carry[3] ),.SO(N305));
  HADDX1 desc328(.A0(N295),.B0(\add_90_I13_L14036_C129/carry[3] ),.C1(\add_90_I13_L14036_C129/carry[4] ),.SO(N306));
  HADDX1 desc329(.A0(N296),.B0(\add_90_I13_L14036_C129/carry[4] ),.C1(\add_90_I13_L14036_C129/carry[5] ),.SO(N307));
  HADDX1 desc330(.A0(N276),.B0(N275),.C1(\add_90_I12_L14036_C129/carry[2] ),.SO(N287));
  HADDX1 desc331(.A0(N277),.B0(\add_90_I12_L14036_C129/carry[2] ),.C1(\add_90_I12_L14036_C129/carry[3] ),.SO(N288));
  HADDX1 desc332(.A0(N278),.B0(\add_90_I12_L14036_C129/carry[3] ),.C1(\add_90_I12_L14036_C129/carry[4] ),.SO(N289));
  HADDX1 desc333(.A0(N279),.B0(\add_90_I12_L14036_C129/carry[4] ),.C1(\add_90_I12_L14036_C129/carry[5] ),.SO(N290));
  HADDX1 desc334(.A0(N259),.B0(N258),.C1(\add_90_I11_L14036_C129/carry[2] ),.SO(N270));
  HADDX1 desc335(.A0(N260),.B0(\add_90_I11_L14036_C129/carry[2] ),.C1(\add_90_I11_L14036_C129/carry[3] ),.SO(N271));
  HADDX1 desc336(.A0(N261),.B0(\add_90_I11_L14036_C129/carry[3] ),.C1(\add_90_I11_L14036_C129/carry[4] ),.SO(N272));
  HADDX1 desc337(.A0(N262),.B0(\add_90_I11_L14036_C129/carry[4] ),.C1(\add_90_I11_L14036_C129/carry[5] ),.SO(N273));
  HADDX1 desc338(.A0(N242),.B0(N241),.C1(\add_90_I10_L14036_C129/carry[2] ),.SO(N253));
  HADDX1 desc339(.A0(N243),.B0(\add_90_I10_L14036_C129/carry[2] ),.C1(\add_90_I10_L14036_C129/carry[3] ),.SO(N254));
  HADDX1 desc340(.A0(N244),.B0(\add_90_I10_L14036_C129/carry[3] ),.C1(\add_90_I10_L14036_C129/carry[4] ),.SO(N255));
  HADDX1 desc341(.A0(N245),.B0(\add_90_I10_L14036_C129/carry[4] ),.C1(\add_90_I10_L14036_C129/carry[5] ),.SO(N256));
  HADDX1 desc342(.A0(N225),.B0(N224),.C1(\add_90_I9_L14036_C129/carry[2] ),.SO(N236));
  HADDX1 desc343(.A0(N226),.B0(\add_90_I9_L14036_C129/carry[2] ),.C1(\add_90_I9_L14036_C129/carry[3] ),.SO(N237));
  HADDX1 desc344(.A0(N227),.B0(\add_90_I9_L14036_C129/carry[3] ),.C1(\add_90_I9_L14036_C129/carry[4] ),.SO(N238));
  HADDX1 desc345(.A0(N228),.B0(\add_90_I9_L14036_C129/carry[4] ),.C1(\add_90_I9_L14036_C129/carry[5] ),.SO(N239));
  HADDX1 desc346(.A0(N208),.B0(N207),.C1(\add_90_I8_L14036_C129/carry[2] ),.SO(N219));
  HADDX1 desc347(.A0(N209),.B0(\add_90_I8_L14036_C129/carry[2] ),.C1(\add_90_I8_L14036_C129/carry[3] ),.SO(N220));
  HADDX1 desc348(.A0(N210),.B0(\add_90_I8_L14036_C129/carry[3] ),.C1(\add_90_I8_L14036_C129/carry[4] ),.SO(N221));
  HADDX1 desc349(.A0(N211),.B0(\add_90_I8_L14036_C129/carry[4] ),.C1(\add_90_I8_L14036_C129/carry[5] ),.SO(N222));
  HADDX1 desc350(.A0(N191),.B0(N190),.C1(\add_90_I7_L14036_C129/carry[2] ),.SO(N202));
  HADDX1 desc351(.A0(N192),.B0(\add_90_I7_L14036_C129/carry[2] ),.C1(\add_90_I7_L14036_C129/carry[3] ),.SO(N203));
  HADDX1 desc352(.A0(N193),.B0(\add_90_I7_L14036_C129/carry[3] ),.C1(\add_90_I7_L14036_C129/carry[4] ),.SO(N204));
  HADDX1 desc353(.A0(N194),.B0(\add_90_I7_L14036_C129/carry[4] ),.C1(N206),.SO(N205));
  HADDX1 desc354(.A0(N175),.B0(N174),.C1(\add_90_I6_L14036_C129/carry[2] ),.SO(N185));
  HADDX1 desc355(.A0(N176),.B0(\add_90_I6_L14036_C129/carry[2] ),.C1(\add_90_I6_L14036_C129/carry[3] ),.SO(N186));
  HADDX1 desc356(.A0(N177),.B0(\add_90_I6_L14036_C129/carry[3] ),.C1(N188),.SO(N187));
  HADDX1 desc357(.A0(\add_90_I5_L14036_C129/A[1] ),.B0(N160),.C1(\add_90_I5_L14036_C129/carry[2] ),.SO(N170));
  HADDX1 desc358(.A0(N162),.B0(\add_90_I5_L14036_C129/carry[2] ),.C1(N172),.SO(N171));
  FADDX1 desc359(.A(\sub_0_root_add_0_root_sub_132/A[1] ),.B(n35),.CI(\sub_0_root_add_0_root_sub_132/carry[1] ),.CO(\sub_0_root_add_0_root_sub_132/carry[2] ),.S(s_exp10[1:1]));
  FADDX1 desc360(.A(\sub_0_root_add_0_root_sub_132/A[2] ),.B(n149),.CI(\sub_0_root_add_0_root_sub_132/carry[2] ),.CO(\sub_0_root_add_0_root_sub_132/carry[3] ),.S(s_exp10[2:2]));
  FADDX1 desc361(.A(\sub_0_root_add_0_root_sub_132/A[3] ),.B(n34),.CI(\sub_0_root_add_0_root_sub_132/carry[3] ),.CO(\sub_0_root_add_0_root_sub_132/carry[4] ),.S(s_exp10[3:3]));
  FADDX1 desc362(.A(\sub_0_root_add_0_root_sub_132/A[4] ),.B(n37),.CI(\sub_0_root_add_0_root_sub_132/carry[4] ),.CO(\sub_0_root_add_0_root_sub_132/carry[5] ),.S(s_exp10[4:4]));
  FADDX1 desc363(.A(\sub_0_root_add_0_root_sub_132/A[5] ),.B(n38),.CI(\sub_0_root_add_0_root_sub_132/carry[5] ),.CO(\sub_0_root_add_0_root_sub_132/carry[6] ),.S(s_exp10[5:5]));
  NBUFFX2 U4(.INP(s_shl1[5:5]),.Z(n28));
  NOR2X0 U5(.IN1(n283),.IN2(n11),.QN(n153));
  NAND2X0 U6(.IN1(n257),.IN2(n302),.QN(n258));
  NAND2X0 U7(.IN1(n102),.IN2(n104),.QN(n259));
  NAND2X0 U8(.IN1(n222),.IN2(n103),.QN(n221));
  NAND2X0 U10(.IN1(n157),.IN2(n100),.QN(n220));
  INVX0 U11(.INP(n382),.ZN(n77));
  INVX0 U12(.INP(n389),.ZN(n78));
  INVX0 U13(.INP(n396),.ZN(n79));
  NOR2X0 U14(.IN1(n48),.IN2(s_exp10[8:8]),.QN(n155));
  INVX0 U15(.INP(n153),.ZN(n48));
  INVX0 U16(.INP(n237),.ZN(\add_90_I5_L14036_C129/A[1] ));
  INVX0 U17(.INP(n149),.ZN(\sub_0_root_add_0_root_sub_132/B[2] ));
  INVX0 U18(.INP(n150),.ZN(\sub_0_root_add_0_root_sub_132/B[5] ));
  AND2X1 U19(.IN1(n148),.IN2(n60),.Q(n21));
  AND2X1 U20(.IN1(n148),.IN2(n60),.Q(n114));
  INVX0 U21(.INP(n124),.ZN(n57));
  INVX0 U22(.INP(n277),.ZN(n318));
  INVX0 U23(.INP(n278),.ZN(n311));
  NAND2X1 U24(.IN1(n311),.IN2(n178),.QN(n176));
  INVX0 U25(.INP(n221),.ZN(n102));
  INVX0 U26(.INP(n117),.ZN(n325));
  INVX0 U27(.INP(n220),.ZN(n86));
  INVX0 U28(.INP(n411),.ZN(n80));
  INVX0 U29(.INP(n375),.ZN(n76));
  INVX0 U30(.INP(n376),.ZN(n65));
  INVX0 U31(.INP(n384),.ZN(n66));
  INVX0 U32(.INP(n391),.ZN(n67));
  INVX0 U33(.INP(n398),.ZN(n68));
  INVX0 U34(.INP(n405),.ZN(n69));
  INVX0 U36(.INP(n364),.ZN(n63));
  INVX0 U37(.INP(n370),.ZN(n64));
  INVX0 U38(.INP(n369),.ZN(n75));
  INVX0 U39(.INP(n414),.ZN(n74));
  INVX0 U40(.INP(n345),.ZN(n81));
  INVX0 U41(.INP(n425),.ZN(n72));
  INVX0 U42(.INP(n362),.ZN(n83));
  INVX0 U43(.INP(n355),.ZN(n82));
  NOR2X0 U44(.IN1(n334),.IN2(n24),.QN(n414));
  NOR2X0 U45(.IN1(n365),.IN2(n24),.QN(n423));
  NOR2X0 U46(.IN1(\sub_0_root_add_0_root_sub_132/A[8] ),.IN2(\sub_0_root_add_0_root_sub_132/carry[8] ),.QN(n11));
  INVX0 U47(.INP(N396),.ZN(n95));
  INVX0 U48(.INP(N447),.ZN(n92));
  NOR2X0 U49(.IN1(n231),.IN2(n232),.QN(n230));
  INVX0 U50(.INP(N397),.ZN(n91));
  INVX0 U51(.INP(N448),.ZN(n88));
  NOR2X0 U52(.IN1(n216),.IN2(n217),.QN(n215));
  INVX0 U53(.INP(N399),.ZN(n52));
  INVX0 U54(.INP(N450),.ZN(n49));
  NOR2X0 U55(.IN1(n179),.IN2(n180),.QN(n177));
  NAND2X0 U56(.IN1(n157),.IN2(n158),.QN(n150));
  NOR2X0 U57(.IN1(n247),.IN2(n248),.QN(n246));
  INVX0 U58(.INP(N445),.ZN(N456));
  INVX0 U59(.INP(N241),.ZN(N252));
  INVX0 U60(.INP(N343),.ZN(N354));
  INVX0 U61(.INP(n19),.ZN(n304));
  INVX0 U62(.INP(N398),.ZN(n56));
  INVX0 U63(.INP(N449),.ZN(n53));
  NOR2X0 U64(.IN1(n203),.IN2(n204),.QN(n202));
  NOR2X0 U65(.IN1(n272),.IN2(n273),.QN(n271));
  INVX0 U66(.INP(N530),.ZN(N541));
  AND2X1 U67(.IN1(N206),.IN2(n126),.Q(n12));
  INVX0 U68(.INP(s_zeros[0:0]),.ZN(n36));
  AND2X1 U69(.IN1(n148),.IN2(s_fracto28_rnd[27:27]),.Q(n113));
  INVX0 U70(.INP(n17),.ZN(n310));
  OR2X1 U71(.IN1(n118),.IN2(n13),.Q(s_output_o[22:22]));
  AND3X1 U72(.IN1(n127),.IN2(n125),.IN3(n124),.Q(n13));
  INVX0 U73(.INP(N430),.ZN(n93));
  INVX0 U74(.INP(N429),.ZN(n97));
  INVX0 U75(.INP(N431),.ZN(n89));
  INVX0 U76(.INP(N446),.ZN(n96));
  INVX0 U77(.INP(n16),.ZN(n317));
  INVX0 U78(.INP(s_fracto28_rnd[27:27]),.ZN(n60));
  NAND2X1 U79(.IN1(n295),.IN2(n296),.QN(n152));
  INVX0 U80(.INP(N413),.ZN(n94));
  INVX0 U81(.INP(N412),.ZN(n98));
  INVX0 U82(.INP(N414),.ZN(n90));
  INVX0 U83(.INP(N415),.ZN(n55));
  INVX0 U84(.INP(N416),.ZN(n51));
  INVX0 U85(.INP(N432),.ZN(n54));
  INVX0 U86(.INP(N433),.ZN(n50));
  INVX0 U87(.INP(N395),.ZN(n99));
  NOR2X0 U88(.IN1(n275),.IN2(n276),.QN(n183));
  NOR2X0 U89(.IN1(n266),.IN2(n170),.QN(n169));
  NOR2X0 U90(.IN1(n274),.IN2(n16),.QN(n181));
  NAND2X1 U91(.IN1(n311),.IN2(n316),.QN(n178));
  NOR2X0 U92(.IN1(n279),.IN2(n17),.QN(n185));
  NOR2X0 U93(.IN1(n264),.IN2(n265),.QN(n189));
  NAND2X1 U94(.IN1(n279),.IN2(n313),.QN(n280));
  NAND2X1 U95(.IN1(n274),.IN2(n320),.QN(n275));
  NAND2X1 U96(.IN1(n263),.IN2(n306),.QN(n264));
  NAND2X1 U97(.IN1(n265),.IN2(n308),.QN(n266));
  NAND2X1 U98(.IN1(n279),.IN2(n280),.QN(n175));
  NAND2X1 U99(.IN1(n281),.IN2(n278),.QN(n187));
  NAND2X1 U100(.IN1(n281),.IN2(n315),.QN(n278));
  NOR2X0 U101(.IN1(n258),.IN2(n160),.QN(n159));
  NOR2X0 U102(.IN1(n259),.IN2(n257),.QN(n164));
  NOR2X0 U103(.IN1(n263),.IN2(n19),.QN(n188));
  NAND2X1 U104(.IN1(n129),.IN2(n130),.QN(n117));
  INVX0 U105(.INP(n160),.ZN(n101));
  NAND2X0 U106(.IN1(n193),.IN2(N190),.QN(n254));
  NOR2X0 U107(.IN1(n32),.IN2(n87),.QN(N998));
  NOR2X0 U108(.IN1(n444),.IN2(n28),.QN(N1026));
  INVX0 U109(.INP(n413),.ZN(n70));
  INVX0 U110(.INP(n422),.ZN(n71));
  INVX0 U111(.INP(n433),.ZN(n73));
  INVX0 U112(.INP(n442),.ZN(n61));
  NAND2X1 U113(.IN1(n406),.IN2(n6),.QN(n450));
  NAND2X1 U114(.IN1(n414),.IN2(n6),.QN(n357));
  INVX0 U115(.INP(N1093),.ZN(n59));
  NAND2X1 U116(.IN1(N1095),.IN2(N1094),.QN(n301));
  NAND2X1 U117(.IN1(n423),.IN2(n6),.QN(n379));
  NAND2X1 U118(.IN1(n341),.IN2(n7),.QN(n365));
  INVX0 U119(.INP(n333),.ZN(n84));
  INVX0 U120(.INP(n43),.ZN(n47));
  INVX0 U121(.INP(n41),.ZN(n45));
  INVX0 U122(.INP(n42),.ZN(n46));
  NAND2X1 U123(.IN1(n350),.IN2(n9),.QN(n377));
  INVX0 U124(.INP(n14),.ZN(n58));
  INVX0 U125(.INP(n9),.ZN(n24));
  INVX0 U126(.INP(n8),.ZN(n22));
  INVX0 U127(.INP(n7),.ZN(n23));
  INVX0 U128(.INP(s_zeros[4:4]),.ZN(n37));
  INVX0 U129(.INP(s_zeros[3:3]),.ZN(n34));
  INVX0 U130(.INP(s_zeros[1:1]),.ZN(n35));
  NOR2X0 U131(.IN1(n288),.IN2(fract_28_i[23:23]),.QN(n286));
  NAND2X0 U132(.IN1(n193),.IN2(N191),.QN(n235));
  NOR2X0 U133(.IN1(fract_28_i[25:25]),.IN2(fract_28_i[26:26]),.QN(n282));
  INVX0 U134(.INP(\sub_0_root_add_0_root_sub_132/B[5] ),.ZN(n38));
  INVX0 U135(.INP(exp_i[0:0]),.ZN(N920));
  NBUFFX2 U136(.INP(fract_28_i[17:17]),.Z(n20));
  NBUFFX2 U137(.INP(fract_28_i[17:17]),.Z(n19));
  INVX0 U138(.INP(N174),.ZN(N184));
  INVX0 U139(.INP(N377),.ZN(N388));
  INVX0 U140(.INP(N394),.ZN(N405));
  INVX0 U141(.INP(N411),.ZN(N422));
  INVX0 U142(.INP(N428),.ZN(N439));
  INVX0 U169(.INP(N496),.ZN(N507));
  INVX0 U206(.INP(N479),.ZN(N490));
  INVX0 U207(.INP(N207),.ZN(N218));
  INVX0 U432(.INP(N326),.ZN(N337));
  INVX0 U438(.INP(N190),.ZN(N201));
  INVX0 U439(.INP(N258),.ZN(N269));
  INVX0 U444(.INP(N224),.ZN(N235));
  INVX0 U449(.INP(N309),.ZN(N320));
  INVX0 U497(.INP(N292),.ZN(N303));
  INVX0 U498(.INP(N275),.ZN(N286));
  INVX0 U499(.INP(N513),.ZN(N524));
  INVX0 U500(.INP(fract_28_i[24:24]),.ZN(n100));
  NOR2X0 U501(.IN1(fract_28_i[27:27]),.IN2(fract_28_i[26:26]),.QN(n252));
  INVX0 U502(.INP(N160),.ZN(N169));
  INVX0 U503(.INP(N462),.ZN(N473));
  INVX0 U504(.INP(N360),.ZN(N371));
  NBUFFX2 U505(.INP(fract_28_i[11:11]),.Z(n18));
  NBUFFX2 U506(.INP(fract_28_i[11:11]),.Z(n17));
  INVX0 U507(.INP(fract_28_i[19:19]),.ZN(n302));
  INVX0 U508(.INP(fract_28_i[20:20]),.ZN(n126));
  INVX0 U509(.INP(fract_28_i[21:21]),.ZN(n104));
  INVX0 U510(.INP(fract_28_i[18:18]),.ZN(n303));
  INVX0 U511(.INP(fract_28_i[22:22]),.ZN(n103));
  NOR2X0 U512(.IN1(n323),.IN2(n87),.QN(n112));
  NBUFFX2 U513(.INP(fract_28_i[5:5]),.Z(n16));
  INVX0 U514(.INP(fract_28_i[15:15]),.ZN(n306));
  INVX0 U515(.INP(fract_28_i[13:13]),.ZN(n308));
  INVX0 U516(.INP(fract_28_i[27:27]),.ZN(n87));
  INVX0 U517(.INP(fract_28_i[14:14]),.ZN(n307));
  INVX0 U518(.INP(fract_28_i[12:12]),.ZN(n309));
  INVX0 U519(.INP(fract_28_i[16:16]),.ZN(n305));
  INVX0 U520(.INP(fract_28_i[10:10]),.ZN(n312));
  NAND2X1 U521(.IN1(n105),.IN2(n106),.QN(s_roundup));
  INVX0 U522(.INP(rmode_i[1:1]),.ZN(n326));
  INVX0 U523(.INP(fract_28_i[0:0]),.ZN(n323));
  INVX0 U524(.INP(rmode_i[0:0]),.ZN(n327));
  NAND2X1 U525(.IN1(n39),.IN2(n107),.QN(n111));
  NAND2X0 U526(.IN1(rmode_i[1:1]),.IN2(n327),.QN(n110));
  NOR2X0 U527(.IN1(fract_28_i[10:10]),.IN2(n17),.QN(n279));
  NOR2X0 U528(.IN1(n266),.IN2(fract_28_i[12:12]),.QN(n170));
  NOR2X0 U529(.IN1(n280),.IN2(fract_28_i[8:8]),.QN(n281));
  NOR2X0 U530(.IN1(fract_28_i[4:4]),.IN2(n16),.QN(n274));
  NOR2X0 U531(.IN1(fract_28_i[16:16]),.IN2(n19),.QN(n263));
  NOR2X0 U532(.IN1(n264),.IN2(fract_28_i[14:14]),.QN(n265));
  INVX0 U533(.INP(fract_28_i[9:9]),.ZN(n313));
  INVX0 U534(.INP(fract_28_i[7:7]),.ZN(n315));
  NOR2X0 U535(.IN1(n275),.IN2(fract_28_i[2:2]),.QN(n276));
  INVX0 U536(.INP(fract_28_i[8:8]),.ZN(n314));
  NOR2X0 U537(.IN1(n292),.IN2(n293),.QN(n129));
  NOR2X0 U538(.IN1(n258),.IN2(fract_28_i[18:18]),.QN(n160));
  NOR2X0 U539(.IN1(n259),.IN2(fract_28_i[20:20]),.QN(n257));
  INVX0 U540(.INP(fract_28_i[3:3]),.ZN(n320));
  INVX0 U541(.INP(fract_28_i[6:6]),.ZN(n316));
  INVX0 U542(.INP(fract_28_i[4:4]),.ZN(n319));
  NOR2X0 U543(.IN1(fract_28_i[23:23]),.IN2(fract_28_i[24:24]),.QN(n222));
  INVX0 U544(.INP(n115),.ZN(n324));
  NAND2X1 U545(.IN1(n118),.IN2(n119),.QN(n115));
  INVX0 U546(.INP(fract_28_i[1:1]),.ZN(n322));
  INVX0 U547(.INP(fract_28_i[2:2]),.ZN(n321));
  NOR2X0 U548(.IN1(n28),.IN2(n359),.QN(N1015));
  NOR2X0 U549(.IN1(n28),.IN2(n366),.QN(N1016));
  NOR2X0 U550(.IN1(n28),.IN2(n372),.QN(N1017));
  NOR2X0 U551(.IN1(n28),.IN2(n378),.QN(N1018));
  NOR2X0 U552(.IN1(n28),.IN2(n386),.QN(N1019));
  NOR2X0 U553(.IN1(n28),.IN2(n393),.QN(N1020));
  NOR2X0 U554(.IN1(n28),.IN2(n400),.QN(N1021));
  NOR2X0 U555(.IN1(n28),.IN2(n407),.QN(N1022));
  NOR2X0 U556(.IN1(n28),.IN2(n416),.QN(N1023));
  NOR2X0 U557(.IN1(n28),.IN2(n435),.QN(N1025));
  NOR2X0 U558(.IN1(n28),.IN2(n426),.QN(N1024));
  INVX0 U559(.INP(n352),.ZN(n62));
  NOR2X0 U560(.IN1(n290),.IN2(n291),.QN(n121));
  NAND2X1 U561(.IN1(fract_28_i[0:0]),.IN2(n8),.QN(n329));
  NOR2X0 U562(.IN1(s_expo9_1[7:7]),.IN2(\sub_172_aco/carry[7] ),.QN(n14));
  OR2X1 U563(.IN1(s_fracto28_1[27:27]),.IN2(s_fracto28_1[26:26]),.Q(n15));
  INVX0 U564(.INP(n328),.ZN(n85));
  INVX0 U565(.INP(\s_shr1[0] ),.ZN(n33));
  NBUFFX2 U566(.INP(s_shl1[4:4]),.Z(n27));
  NBUFFX2 U567(.INP(s_shl1[4:4]),.Z(n26));
  NBUFFX2 U568(.INP(s_shl1[5:5]),.Z(n29));
  INVX0 U569(.INP(n6),.ZN(n25));
  INVX0 U570(.INP(n33),.ZN(n32));
  XNOR2X1 U571(.IN1(\sub_172_aco/carry[7] ),.IN2(s_expo9_1[7:7]),.Q(s_expo9_2[7:7]));
  OR2X1 U572(.IN1(s_expo9_1[6:6]),.IN2(\sub_172_aco/carry[6] ),.Q(\sub_172_aco/carry[7] ));
  XNOR2X1 U573(.IN1(\sub_172_aco/carry[6] ),.IN2(s_expo9_1[6:6]),.Q(s_expo9_2[6:6]));
  OR2X1 U574(.IN1(s_expo9_1[5:5]),.IN2(\sub_172_aco/carry[5] ),.Q(\sub_172_aco/carry[6] ));
  XNOR2X1 U575(.IN1(\sub_172_aco/carry[5] ),.IN2(s_expo9_1[5:5]),.Q(s_expo9_2[5:5]));
  OR2X1 U576(.IN1(s_expo9_1[4:4]),.IN2(\sub_172_aco/carry[4] ),.Q(\sub_172_aco/carry[5] ));
  XNOR2X1 U577(.IN1(\sub_172_aco/carry[4] ),.IN2(s_expo9_1[4:4]),.Q(s_expo9_2[4:4]));
  OR2X1 U578(.IN1(s_expo9_1[3:3]),.IN2(\sub_172_aco/carry[3] ),.Q(\sub_172_aco/carry[4] ));
  XNOR2X1 U579(.IN1(\sub_172_aco/carry[3] ),.IN2(s_expo9_1[3:3]),.Q(s_expo9_2[3:3]));
  OR2X1 U580(.IN1(s_expo9_1[2:2]),.IN2(\sub_172_aco/carry[2] ),.Q(\sub_172_aco/carry[3] ));
  XNOR2X1 U581(.IN1(\sub_172_aco/carry[2] ),.IN2(s_expo9_1[2:2]),.Q(s_expo9_2[2:2]));
  OR2X1 U582(.IN1(s_expo9_1[1:1]),.IN2(\sub_172_aco/carry[1] ),.Q(\sub_172_aco/carry[2] ));
  XNOR2X1 U583(.IN1(\sub_172_aco/carry[1] ),.IN2(s_expo9_1[1:1]),.Q(s_expo9_2[1:1]));
  OR2X1 U584(.IN1(s_expo9_1[0:0]),.IN2(n15),.Q(\sub_172_aco/carry[1] ));
  XNOR2X1 U585(.IN1(n15),.IN2(s_expo9_1[0:0]),.Q(s_expo9_2[0:0]));
  XNOR2X1 U586(.IN1(\sub_0_root_add_0_root_sub_132/carry[8] ),.IN2(\sub_0_root_add_0_root_sub_132/A[8] ),.Q(s_exp10[8:8]));
  OR2X1 U587(.IN1(\sub_0_root_add_0_root_sub_132/A[7] ),.IN2(\sub_0_root_add_0_root_sub_132/carry[7] ),.Q(\sub_0_root_add_0_root_sub_132/carry[8] ));
  XNOR2X1 U588(.IN1(\sub_0_root_add_0_root_sub_132/carry[7] ),.IN2(\sub_0_root_add_0_root_sub_132/A[7] ),.Q(s_exp10[7:7]));
  OR2X1 U589(.IN1(\sub_0_root_add_0_root_sub_132/A[6] ),.IN2(\sub_0_root_add_0_root_sub_132/carry[6] ),.Q(\sub_0_root_add_0_root_sub_132/carry[7] ));
  XNOR2X1 U590(.IN1(\sub_0_root_add_0_root_sub_132/carry[6] ),.IN2(\sub_0_root_add_0_root_sub_132/A[6] ),.Q(s_exp10[6:6]));
  OR2X1 U591(.IN1(\sub_0_root_add_0_root_sub_132/A[0] ),.IN2(n36),.Q(\sub_0_root_add_0_root_sub_132/carry[1] ));
  XNOR2X1 U592(.IN1(n36),.IN2(\sub_0_root_add_0_root_sub_132/A[0] ),.Q(s_exp10[0:0]));
  AND2X1 U593(.IN1(\add_1_root_add_0_root_sub_132/carry[7] ),.IN2(exp_i[7:7]),.Q(\sub_0_root_add_0_root_sub_132/A[8] ));
  XOR2X1 U594(.IN1(exp_i[7:7]),.IN2(\add_1_root_add_0_root_sub_132/carry[7] ),.Q(\sub_0_root_add_0_root_sub_132/A[7] ));
  AND2X1 U595(.IN1(exp_i[6:6]),.IN2(\add_1_root_add_0_root_sub_132/carry[6] ),.Q(\add_1_root_add_0_root_sub_132/carry[7] ));
  XOR2X1 U596(.IN1(exp_i[6:6]),.IN2(\add_1_root_add_0_root_sub_132/carry[6] ),.Q(\sub_0_root_add_0_root_sub_132/A[6] ));
  AND2X1 U597(.IN1(exp_i[5:5]),.IN2(\add_1_root_add_0_root_sub_132/carry[5] ),.Q(\add_1_root_add_0_root_sub_132/carry[6] ));
  XOR2X1 U598(.IN1(exp_i[5:5]),.IN2(\add_1_root_add_0_root_sub_132/carry[5] ),.Q(\sub_0_root_add_0_root_sub_132/A[5] ));
  AND2X1 U599(.IN1(exp_i[4:4]),.IN2(\add_1_root_add_0_root_sub_132/carry[4] ),.Q(\add_1_root_add_0_root_sub_132/carry[5] ));
  XOR2X1 U600(.IN1(exp_i[4:4]),.IN2(\add_1_root_add_0_root_sub_132/carry[4] ),.Q(\sub_0_root_add_0_root_sub_132/A[4] ));
  AND2X1 U601(.IN1(exp_i[3:3]),.IN2(\add_1_root_add_0_root_sub_132/carry[3] ),.Q(\add_1_root_add_0_root_sub_132/carry[4] ));
  XOR2X1 U602(.IN1(exp_i[3:3]),.IN2(\add_1_root_add_0_root_sub_132/carry[3] ),.Q(\sub_0_root_add_0_root_sub_132/A[3] ));
  AND2X1 U603(.IN1(exp_i[2:2]),.IN2(\add_1_root_add_0_root_sub_132/carry[2] ),.Q(\add_1_root_add_0_root_sub_132/carry[3] ));
  XOR2X1 U604(.IN1(exp_i[2:2]),.IN2(\add_1_root_add_0_root_sub_132/carry[2] ),.Q(\sub_0_root_add_0_root_sub_132/A[2] ));
  AND2X1 U605(.IN1(exp_i[1:1]),.IN2(\add_1_root_add_0_root_sub_132/carry[1] ),.Q(\add_1_root_add_0_root_sub_132/carry[2] ));
  XOR2X1 U606(.IN1(exp_i[1:1]),.IN2(\add_1_root_add_0_root_sub_132/carry[1] ),.Q(\sub_0_root_add_0_root_sub_132/A[1] ));
  AND2X1 U607(.IN1(fract_28_i[27:27]),.IN2(exp_i[0:0]),.Q(\add_1_root_add_0_root_sub_132/carry[1] ));
  XOR2X1 U608(.IN1(fract_28_i[27:27]),.IN2(exp_i[0:0]),.Q(\sub_0_root_add_0_root_sub_132/A[0] ));
  XOR2X1 U609(.IN1(\add_90_I8_L14036_C129/carry[5] ),.IN2(n12),.Q(N223));
  XOR2X1 U610(.IN1(\add_90_I9_L14036_C129/carry[5] ),.IN2(N229),.Q(N240));
  XOR2X1 U611(.IN1(\add_90_I10_L14036_C129/carry[5] ),.IN2(N246),.Q(N257));
  XOR2X1 U612(.IN1(\add_90_I11_L14036_C129/carry[5] ),.IN2(N263),.Q(N274));
  XOR2X1 U613(.IN1(\add_90_I12_L14036_C129/carry[5] ),.IN2(N280),.Q(N291));
  XOR2X1 U614(.IN1(\add_90_I13_L14036_C129/carry[5] ),.IN2(N297),.Q(N308));
  XOR2X1 U615(.IN1(\add_90_I14_L14036_C129/carry[5] ),.IN2(N314),.Q(N325));
  XOR2X1 U616(.IN1(\add_90_I15_L14036_C129/carry[5] ),.IN2(N331),.Q(N342));
  XOR2X1 U617(.IN1(\add_90_I16_L14036_C129/carry[5] ),.IN2(N348),.Q(N359));
  XOR2X1 U618(.IN1(\add_90_I17_L14036_C129/carry[5] ),.IN2(N365),.Q(N376));
  XOR2X1 U619(.IN1(\add_90_I18_L14036_C129/carry[5] ),.IN2(N382),.Q(N393));
  XOR2X1 U620(.IN1(\add_90_I19_L14036_C129/carry[5] ),.IN2(N399),.Q(N410));
  XOR2X1 U621(.IN1(\add_90_I20_L14036_C129/carry[5] ),.IN2(N416),.Q(N427));
  XOR2X1 U622(.IN1(\add_90_I21_L14036_C129/carry[5] ),.IN2(N433),.Q(N444));
  XOR2X1 U623(.IN1(\add_90_I22_L14036_C129/carry[5] ),.IN2(N450),.Q(N461));
  XOR2X1 U624(.IN1(\add_90_I23_L14036_C129/carry[5] ),.IN2(N467),.Q(N478));
  XOR2X1 U625(.IN1(\add_90_I24_L14036_C129/carry[5] ),.IN2(N484),.Q(N495));
  XOR2X1 U626(.IN1(\add_90_I25_L14036_C129/carry[5] ),.IN2(N501),.Q(N512));
  XOR2X1 U627(.IN1(\add_90_I26_L14036_C129/carry[5] ),.IN2(N518),.Q(N529));
  XOR2X1 U628(.IN1(\add_90_I27_L14036_C129/carry[5] ),.IN2(N535),.Q(N546));
  NOR2X0 U629(.IN1(exp_i[1:1]),.IN2(exp_i[0:0]),.QN(n41));
  AO21X1 U630(.IN1(exp_i[1:1]),.IN2(exp_i[0:0]),.IN3(n41),.Q(N921));
  NOR2X0 U631(.IN1(n45),.IN2(exp_i[2:2]),.QN(n42));
  AO21X1 U632(.IN1(exp_i[2:2]),.IN2(n45),.IN3(n42),.Q(N922));
  NOR2X0 U633(.IN1(n46),.IN2(exp_i[3:3]),.QN(n43));
  AO21X1 U634(.IN1(exp_i[3:3]),.IN2(n46),.IN3(n43),.Q(N923));
  XNOR2X1 U635(.IN1(exp_i[4:4]),.IN2(n47),.Q(N924));
  NOR2X0 U636(.IN1(exp_i[4:4]),.IN2(n47),.QN(n44));
  XOR2X1 U637(.IN1(exp_i[5:5]),.IN2(n44),.Q(N925));
  AND2X1 U638(.IN1(N188),.IN2(n104),.Q(N194));
  MUX21X1 U639(.IN1(fract_28_i[0:0]),.IN2(fract_28_i[1:1]),.S(n32),.Q(N971));
  MUX21X1 U640(.IN1(fract_28_i[10:10]),.IN2(n18),.S(n32),.Q(N981));
  MUX21X1 U641(.IN1(n18),.IN2(fract_28_i[12:12]),.S(n32),.Q(N982));
  MUX21X1 U642(.IN1(fract_28_i[12:12]),.IN2(fract_28_i[13:13]),.S(n32),.Q(N983));
  MUX21X1 U643(.IN1(fract_28_i[13:13]),.IN2(fract_28_i[14:14]),.S(n32),.Q(N984));
  MUX21X1 U644(.IN1(fract_28_i[14:14]),.IN2(fract_28_i[15:15]),.S(n32),.Q(N985));
  MUX21X1 U645(.IN1(fract_28_i[15:15]),.IN2(fract_28_i[16:16]),.S(n32),.Q(N986));
  MUX21X1 U646(.IN1(fract_28_i[16:16]),.IN2(n20),.S(n32),.Q(N987));
  MUX21X1 U647(.IN1(n20),.IN2(fract_28_i[18:18]),.S(n32),.Q(N988));
  MUX21X1 U648(.IN1(fract_28_i[18:18]),.IN2(fract_28_i[19:19]),.S(n32),.Q(N989));
  MUX21X1 U649(.IN1(fract_28_i[19:19]),.IN2(fract_28_i[20:20]),.S(n32),.Q(N990));
  MUX21X1 U650(.IN1(fract_28_i[1:1]),.IN2(fract_28_i[2:2]),.S(n32),.Q(N972));
  MUX21X1 U651(.IN1(fract_28_i[20:20]),.IN2(fract_28_i[21:21]),.S(n32),.Q(N991));
  MUX21X1 U652(.IN1(fract_28_i[21:21]),.IN2(fract_28_i[22:22]),.S(n32),.Q(N992));
  MUX21X1 U653(.IN1(fract_28_i[22:22]),.IN2(fract_28_i[23:23]),.S(n32),.Q(N993));
  MUX21X1 U654(.IN1(fract_28_i[23:23]),.IN2(fract_28_i[24:24]),.S(n32),.Q(N994));
  MUX21X1 U655(.IN1(fract_28_i[24:24]),.IN2(fract_28_i[25:25]),.S(n32),.Q(N995));
  MUX21X1 U656(.IN1(fract_28_i[25:25]),.IN2(fract_28_i[26:26]),.S(\s_shr1[0] ),.Q(N996));
  MUX21X1 U657(.IN1(fract_28_i[26:26]),.IN2(fract_28_i[27:27]),.S(\s_shr1[0] ),.Q(N997));
  MUX21X1 U658(.IN1(fract_28_i[2:2]),.IN2(fract_28_i[3:3]),.S(\s_shr1[0] ),.Q(N973));
  MUX21X1 U659(.IN1(fract_28_i[3:3]),.IN2(fract_28_i[4:4]),.S(\s_shr1[0] ),.Q(N974));
  MUX21X1 U660(.IN1(fract_28_i[4:4]),.IN2(n16),.S(\s_shr1[0] ),.Q(N975));
  MUX21X1 U661(.IN1(n16),.IN2(fract_28_i[6:6]),.S(\s_shr1[0] ),.Q(N976));
  MUX21X1 U662(.IN1(fract_28_i[6:6]),.IN2(fract_28_i[7:7]),.S(\s_shr1[0] ),.Q(N977));
  MUX21X1 U663(.IN1(fract_28_i[7:7]),.IN2(fract_28_i[8:8]),.S(\s_shr1[0] ),.Q(N978));
  MUX21X1 U664(.IN1(fract_28_i[8:8]),.IN2(fract_28_i[9:9]),.S(\s_shr1[0] ),.Q(N979));
  MUX21X1 U665(.IN1(fract_28_i[9:9]),.IN2(fract_28_i[10:10]),.S(\s_shr1[0] ),.Q(N980));
  OR2X1 U666(.IN1(n329),.IN2(n5),.Q(n334));
  NOR3X0 U667(.IN1(n357),.IN2(n28),.IN3(n27),.QN(N999));
  MUX21X1 U668(.IN1(fract_28_i[10:10]),.IN2(fract_28_i[9:9]),.S(n22),.Q(n330));
  MUX21X1 U669(.IN1(fract_28_i[8:8]),.IN2(fract_28_i[7:7]),.S(n22),.Q(n332));
  MUX21X1 U670(.IN1(n330),.IN2(n332),.S(n5),.Q(n344));
  MUX21X1 U671(.IN1(fract_28_i[6:6]),.IN2(n16),.S(n22),.Q(n331));
  MUX21X1 U672(.IN1(fract_28_i[4:4]),.IN2(fract_28_i[3:3]),.S(n22),.Q(n333));
  MUX21X1 U673(.IN1(n331),.IN2(n333),.S(n5),.Q(n345));
  MUX21X1 U674(.IN1(n344),.IN2(n345),.S(n24),.Q(n369));
  MUX21X1 U675(.IN1(fract_28_i[2:2]),.IN2(fract_28_i[1:1]),.S(n22),.Q(n328));
  MUX21X1 U676(.IN1(n85),.IN2(n329),.S(n23),.Q(n346));
  OR2X1 U677(.IN1(n346),.IN2(n3),.Q(n371));
  MUX21X1 U678(.IN1(n75),.IN2(n371),.S(n25),.Q(n434));
  NOR3X0 U679(.IN1(n434),.IN2(n28),.IN3(n27),.QN(N1009));
  MUX21X1 U680(.IN1(n18),.IN2(fract_28_i[10:10]),.S(n22),.Q(n336));
  MUX21X1 U681(.IN1(fract_28_i[9:9]),.IN2(fract_28_i[8:8]),.S(n22),.Q(n338));
  MUX21X1 U682(.IN1(n336),.IN2(n338),.S(n23),.Q(n349));
  MUX21X1 U683(.IN1(fract_28_i[7:7]),.IN2(fract_28_i[6:6]),.S(n22),.Q(n337));
  MUX21X1 U684(.IN1(n16),.IN2(fract_28_i[4:4]),.S(n22),.Q(n340));
  MUX21X1 U685(.IN1(n337),.IN2(n340),.S(n23),.Q(n351));
  MUX21X1 U686(.IN1(n349),.IN2(n351),.S(n3),.Q(n375));
  MUX21X1 U687(.IN1(fract_28_i[3:3]),.IN2(fract_28_i[2:2]),.S(n22),.Q(n339));
  MUX21X1 U688(.IN1(fract_28_i[1:1]),.IN2(fract_28_i[0:0]),.S(n22),.Q(n341));
  MUX21X1 U689(.IN1(n339),.IN2(n341),.S(n23),.Q(n350));
  MUX21X1 U690(.IN1(n76),.IN2(n377),.S(n2),.Q(n443));
  NOR3X0 U691(.IN1(n443),.IN2(n29),.IN3(n27),.QN(N1010));
  MUX21X1 U692(.IN1(fract_28_i[12:12]),.IN2(n18),.S(n22),.Q(n343));
  MUX21X1 U693(.IN1(n343),.IN2(n330),.S(n23),.Q(n354));
  MUX21X1 U694(.IN1(n332),.IN2(n331),.S(n23),.Q(n355));
  MUX21X1 U695(.IN1(n354),.IN2(n355),.S(n3),.Q(n382));
  MUX21X1 U696(.IN1(n84),.IN2(n85),.S(n23),.Q(n356));
  MUX21X1 U697(.IN1(n356),.IN2(n334),.S(n3),.Q(n385));
  MUX21X1 U698(.IN1(n77),.IN2(n385),.S(n2),.Q(n335));
  NOR3X0 U699(.IN1(n335),.IN2(n29),.IN3(n27),.QN(N1011));
  MUX21X1 U700(.IN1(fract_28_i[13:13]),.IN2(fract_28_i[12:12]),.S(n4),.Q(n348));
  MUX21X1 U701(.IN1(n348),.IN2(n336),.S(n23),.Q(n361));
  MUX21X1 U702(.IN1(n338),.IN2(n337),.S(n23),.Q(n363));
  MUX21X1 U703(.IN1(n361),.IN2(n363),.S(n3),.Q(n389));
  MUX21X1 U704(.IN1(n340),.IN2(n339),.S(n23),.Q(n362));
  MUX21X1 U705(.IN1(n83),.IN2(n365),.S(n3),.Q(n392));
  MUX21X1 U706(.IN1(n78),.IN2(n392),.S(n2),.Q(n342));
  NOR3X0 U707(.IN1(n27),.IN2(n29),.IN3(n342),.QN(N1012));
  MUX21X1 U708(.IN1(fract_28_i[14:14]),.IN2(fract_28_i[13:13]),.S(n4),.Q(n353));
  MUX21X1 U709(.IN1(n353),.IN2(n343),.S(n23),.Q(n368));
  MUX21X1 U710(.IN1(n368),.IN2(n344),.S(n3),.Q(n396));
  MUX21X1 U711(.IN1(n81),.IN2(n346),.S(n3),.Q(n399));
  MUX21X1 U712(.IN1(n79),.IN2(n399),.S(n2),.Q(n347));
  NOR3X0 U713(.IN1(n27),.IN2(n29),.IN3(n347),.QN(N1013));
  MUX21X1 U714(.IN1(fract_28_i[15:15]),.IN2(fract_28_i[14:14]),.S(n4),.Q(n360));
  MUX21X1 U715(.IN1(n360),.IN2(n348),.S(n23),.Q(n374));
  MUX21X1 U716(.IN1(n374),.IN2(n349),.S(n3),.Q(n403));
  MUX21X1 U717(.IN1(n351),.IN2(n350),.S(n24),.Q(n406));
  MUX21X1 U718(.IN1(n403),.IN2(n406),.S(n2),.Q(n352));
  NOR3X0 U719(.IN1(n27),.IN2(n29),.IN3(n62),.QN(N1014));
  MUX21X1 U720(.IN1(fract_28_i[16:16]),.IN2(fract_28_i[15:15]),.S(n4),.Q(n367));
  MUX21X1 U721(.IN1(n367),.IN2(n353),.S(n5),.Q(n381));
  MUX21X1 U722(.IN1(n381),.IN2(n354),.S(n24),.Q(n411));
  MUX21X1 U723(.IN1(n82),.IN2(n356),.S(n24),.Q(n415));
  MUX21X1 U724(.IN1(n80),.IN2(n415),.S(n25),.Q(n358));
  MUX21X1 U725(.IN1(n358),.IN2(n357),.S(n26),.Q(n359));
  MUX21X1 U726(.IN1(n20),.IN2(fract_28_i[16:16]),.S(n4),.Q(n373));
  MUX21X1 U727(.IN1(n373),.IN2(n360),.S(n5),.Q(n388));
  MUX21X1 U728(.IN1(n388),.IN2(n361),.S(n24),.Q(n420));
  MUX21X1 U729(.IN1(n363),.IN2(n362),.S(n24),.Q(n424));
  MUX21X1 U730(.IN1(n420),.IN2(n424),.S(n2),.Q(n364));
  MUX21X1 U731(.IN1(n63),.IN2(n379),.S(n26),.Q(n366));
  MUX21X1 U732(.IN1(fract_28_i[18:18]),.IN2(n20),.S(n4),.Q(n380));
  MUX21X1 U733(.IN1(n380),.IN2(n367),.S(n5),.Q(n395));
  MUX21X1 U734(.IN1(n395),.IN2(n368),.S(n24),.Q(n431));
  MUX21X1 U735(.IN1(n431),.IN2(n369),.S(n2),.Q(n370));
  OR2X1 U736(.IN1(n371),.IN2(n2),.Q(n445));
  MUX21X1 U737(.IN1(n64),.IN2(n445),.S(n26),.Q(n372));
  MUX21X1 U738(.IN1(fract_28_i[19:19]),.IN2(fract_28_i[18:18]),.S(n4),.Q(n387));
  MUX21X1 U739(.IN1(n387),.IN2(n373),.S(n5),.Q(n402));
  MUX21X1 U740(.IN1(n402),.IN2(n374),.S(n24),.Q(n441));
  MUX21X1 U741(.IN1(n441),.IN2(n375),.S(n25),.Q(n376));
  OR2X1 U742(.IN1(n377),.IN2(n2),.Q(n446));
  MUX21X1 U743(.IN1(n65),.IN2(n446),.S(n26),.Q(n378));
  NOR3X0 U744(.IN1(n379),.IN2(n29),.IN3(n27),.QN(N1000));
  MUX21X1 U745(.IN1(fract_28_i[20:20]),.IN2(fract_28_i[19:19]),.S(n4),.Q(n394));
  MUX21X1 U746(.IN1(n394),.IN2(n380),.S(n5),.Q(n409));
  MUX21X1 U747(.IN1(n409),.IN2(n381),.S(n24),.Q(n383));
  MUX21X1 U748(.IN1(n383),.IN2(n382),.S(n25),.Q(n384));
  OR2X1 U749(.IN1(n385),.IN2(n2),.Q(n447));
  MUX21X1 U750(.IN1(n66),.IN2(n447),.S(n26),.Q(n386));
  MUX21X1 U751(.IN1(fract_28_i[21:21]),.IN2(fract_28_i[20:20]),.S(n4),.Q(n401));
  MUX21X1 U752(.IN1(n401),.IN2(n387),.S(n5),.Q(n418));
  MUX21X1 U753(.IN1(n418),.IN2(n388),.S(n24),.Q(n390));
  MUX21X1 U754(.IN1(n390),.IN2(n389),.S(n25),.Q(n391));
  OR2X1 U755(.IN1(n392),.IN2(n2),.Q(n448));
  MUX21X1 U756(.IN1(n67),.IN2(n448),.S(n26),.Q(n393));
  MUX21X1 U757(.IN1(fract_28_i[22:22]),.IN2(fract_28_i[21:21]),.S(n4),.Q(n408));
  MUX21X1 U758(.IN1(n408),.IN2(n394),.S(n5),.Q(n429));
  MUX21X1 U759(.IN1(n429),.IN2(n395),.S(n24),.Q(n397));
  MUX21X1 U760(.IN1(n397),.IN2(n396),.S(n25),.Q(n398));
  OR2X1 U761(.IN1(n399),.IN2(n2),.Q(n449));
  MUX21X1 U762(.IN1(n68),.IN2(n449),.S(n26),.Q(n400));
  MUX21X1 U763(.IN1(fract_28_i[23:23]),.IN2(fract_28_i[22:22]),.S(n4),.Q(n417));
  MUX21X1 U764(.IN1(n417),.IN2(n401),.S(n5),.Q(n438));
  MUX21X1 U765(.IN1(n438),.IN2(n402),.S(n24),.Q(n404));
  MUX21X1 U766(.IN1(n404),.IN2(n403),.S(n25),.Q(n405));
  MUX21X1 U767(.IN1(n69),.IN2(n450),.S(n26),.Q(n407));
  MUX21X1 U768(.IN1(fract_28_i[24:24]),.IN2(fract_28_i[23:23]),.S(n4),.Q(n427));
  MUX21X1 U769(.IN1(n427),.IN2(n408),.S(n5),.Q(n410));
  MUX21X1 U770(.IN1(n410),.IN2(n409),.S(n24),.Q(n412));
  MUX21X1 U771(.IN1(n412),.IN2(n411),.S(n25),.Q(n413));
  MUX21X1 U772(.IN1(n415),.IN2(n74),.S(n25),.Q(n451));
  MUX21X1 U773(.IN1(n70),.IN2(n451),.S(n26),.Q(n416));
  MUX21X1 U774(.IN1(fract_28_i[25:25]),.IN2(fract_28_i[24:24]),.S(n4),.Q(n436));
  MUX21X1 U775(.IN1(n436),.IN2(n417),.S(n5),.Q(n419));
  MUX21X1 U776(.IN1(n419),.IN2(n418),.S(n24),.Q(n421));
  MUX21X1 U777(.IN1(n421),.IN2(n420),.S(n25),.Q(n422));
  MUX21X1 U778(.IN1(n424),.IN2(n423),.S(n25),.Q(n425));
  MUX21X1 U779(.IN1(n71),.IN2(n72),.S(n26),.Q(n426));
  MUX21X1 U780(.IN1(fract_28_i[26:26]),.IN2(fract_28_i[25:25]),.S(n4),.Q(n428));
  MUX21X1 U781(.IN1(n428),.IN2(n427),.S(n5),.Q(n430));
  MUX21X1 U782(.IN1(n430),.IN2(n429),.S(n24),.Q(n432));
  MUX21X1 U783(.IN1(n432),.IN2(n431),.S(n25),.Q(n433));
  MUX21X1 U784(.IN1(n73),.IN2(n434),.S(n26),.Q(n435));
  MUX21X1 U785(.IN1(fract_28_i[27:27]),.IN2(fract_28_i[26:26]),.S(n4),.Q(n437));
  MUX21X1 U786(.IN1(n437),.IN2(n436),.S(n5),.Q(n439));
  MUX21X1 U787(.IN1(n439),.IN2(n438),.S(n24),.Q(n440));
  MUX21X1 U788(.IN1(n441),.IN2(n440),.S(n6),.Q(n442));
  MUX21X1 U789(.IN1(n61),.IN2(n443),.S(n26),.Q(n444));
  NOR3X0 U790(.IN1(n27),.IN2(n29),.IN3(n445),.QN(N1001));
  NOR3X0 U791(.IN1(n27),.IN2(n29),.IN3(n446),.QN(N1002));
  NOR3X0 U792(.IN1(n27),.IN2(n29),.IN3(n447),.QN(N1003));
  NOR3X0 U793(.IN1(n448),.IN2(n29),.IN3(n27),.QN(N1004));
  NOR3X0 U794(.IN1(n449),.IN2(n29),.IN3(n27),.QN(N1005));
  NOR3X0 U795(.IN1(n450),.IN2(n29),.IN3(n27),.QN(N1006));
  NOR3X0 U796(.IN1(n27),.IN2(n29),.IN3(n451),.QN(N1007));
  NOR3X0 U797(.IN1(n72),.IN2(n29),.IN3(n27),.QN(N1008));
endmodule
module pre_norm_mul_DW01_add_1_inj (A,B,CI,SUM,CO);
input [9:0] A ;
input [9:0] B ;
output [9:0] SUM ;
input CI ;
output CO ;
wire [9:1] carry ;
// instances
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(SUM[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(carry[1:1]),.CO(carry[2:2]),.S(SUM[1:1]));
  FADDX1 U1_0(.A(A[0:0]),.B(B[0:0]),.CI(CI),.CO(carry[1:1]),.S(SUM[0:0]));
endmodule
module pre_norm_mul_inj (clk_i,opa_i,opb_i,exp_10_o,fracta_24_o,fractb_24_o);
input [31:0] opa_i ;
input [31:0] opb_i ;
output [9:0] exp_10_o ;
output [23:0] fracta_24_o ;
output [23:0] fractb_24_o ;
input clk_i ;
wire \opa_i[22]  ;
wire \opa_i[21]  ;
wire \opa_i[20]  ;
wire \opa_i[19]  ;
wire \opa_i[18]  ;
wire \opa_i[17]  ;
wire \opa_i[16]  ;
wire \opa_i[15]  ;
wire \opa_i[14]  ;
wire \opa_i[13]  ;
wire \opa_i[12]  ;
wire \opa_i[11]  ;
wire \opa_i[10]  ;
wire \opa_i[9]  ;
wire \opa_i[8]  ;
wire \opa_i[7]  ;
wire \opa_i[6]  ;
wire \opa_i[5]  ;
wire \opa_i[4]  ;
wire \opa_i[3]  ;
wire \opa_i[2]  ;
wire \opa_i[1]  ;
wire \opa_i[0]  ;
wire \opb_i[22]  ;
wire \opb_i[21]  ;
wire \opb_i[20]  ;
wire \opb_i[19]  ;
wire \opb_i[18]  ;
wire \opb_i[17]  ;
wire \opb_i[16]  ;
wire \opb_i[15]  ;
wire \opb_i[14]  ;
wire \opb_i[13]  ;
wire \opb_i[12]  ;
wire \opb_i[11]  ;
wire \opb_i[10]  ;
wire \opb_i[9]  ;
wire \opb_i[8]  ;
wire \opb_i[7]  ;
wire \opb_i[6]  ;
wire \opb_i[5]  ;
wire \opb_i[4]  ;
wire \opb_i[3]  ;
wire \opb_i[2]  ;
wire \opb_i[1]  ;
wire \opb_i[0]  ;
wire N6 ;
wire N13 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire \add_0_root_add_1_root_sub_101/carry[8]  ;
wire \add_0_root_add_1_root_sub_101/carry[7]  ;
wire \add_0_root_add_1_root_sub_101/carry[6]  ;
wire \add_0_root_add_1_root_sub_101/carry[5]  ;
wire \add_0_root_add_1_root_sub_101/carry[4]  ;
wire \add_0_root_add_1_root_sub_101/carry[3]  ;
wire \add_0_root_add_1_root_sub_101/carry[2]  ;
wire \add_0_root_add_1_root_sub_101/carry[1]  ;
wire \add_0_root_add_1_root_sub_101/B[0]  ;
wire \add_0_root_add_1_root_sub_101/B[1]  ;
wire \add_0_root_add_1_root_sub_101/B[2]  ;
wire \add_0_root_add_1_root_sub_101/B[3]  ;
wire \add_0_root_add_1_root_sub_101/B[4]  ;
wire \add_0_root_add_1_root_sub_101/B[5]  ;
wire \add_0_root_add_1_root_sub_101/B[6]  ;
wire \add_0_root_add_1_root_sub_101/B[7]  ;
wire \add_0_root_add_1_root_sub_101/B[8]  ;
wire \add_0_root_add_1_root_sub_101/A[1]  ;
wire n1 ;
wire n2 ;
wire [9:0] s_exp_10_o ;
wire SYNOPSYS_UNCONNECTED__0 ;
// instances
  DFFX1 desc364(.D(n1),.CLK(clk_i),.Q(exp_10_o[9:9]));
  DFFX1 desc365(.D(s_exp_10_o[8:8]),.CLK(clk_i),.Q(exp_10_o[8:8]));
  DFFX1 desc366(.D(s_exp_10_o[7:7]),.CLK(clk_i),.Q(exp_10_o[7:7]));
  DFFX1 desc367(.D(s_exp_10_o[6:6]),.CLK(clk_i),.Q(exp_10_o[6:6]));
  DFFX1 desc368(.D(s_exp_10_o[5:5]),.CLK(clk_i),.Q(exp_10_o[5:5]));
  DFFX1 desc369(.D(s_exp_10_o[4:4]),.CLK(clk_i),.Q(exp_10_o[4:4]));
  DFFX1 desc370(.D(s_exp_10_o[3:3]),.CLK(clk_i),.Q(exp_10_o[3:3]));
  DFFX1 desc371(.D(s_exp_10_o[2:2]),.CLK(clk_i),.Q(exp_10_o[2:2]));
  DFFX1 desc372(.D(s_exp_10_o[1:1]),.CLK(clk_i),.Q(exp_10_o[1:1]));
  DFFX1 desc373(.D(s_exp_10_o[0:0]),.CLK(clk_i),.Q(exp_10_o[0:0]));
  NOR4X0 U7(.IN1(opa_i[30:30]),.IN2(opa_i[29:29]),.IN3(opa_i[28:28]),.IN4(opa_i[27:27]),.QN(n4));
  NOR4X0 U8(.IN1(opa_i[26:26]),.IN2(opa_i[25:25]),.IN3(opa_i[24:24]),.IN4(opa_i[23:23]),.QN(n3));
  NOR4X0 U9(.IN1(opb_i[30:30]),.IN2(opb_i[29:29]),.IN3(opb_i[28:28]),.IN4(opb_i[27:27]),.QN(n6));
  NOR4X0 U10(.IN1(opb_i[26:26]),.IN2(opb_i[25:25]),.IN3(opb_i[24:24]),.IN4(opb_i[23:23]),.QN(n5));
  pre_norm_mul_DW01_add_1_inj add_1_root_add_1_root_sub_101(.A({1'b0,1'b0,opb_i[30:23]}),.B({1'b0,1'b0,opa_i[30:23]}),.CI(n2),.SUM({SYNOPSYS_UNCONNECTED__0,\add_0_root_add_1_root_sub_101/B[8] ,\add_0_root_add_1_root_sub_101/B[7] ,\add_0_root_add_1_root_sub_101/B[6] ,\add_0_root_add_1_root_sub_101/B[5] ,\add_0_root_add_1_root_sub_101/B[4] ,\add_0_root_add_1_root_sub_101/B[3] ,\add_0_root_add_1_root_sub_101/B[2] ,\add_0_root_add_1_root_sub_101/B[1] ,\add_0_root_add_1_root_sub_101/B[0] }));
  FADDX1 desc374(.A(\add_0_root_add_1_root_sub_101/A[1] ),.B(\add_0_root_add_1_root_sub_101/B[1] ),.CI(\add_0_root_add_1_root_sub_101/carry[1] ),.CO(\add_0_root_add_1_root_sub_101/carry[2] ),.S(s_exp_10_o[1:1]));
  NOR2X0 U3(.IN1(\add_0_root_add_1_root_sub_101/B[8] ),.IN2(\add_0_root_add_1_root_sub_101/carry[8] ),.QN(n1));
  INVX0 U4(.INP(N13),.ZN(\add_0_root_add_1_root_sub_101/A[1] ));
  INVX0 U5(.INP(N6),.ZN(n2));
  NAND2X0 U6(.IN1(n3),.IN2(n4),.QN(N6));
  NAND2X1 U11(.IN1(n5),.IN2(n6),.QN(N13));
  XNOR2X1 U12(.IN1(\add_0_root_add_1_root_sub_101/carry[8] ),.IN2(\add_0_root_add_1_root_sub_101/B[8] ),.Q(s_exp_10_o[8:8]));
  OR2X1 U13(.IN1(\add_0_root_add_1_root_sub_101/B[7] ),.IN2(\add_0_root_add_1_root_sub_101/carry[7] ),.Q(\add_0_root_add_1_root_sub_101/carry[8] ));
  XNOR2X1 U14(.IN1(\add_0_root_add_1_root_sub_101/carry[7] ),.IN2(\add_0_root_add_1_root_sub_101/B[7] ),.Q(s_exp_10_o[7:7]));
  AND2X1 U15(.IN1(\add_0_root_add_1_root_sub_101/B[6] ),.IN2(\add_0_root_add_1_root_sub_101/carry[6] ),.Q(\add_0_root_add_1_root_sub_101/carry[7] ));
  XOR2X1 U16(.IN1(\add_0_root_add_1_root_sub_101/B[6] ),.IN2(\add_0_root_add_1_root_sub_101/carry[6] ),.Q(s_exp_10_o[6:6]));
  AND2X1 U17(.IN1(\add_0_root_add_1_root_sub_101/B[5] ),.IN2(\add_0_root_add_1_root_sub_101/carry[5] ),.Q(\add_0_root_add_1_root_sub_101/carry[6] ));
  XOR2X1 U18(.IN1(\add_0_root_add_1_root_sub_101/B[5] ),.IN2(\add_0_root_add_1_root_sub_101/carry[5] ),.Q(s_exp_10_o[5:5]));
  AND2X1 U19(.IN1(\add_0_root_add_1_root_sub_101/B[4] ),.IN2(\add_0_root_add_1_root_sub_101/carry[4] ),.Q(\add_0_root_add_1_root_sub_101/carry[5] ));
  XOR2X1 U20(.IN1(\add_0_root_add_1_root_sub_101/B[4] ),.IN2(\add_0_root_add_1_root_sub_101/carry[4] ),.Q(s_exp_10_o[4:4]));
  AND2X1 U21(.IN1(\add_0_root_add_1_root_sub_101/B[3] ),.IN2(\add_0_root_add_1_root_sub_101/carry[3] ),.Q(\add_0_root_add_1_root_sub_101/carry[4] ));
  XOR2X1 U22(.IN1(\add_0_root_add_1_root_sub_101/B[3] ),.IN2(\add_0_root_add_1_root_sub_101/carry[3] ),.Q(s_exp_10_o[3:3]));
  AND2X1 U23(.IN1(\add_0_root_add_1_root_sub_101/B[2] ),.IN2(\add_0_root_add_1_root_sub_101/carry[2] ),.Q(\add_0_root_add_1_root_sub_101/carry[3] ));
  XOR2X1 U24(.IN1(\add_0_root_add_1_root_sub_101/B[2] ),.IN2(\add_0_root_add_1_root_sub_101/carry[2] ),.Q(s_exp_10_o[2:2]));
  AND2X1 U25(.IN1(N13),.IN2(\add_0_root_add_1_root_sub_101/B[0] ),.Q(\add_0_root_add_1_root_sub_101/carry[1] ));
  XOR2X1 U26(.IN1(N13),.IN2(\add_0_root_add_1_root_sub_101/B[0] ),.Q(s_exp_10_o[0:0]));
assign fracta_24_o[22:22]=\opa_i[22] ;
assign \opa_i[22] =opa_i[22:22];
assign fracta_24_o[21:21]=\opa_i[21] ;
assign \opa_i[21] =opa_i[21:21];
assign fracta_24_o[20:20]=\opa_i[20] ;
assign \opa_i[20] =opa_i[20:20];
assign fracta_24_o[19:19]=\opa_i[19] ;
assign \opa_i[19] =opa_i[19:19];
assign fracta_24_o[18:18]=\opa_i[18] ;
assign \opa_i[18] =opa_i[18:18];
assign fracta_24_o[17:17]=\opa_i[17] ;
assign \opa_i[17] =opa_i[17:17];
assign fracta_24_o[16:16]=\opa_i[16] ;
assign \opa_i[16] =opa_i[16:16];
assign fracta_24_o[15:15]=\opa_i[15] ;
assign \opa_i[15] =opa_i[15:15];
assign fracta_24_o[14:14]=\opa_i[14] ;
assign \opa_i[14] =opa_i[14:14];
assign fracta_24_o[13:13]=\opa_i[13] ;
assign \opa_i[13] =opa_i[13:13];
assign fracta_24_o[12:12]=\opa_i[12] ;
assign \opa_i[12] =opa_i[12:12];
assign fracta_24_o[11:11]=\opa_i[11] ;
assign \opa_i[11] =opa_i[11:11];
assign fracta_24_o[10:10]=\opa_i[10] ;
assign \opa_i[10] =opa_i[10:10];
assign fracta_24_o[9:9]=\opa_i[9] ;
assign \opa_i[9] =opa_i[9:9];
assign fracta_24_o[8:8]=\opa_i[8] ;
assign \opa_i[8] =opa_i[8:8];
assign fracta_24_o[7:7]=\opa_i[7] ;
assign \opa_i[7] =opa_i[7:7];
assign fracta_24_o[6:6]=\opa_i[6] ;
assign \opa_i[6] =opa_i[6:6];
assign fracta_24_o[5:5]=\opa_i[5] ;
assign \opa_i[5] =opa_i[5:5];
assign fracta_24_o[4:4]=\opa_i[4] ;
assign \opa_i[4] =opa_i[4:4];
assign fracta_24_o[3:3]=\opa_i[3] ;
assign \opa_i[3] =opa_i[3:3];
assign fracta_24_o[2:2]=\opa_i[2] ;
assign \opa_i[2] =opa_i[2:2];
assign fracta_24_o[1:1]=\opa_i[1] ;
assign \opa_i[1] =opa_i[1:1];
assign fracta_24_o[0:0]=\opa_i[0] ;
assign \opa_i[0] =opa_i[0:0];
assign fractb_24_o[22:22]=\opb_i[22] ;
assign \opb_i[22] =opb_i[22:22];
assign fractb_24_o[21:21]=\opb_i[21] ;
assign \opb_i[21] =opb_i[21:21];
assign fractb_24_o[20:20]=\opb_i[20] ;
assign \opb_i[20] =opb_i[20:20];
assign fractb_24_o[19:19]=\opb_i[19] ;
assign \opb_i[19] =opb_i[19:19];
assign fractb_24_o[18:18]=\opb_i[18] ;
assign \opb_i[18] =opb_i[18:18];
assign fractb_24_o[17:17]=\opb_i[17] ;
assign \opb_i[17] =opb_i[17:17];
assign fractb_24_o[16:16]=\opb_i[16] ;
assign \opb_i[16] =opb_i[16:16];
assign fractb_24_o[15:15]=\opb_i[15] ;
assign \opb_i[15] =opb_i[15:15];
assign fractb_24_o[14:14]=\opb_i[14] ;
assign \opb_i[14] =opb_i[14:14];
assign fractb_24_o[13:13]=\opb_i[13] ;
assign \opb_i[13] =opb_i[13:13];
assign fractb_24_o[12:12]=\opb_i[12] ;
assign \opb_i[12] =opb_i[12:12];
assign fractb_24_o[11:11]=\opb_i[11] ;
assign \opb_i[11] =opb_i[11:11];
assign fractb_24_o[10:10]=\opb_i[10] ;
assign \opb_i[10] =opb_i[10:10];
assign fractb_24_o[9:9]=\opb_i[9] ;
assign \opb_i[9] =opb_i[9:9];
assign fractb_24_o[8:8]=\opb_i[8] ;
assign \opb_i[8] =opb_i[8:8];
assign fractb_24_o[7:7]=\opb_i[7] ;
assign \opb_i[7] =opb_i[7:7];
assign fractb_24_o[6:6]=\opb_i[6] ;
assign \opb_i[6] =opb_i[6:6];
assign fractb_24_o[5:5]=\opb_i[5] ;
assign \opb_i[5] =opb_i[5:5];
assign fractb_24_o[4:4]=\opb_i[4] ;
assign \opb_i[4] =opb_i[4:4];
assign fractb_24_o[3:3]=\opb_i[3] ;
assign \opb_i[3] =opb_i[3:3];
assign fractb_24_o[2:2]=\opb_i[2] ;
assign \opb_i[2] =opb_i[2:2];
assign fractb_24_o[1:1]=\opb_i[1] ;
assign \opb_i[1] =opb_i[1:1];
assign fractb_24_o[0:0]=\opb_i[0] ;
assign \opb_i[0] =opb_i[0:0];
assign fracta_24_o[23:23]=N6;
assign fractb_24_o[23:23]=N13;
endmodule
module mul_24_DW01_add_3_inj (A,B,CI,SUM,CO);
input [23:0] A ;
input [23:0] B ;
output [23:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire [23:1] carry ;
// instances
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(carry[13:13]),.CO(carry[14:14]),.S(SUM[13:13]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(carry[12:12]),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_11(.A(A[11:11]),.B(B[11:11]),.CI(carry[11:11]),.CO(carry[12:12]),.S(SUM[11:11]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(carry[10:10]),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_9(.A(A[9:9]),.B(B[9:9]),.CI(carry[9:9]),.CO(carry[10:10]),.S(SUM[9:9]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(n1),.CO(carry[8:8]),.S(SUM[7:7]));
  AND2X1 U1(.IN1(A[6:6]),.IN2(B[6:6]),.Q(n1));
  AND2X1 U2(.IN1(A[19:19]),.IN2(carry[19:19]),.Q(n2));
  AND2X1 U3(.IN1(A[20:20]),.IN2(n2),.Q(n3));
  AND2X1 U4(.IN1(A[21:21]),.IN2(n3),.Q(n4));
  NAND2X1 U5(.IN1(A[22:22]),.IN2(n4),.QN(n5));
  XNOR2X1 U6(.IN1(A[23:23]),.IN2(n5),.Q(SUM[23:23]));
  XOR2X1 U7(.IN1(A[6:6]),.IN2(B[6:6]),.Q(SUM[6:6]));
  XOR2X1 U8(.IN1(A[19:19]),.IN2(carry[19:19]),.Q(SUM[19:19]));
  XOR2X1 U9(.IN1(A[20:20]),.IN2(n2),.Q(SUM[20:20]));
  XOR2X1 U10(.IN1(A[21:21]),.IN2(n3),.Q(SUM[21:21]));
  XOR2X1 U11(.IN1(A[22:22]),.IN2(n4),.Q(SUM[22:22]));
assign SUM[5:5]=B[5:5];
assign SUM[4:4]=B[4:4];
assign SUM[3:3]=B[3:3];
assign SUM[2:2]=B[2:2];
assign SUM[1:1]=B[1:1];
assign SUM[0:0]=B[0:0];
endmodule
module mul_24_DW_mult_uns_3_inj (a,b,product);
input [5:0] a ;
input [5:0] b ;
output [11:0] product ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
// instances
  FADDX1 U2(.A(n11),.B(n51),.CI(n2),.CO(product[11:11]),.S(product[10:10]));
  FADDX1 U3(.A(n13),.B(n12),.CI(n3),.CO(n2),.S(product[9:9]));
  FADDX1 U4(.A(n17),.B(n14),.CI(n4),.CO(n3),.S(product[8:8]));
  FADDX1 U5(.A(n18),.B(n23),.CI(n5),.CO(n4),.S(product[7:7]));
  FADDX1 U6(.A(n24),.B(n31),.CI(n6),.CO(n5),.S(product[6:6]));
  FADDX1 U7(.A(n32),.B(n39),.CI(n7),.CO(n6),.S(product[5:5]));
  FADDX1 U8(.A(n40),.B(n45),.CI(n8),.CO(n7),.S(product[4:4]));
  FADDX1 U9(.A(n46),.B(n49),.CI(n9),.CO(n8),.S(product[3:3]));
  FADDX1 U10(.A(n50),.B(n74),.CI(n10),.CO(n9),.S(product[2:2]));
  HADDX1 U11(.A0(n80),.B0(n85),.C1(n10),.SO(product[1:1]));
  FADDX1 U12(.A(n52),.B(n57),.CI(n15),.CO(n11),.S(n12));
  FADDX1 U13(.A(n16),.B(n21),.CI(n19),.CO(n13),.S(n14));
  FADDX1 U14(.A(n53),.B(n63),.CI(n58),.CO(n15),.S(n16));
  FADDX1 U15(.A(n25),.B(n22),.CI(n20),.CO(n17),.S(n18));
  FADDX1 U16(.A(n29),.B(n64),.CI(n27),.CO(n19),.S(n20));
  FADDX1 U17(.A(n54),.B(n69),.CI(n59),.CO(n21),.S(n22));
  FADDX1 U18(.A(n33),.B(n28),.CI(n26),.CO(n23),.S(n24));
  FADDX1 U19(.A(n37),.B(n30),.CI(n35),.CO(n25),.S(n26));
  FADDX1 U20(.A(n70),.B(n65),.CI(n75),.CO(n27),.S(n28));
  HADDX1 U21(.A0(n60),.B0(n55),.C1(n29),.SO(n30));
  FADDX1 U22(.A(n36),.B(n41),.CI(n34),.CO(n31),.S(n32));
  FADDX1 U23(.A(n38),.B(n81),.CI(n43),.CO(n33),.S(n34));
  FADDX1 U24(.A(n66),.B(n71),.CI(n76),.CO(n35),.S(n36));
  HADDX1 U25(.A0(n61),.B0(n56),.C1(n37),.SO(n38));
  FADDX1 U26(.A(n47),.B(n44),.CI(n42),.CO(n39),.S(n40));
  FADDX1 U27(.A(n72),.B(n82),.CI(n77),.CO(n41),.S(n42));
  HADDX1 U28(.A0(n67),.B0(n62),.C1(n43),.SO(n44));
  FADDX1 U29(.A(n78),.B(n83),.CI(n48),.CO(n45),.S(n46));
  HADDX1 U30(.A0(n73),.B0(n68),.C1(n47),.SO(n48));
  HADDX1 U31(.A0(n84),.B0(n79),.C1(n49),.SO(n50));
  INVX0 U82(.INP(a[0:0]),.ZN(n131));
  INVX0 U83(.INP(b[1:1]),.ZN(n136));
  INVX0 U84(.INP(b[0:0]),.ZN(n137));
  INVX0 U85(.INP(b[2:2]),.ZN(n135));
  INVX0 U86(.INP(b[5:5]),.ZN(n132));
  INVX0 U87(.INP(b[3:3]),.ZN(n134));
  INVX0 U88(.INP(b[4:4]),.ZN(n133));
  INVX0 U89(.INP(a[1:1]),.ZN(n130));
  INVX0 U90(.INP(a[2:2]),.ZN(n129));
  INVX0 U91(.INP(a[3:3]),.ZN(n128));
  INVX0 U92(.INP(a[5:5]),.ZN(n126));
  INVX0 U93(.INP(a[4:4]),.ZN(n127));
  NOR2X0 U94(.IN1(n131),.IN2(n137),.QN(product[0:0]));
  NOR2X0 U95(.IN1(n131),.IN2(n136),.QN(n85));
  NOR2X0 U96(.IN1(n131),.IN2(n135),.QN(n84));
  NOR2X0 U97(.IN1(n131),.IN2(n134),.QN(n83));
  NOR2X0 U98(.IN1(n131),.IN2(n133),.QN(n82));
  NOR2X0 U99(.IN1(n131),.IN2(n132),.QN(n81));
  NOR2X0 U100(.IN1(n137),.IN2(n130),.QN(n80));
  NOR2X0 U101(.IN1(n136),.IN2(n130),.QN(n79));
  NOR2X0 U102(.IN1(n135),.IN2(n130),.QN(n78));
  NOR2X0 U103(.IN1(n134),.IN2(n130),.QN(n77));
  NOR2X0 U104(.IN1(n133),.IN2(n130),.QN(n76));
  NOR2X0 U105(.IN1(n132),.IN2(n130),.QN(n75));
  NOR2X0 U106(.IN1(n137),.IN2(n129),.QN(n74));
  NOR2X0 U107(.IN1(n136),.IN2(n129),.QN(n73));
  NOR2X0 U108(.IN1(n135),.IN2(n129),.QN(n72));
  NOR2X0 U109(.IN1(n134),.IN2(n129),.QN(n71));
  NOR2X0 U110(.IN1(n133),.IN2(n129),.QN(n70));
  NOR2X0 U111(.IN1(n132),.IN2(n129),.QN(n69));
  NOR2X0 U112(.IN1(n137),.IN2(n128),.QN(n68));
  NOR2X0 U113(.IN1(n136),.IN2(n128),.QN(n67));
  NOR2X0 U114(.IN1(n135),.IN2(n128),.QN(n66));
  NOR2X0 U115(.IN1(n134),.IN2(n128),.QN(n65));
  NOR2X0 U116(.IN1(n133),.IN2(n128),.QN(n64));
  NOR2X0 U117(.IN1(n132),.IN2(n128),.QN(n63));
  NOR2X0 U118(.IN1(n137),.IN2(n127),.QN(n62));
  NOR2X0 U119(.IN1(n136),.IN2(n127),.QN(n61));
  NOR2X0 U120(.IN1(n135),.IN2(n127),.QN(n60));
  NOR2X0 U121(.IN1(n134),.IN2(n127),.QN(n59));
  NOR2X0 U122(.IN1(n133),.IN2(n127),.QN(n58));
  NOR2X0 U123(.IN1(n132),.IN2(n127),.QN(n57));
  NOR2X0 U124(.IN1(n137),.IN2(n126),.QN(n56));
  NOR2X0 U125(.IN1(n136),.IN2(n126),.QN(n55));
  NOR2X0 U126(.IN1(n135),.IN2(n126),.QN(n54));
  NOR2X0 U127(.IN1(n134),.IN2(n126),.QN(n53));
  NOR2X0 U128(.IN1(n133),.IN2(n126),.QN(n52));
  NOR2X0 U129(.IN1(n132),.IN2(n126),.QN(n51));
endmodule
module mul_24_DW_mult_uns_2_inj (a,b,product);
input [5:0] a ;
input [5:0] b ;
output [11:0] product ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
// instances
  FADDX1 U2(.A(n11),.B(n51),.CI(n2),.CO(product[11:11]),.S(product[10:10]));
  FADDX1 U3(.A(n13),.B(n12),.CI(n3),.CO(n2),.S(product[9:9]));
  FADDX1 U4(.A(n17),.B(n14),.CI(n4),.CO(n3),.S(product[8:8]));
  FADDX1 U5(.A(n18),.B(n23),.CI(n5),.CO(n4),.S(product[7:7]));
  FADDX1 U6(.A(n24),.B(n31),.CI(n6),.CO(n5),.S(product[6:6]));
  FADDX1 U7(.A(n32),.B(n39),.CI(n7),.CO(n6),.S(product[5:5]));
  FADDX1 U8(.A(n40),.B(n45),.CI(n8),.CO(n7),.S(product[4:4]));
  FADDX1 U9(.A(n46),.B(n49),.CI(n9),.CO(n8),.S(product[3:3]));
  FADDX1 U10(.A(n50),.B(n74),.CI(n10),.CO(n9),.S(product[2:2]));
  HADDX1 U11(.A0(n80),.B0(n85),.C1(n10),.SO(product[1:1]));
  FADDX1 U12(.A(n52),.B(n57),.CI(n15),.CO(n11),.S(n12));
  FADDX1 U13(.A(n16),.B(n21),.CI(n19),.CO(n13),.S(n14));
  FADDX1 U14(.A(n53),.B(n63),.CI(n58),.CO(n15),.S(n16));
  FADDX1 U15(.A(n25),.B(n22),.CI(n20),.CO(n17),.S(n18));
  FADDX1 U16(.A(n29),.B(n64),.CI(n27),.CO(n19),.S(n20));
  FADDX1 U17(.A(n54),.B(n69),.CI(n59),.CO(n21),.S(n22));
  FADDX1 U18(.A(n33),.B(n28),.CI(n26),.CO(n23),.S(n24));
  FADDX1 U19(.A(n37),.B(n30),.CI(n35),.CO(n25),.S(n26));
  FADDX1 U20(.A(n70),.B(n65),.CI(n75),.CO(n27),.S(n28));
  HADDX1 U21(.A0(n60),.B0(n55),.C1(n29),.SO(n30));
  FADDX1 U22(.A(n36),.B(n41),.CI(n34),.CO(n31),.S(n32));
  FADDX1 U23(.A(n38),.B(n81),.CI(n43),.CO(n33),.S(n34));
  FADDX1 U24(.A(n66),.B(n71),.CI(n76),.CO(n35),.S(n36));
  HADDX1 U25(.A0(n61),.B0(n56),.C1(n37),.SO(n38));
  FADDX1 U26(.A(n47),.B(n44),.CI(n42),.CO(n39),.S(n40));
  FADDX1 U27(.A(n72),.B(n82),.CI(n77),.CO(n41),.S(n42));
  HADDX1 U28(.A0(n67),.B0(n62),.C1(n43),.SO(n44));
  FADDX1 U29(.A(n78),.B(n83),.CI(n48),.CO(n45),.S(n46));
  HADDX1 U30(.A0(n73),.B0(n68),.C1(n47),.SO(n48));
  HADDX1 U31(.A0(n84),.B0(n79),.C1(n49),.SO(n50));
  INVX0 U82(.INP(a[0:0]),.ZN(n131));
  INVX0 U83(.INP(b[1:1]),.ZN(n136));
  INVX0 U84(.INP(b[0:0]),.ZN(n137));
  INVX0 U85(.INP(b[2:2]),.ZN(n135));
  INVX0 U86(.INP(b[5:5]),.ZN(n132));
  INVX0 U87(.INP(b[3:3]),.ZN(n134));
  INVX0 U88(.INP(b[4:4]),.ZN(n133));
  INVX0 U89(.INP(a[1:1]),.ZN(n130));
  INVX0 U90(.INP(a[2:2]),.ZN(n129));
  INVX0 U91(.INP(a[3:3]),.ZN(n128));
  INVX0 U92(.INP(a[5:5]),.ZN(n126));
  INVX0 U93(.INP(a[4:4]),.ZN(n127));
  NOR2X0 U94(.IN1(n131),.IN2(n137),.QN(product[0:0]));
  NOR2X0 U95(.IN1(n131),.IN2(n136),.QN(n85));
  NOR2X0 U96(.IN1(n131),.IN2(n135),.QN(n84));
  NOR2X0 U97(.IN1(n131),.IN2(n134),.QN(n83));
  NOR2X0 U98(.IN1(n131),.IN2(n133),.QN(n82));
  NOR2X0 U99(.IN1(n131),.IN2(n132),.QN(n81));
  NOR2X0 U100(.IN1(n137),.IN2(n130),.QN(n80));
  NOR2X0 U101(.IN1(n136),.IN2(n130),.QN(n79));
  NOR2X0 U102(.IN1(n135),.IN2(n130),.QN(n78));
  NOR2X0 U103(.IN1(n134),.IN2(n130),.QN(n77));
  NOR2X0 U104(.IN1(n133),.IN2(n130),.QN(n76));
  NOR2X0 U105(.IN1(n132),.IN2(n130),.QN(n75));
  NOR2X0 U106(.IN1(n137),.IN2(n129),.QN(n74));
  NOR2X0 U107(.IN1(n136),.IN2(n129),.QN(n73));
  NOR2X0 U108(.IN1(n135),.IN2(n129),.QN(n72));
  NOR2X0 U109(.IN1(n134),.IN2(n129),.QN(n71));
  NOR2X0 U110(.IN1(n133),.IN2(n129),.QN(n70));
  NOR2X0 U111(.IN1(n132),.IN2(n129),.QN(n69));
  NOR2X0 U112(.IN1(n137),.IN2(n128),.QN(n68));
  NOR2X0 U113(.IN1(n136),.IN2(n128),.QN(n67));
  NOR2X0 U114(.IN1(n135),.IN2(n128),.QN(n66));
  NOR2X0 U115(.IN1(n134),.IN2(n128),.QN(n65));
  NOR2X0 U116(.IN1(n133),.IN2(n128),.QN(n64));
  NOR2X0 U117(.IN1(n132),.IN2(n128),.QN(n63));
  NOR2X0 U118(.IN1(n137),.IN2(n127),.QN(n62));
  NOR2X0 U119(.IN1(n136),.IN2(n127),.QN(n61));
  NOR2X0 U120(.IN1(n135),.IN2(n127),.QN(n60));
  NOR2X0 U121(.IN1(n134),.IN2(n127),.QN(n59));
  NOR2X0 U122(.IN1(n133),.IN2(n127),.QN(n58));
  NOR2X0 U123(.IN1(n132),.IN2(n127),.QN(n57));
  NOR2X0 U124(.IN1(n137),.IN2(n126),.QN(n56));
  NOR2X0 U125(.IN1(n136),.IN2(n126),.QN(n55));
  NOR2X0 U126(.IN1(n135),.IN2(n126),.QN(n54));
  NOR2X0 U127(.IN1(n134),.IN2(n126),.QN(n53));
  NOR2X0 U128(.IN1(n133),.IN2(n126),.QN(n52));
  NOR2X0 U129(.IN1(n132),.IN2(n126),.QN(n51));
endmodule
module mul_24_DW_mult_uns_1_inj (a,b,product);
input [5:0] a ;
input [5:0] b ;
output [11:0] product ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
// instances
  FADDX1 U2(.A(n11),.B(n51),.CI(n2),.CO(product[11:11]),.S(product[10:10]));
  FADDX1 U3(.A(n13),.B(n12),.CI(n3),.CO(n2),.S(product[9:9]));
  FADDX1 U4(.A(n17),.B(n14),.CI(n4),.CO(n3),.S(product[8:8]));
  FADDX1 U5(.A(n18),.B(n23),.CI(n5),.CO(n4),.S(product[7:7]));
  FADDX1 U6(.A(n24),.B(n31),.CI(n6),.CO(n5),.S(product[6:6]));
  FADDX1 U7(.A(n32),.B(n39),.CI(n7),.CO(n6),.S(product[5:5]));
  FADDX1 U8(.A(n40),.B(n45),.CI(n8),.CO(n7),.S(product[4:4]));
  FADDX1 U9(.A(n46),.B(n49),.CI(n9),.CO(n8),.S(product[3:3]));
  FADDX1 U10(.A(n50),.B(n74),.CI(n10),.CO(n9),.S(product[2:2]));
  HADDX1 U11(.A0(n80),.B0(n85),.C1(n10),.SO(product[1:1]));
  FADDX1 U12(.A(n52),.B(n57),.CI(n15),.CO(n11),.S(n12));
  FADDX1 U13(.A(n16),.B(n21),.CI(n19),.CO(n13),.S(n14));
  FADDX1 U14(.A(n53),.B(n63),.CI(n58),.CO(n15),.S(n16));
  FADDX1 U15(.A(n25),.B(n22),.CI(n20),.CO(n17),.S(n18));
  FADDX1 U16(.A(n29),.B(n64),.CI(n27),.CO(n19),.S(n20));
  FADDX1 U17(.A(n54),.B(n69),.CI(n59),.CO(n21),.S(n22));
  FADDX1 U18(.A(n33),.B(n28),.CI(n26),.CO(n23),.S(n24));
  FADDX1 U19(.A(n37),.B(n30),.CI(n35),.CO(n25),.S(n26));
  FADDX1 U20(.A(n70),.B(n65),.CI(n75),.CO(n27),.S(n28));
  HADDX1 U21(.A0(n60),.B0(n55),.C1(n29),.SO(n30));
  FADDX1 U22(.A(n36),.B(n41),.CI(n34),.CO(n31),.S(n32));
  FADDX1 U23(.A(n38),.B(n81),.CI(n43),.CO(n33),.S(n34));
  FADDX1 U24(.A(n66),.B(n71),.CI(n76),.CO(n35),.S(n36));
  HADDX1 U25(.A0(n61),.B0(n56),.C1(n37),.SO(n38));
  FADDX1 U26(.A(n47),.B(n44),.CI(n42),.CO(n39),.S(n40));
  FADDX1 U27(.A(n72),.B(n82),.CI(n77),.CO(n41),.S(n42));
  HADDX1 U28(.A0(n67),.B0(n62),.C1(n43),.SO(n44));
  FADDX1 U29(.A(n78),.B(n83),.CI(n48),.CO(n45),.S(n46));
  HADDX1 U30(.A0(n73),.B0(n68),.C1(n47),.SO(n48));
  HADDX1 U31(.A0(n84),.B0(n79),.C1(n49),.SO(n50));
  INVX0 U82(.INP(a[0:0]),.ZN(n131));
  INVX0 U83(.INP(b[1:1]),.ZN(n136));
  INVX0 U84(.INP(b[0:0]),.ZN(n137));
  INVX0 U85(.INP(b[2:2]),.ZN(n135));
  INVX0 U86(.INP(b[5:5]),.ZN(n132));
  INVX0 U87(.INP(b[3:3]),.ZN(n134));
  INVX0 U88(.INP(b[4:4]),.ZN(n133));
  INVX0 U89(.INP(a[1:1]),.ZN(n130));
  INVX0 U90(.INP(a[2:2]),.ZN(n129));
  INVX0 U91(.INP(a[3:3]),.ZN(n128));
  INVX0 U92(.INP(a[5:5]),.ZN(n126));
  INVX0 U93(.INP(a[4:4]),.ZN(n127));
  NOR2X0 U94(.IN1(n131),.IN2(n137),.QN(product[0:0]));
  NOR2X0 U95(.IN1(n131),.IN2(n136),.QN(n85));
  NOR2X0 U96(.IN1(n131),.IN2(n135),.QN(n84));
  NOR2X0 U97(.IN1(n131),.IN2(n134),.QN(n83));
  NOR2X0 U98(.IN1(n131),.IN2(n133),.QN(n82));
  NOR2X0 U99(.IN1(n131),.IN2(n132),.QN(n81));
  NOR2X0 U100(.IN1(n137),.IN2(n130),.QN(n80));
  NOR2X0 U101(.IN1(n136),.IN2(n130),.QN(n79));
  NOR2X0 U102(.IN1(n135),.IN2(n130),.QN(n78));
  NOR2X0 U103(.IN1(n134),.IN2(n130),.QN(n77));
  NOR2X0 U104(.IN1(n133),.IN2(n130),.QN(n76));
  NOR2X0 U105(.IN1(n132),.IN2(n130),.QN(n75));
  NOR2X0 U106(.IN1(n137),.IN2(n129),.QN(n74));
  NOR2X0 U107(.IN1(n136),.IN2(n129),.QN(n73));
  NOR2X0 U108(.IN1(n135),.IN2(n129),.QN(n72));
  NOR2X0 U109(.IN1(n134),.IN2(n129),.QN(n71));
  NOR2X0 U110(.IN1(n133),.IN2(n129),.QN(n70));
  NOR2X0 U111(.IN1(n132),.IN2(n129),.QN(n69));
  NOR2X0 U112(.IN1(n137),.IN2(n128),.QN(n68));
  NOR2X0 U113(.IN1(n136),.IN2(n128),.QN(n67));
  NOR2X0 U114(.IN1(n135),.IN2(n128),.QN(n66));
  NOR2X0 U115(.IN1(n134),.IN2(n128),.QN(n65));
  NOR2X0 U116(.IN1(n133),.IN2(n128),.QN(n64));
  NOR2X0 U117(.IN1(n132),.IN2(n128),.QN(n63));
  NOR2X0 U118(.IN1(n137),.IN2(n127),.QN(n62));
  NOR2X0 U119(.IN1(n136),.IN2(n127),.QN(n61));
  NOR2X0 U120(.IN1(n135),.IN2(n127),.QN(n60));
  NOR2X0 U121(.IN1(n134),.IN2(n127),.QN(n59));
  NOR2X0 U122(.IN1(n133),.IN2(n127),.QN(n58));
  NOR2X0 U123(.IN1(n132),.IN2(n127),.QN(n57));
  NOR2X0 U124(.IN1(n137),.IN2(n126),.QN(n56));
  NOR2X0 U125(.IN1(n136),.IN2(n126),.QN(n55));
  NOR2X0 U126(.IN1(n135),.IN2(n126),.QN(n54));
  NOR2X0 U127(.IN1(n134),.IN2(n126),.QN(n53));
  NOR2X0 U128(.IN1(n133),.IN2(n126),.QN(n52));
  NOR2X0 U129(.IN1(n132),.IN2(n126),.QN(n51));
endmodule
module mul_24_DW_mult_uns_0_inj (a,b,product);
input [5:0] a ;
input [5:0] b ;
output [11:0] product ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
// instances
  FADDX1 U2(.A(n11),.B(n51),.CI(n2),.CO(product[11:11]),.S(product[10:10]));
  FADDX1 U3(.A(n13),.B(n12),.CI(n3),.CO(n2),.S(product[9:9]));
  FADDX1 U4(.A(n17),.B(n14),.CI(n4),.CO(n3),.S(product[8:8]));
  FADDX1 U5(.A(n18),.B(n23),.CI(n5),.CO(n4),.S(product[7:7]));
  FADDX1 U6(.A(n24),.B(n31),.CI(n6),.CO(n5),.S(product[6:6]));
  FADDX1 U7(.A(n32),.B(n39),.CI(n7),.CO(n6),.S(product[5:5]));
  FADDX1 U8(.A(n40),.B(n45),.CI(n8),.CO(n7),.S(product[4:4]));
  FADDX1 U9(.A(n46),.B(n49),.CI(n9),.CO(n8),.S(product[3:3]));
  FADDX1 U10(.A(n50),.B(n74),.CI(n10),.CO(n9),.S(product[2:2]));
  HADDX1 U11(.A0(n80),.B0(n85),.C1(n10),.SO(product[1:1]));
  FADDX1 U12(.A(n52),.B(n57),.CI(n15),.CO(n11),.S(n12));
  FADDX1 U13(.A(n16),.B(n21),.CI(n19),.CO(n13),.S(n14));
  FADDX1 U14(.A(n53),.B(n63),.CI(n58),.CO(n15),.S(n16));
  FADDX1 U15(.A(n25),.B(n22),.CI(n20),.CO(n17),.S(n18));
  FADDX1 U16(.A(n29),.B(n64),.CI(n27),.CO(n19),.S(n20));
  FADDX1 U17(.A(n54),.B(n69),.CI(n59),.CO(n21),.S(n22));
  FADDX1 U18(.A(n33),.B(n28),.CI(n26),.CO(n23),.S(n24));
  FADDX1 U19(.A(n37),.B(n30),.CI(n35),.CO(n25),.S(n26));
  FADDX1 U20(.A(n70),.B(n65),.CI(n75),.CO(n27),.S(n28));
  HADDX1 U21(.A0(n60),.B0(n55),.C1(n29),.SO(n30));
  FADDX1 U22(.A(n36),.B(n41),.CI(n34),.CO(n31),.S(n32));
  FADDX1 U23(.A(n38),.B(n81),.CI(n43),.CO(n33),.S(n34));
  FADDX1 U24(.A(n66),.B(n71),.CI(n76),.CO(n35),.S(n36));
  HADDX1 U25(.A0(n61),.B0(n56),.C1(n37),.SO(n38));
  FADDX1 U26(.A(n47),.B(n44),.CI(n42),.CO(n39),.S(n40));
  FADDX1 U27(.A(n72),.B(n82),.CI(n77),.CO(n41),.S(n42));
  HADDX1 U28(.A0(n67),.B0(n62),.C1(n43),.SO(n44));
  FADDX1 U29(.A(n78),.B(n83),.CI(n48),.CO(n45),.S(n46));
  HADDX1 U30(.A0(n73),.B0(n68),.C1(n47),.SO(n48));
  HADDX1 U31(.A0(n84),.B0(n79),.C1(n49),.SO(n50));
  INVX0 U82(.INP(a[0:0]),.ZN(n131));
  INVX0 U83(.INP(b[1:1]),.ZN(n136));
  INVX0 U84(.INP(b[0:0]),.ZN(n137));
  INVX0 U85(.INP(b[2:2]),.ZN(n135));
  INVX0 U86(.INP(b[5:5]),.ZN(n132));
  INVX0 U87(.INP(b[3:3]),.ZN(n134));
  INVX0 U88(.INP(b[4:4]),.ZN(n133));
  INVX0 U89(.INP(a[1:1]),.ZN(n130));
  INVX0 U90(.INP(a[2:2]),.ZN(n129));
  INVX0 U91(.INP(a[3:3]),.ZN(n128));
  INVX0 U92(.INP(a[5:5]),.ZN(n126));
  INVX0 U93(.INP(a[4:4]),.ZN(n127));
  NOR2X0 U94(.IN1(n131),.IN2(n137),.QN(product[0:0]));
  NOR2X0 U95(.IN1(n131),.IN2(n136),.QN(n85));
  NOR2X0 U96(.IN1(n131),.IN2(n135),.QN(n84));
  NOR2X0 U97(.IN1(n131),.IN2(n134),.QN(n83));
  NOR2X0 U98(.IN1(n131),.IN2(n133),.QN(n82));
  NOR2X0 U99(.IN1(n131),.IN2(n132),.QN(n81));
  NOR2X0 U100(.IN1(n137),.IN2(n130),.QN(n80));
  NOR2X0 U101(.IN1(n136),.IN2(n130),.QN(n79));
  NOR2X0 U102(.IN1(n135),.IN2(n130),.QN(n78));
  NOR2X0 U103(.IN1(n134),.IN2(n130),.QN(n77));
  NOR2X0 U104(.IN1(n133),.IN2(n130),.QN(n76));
  NOR2X0 U105(.IN1(n132),.IN2(n130),.QN(n75));
  NOR2X0 U106(.IN1(n137),.IN2(n129),.QN(n74));
  NOR2X0 U107(.IN1(n136),.IN2(n129),.QN(n73));
  NOR2X0 U108(.IN1(n135),.IN2(n129),.QN(n72));
  NOR2X0 U109(.IN1(n134),.IN2(n129),.QN(n71));
  NOR2X0 U110(.IN1(n133),.IN2(n129),.QN(n70));
  NOR2X0 U111(.IN1(n132),.IN2(n129),.QN(n69));
  NOR2X0 U112(.IN1(n137),.IN2(n128),.QN(n68));
  NOR2X0 U113(.IN1(n136),.IN2(n128),.QN(n67));
  NOR2X0 U114(.IN1(n135),.IN2(n128),.QN(n66));
  NOR2X0 U115(.IN1(n134),.IN2(n128),.QN(n65));
  NOR2X0 U116(.IN1(n133),.IN2(n128),.QN(n64));
  NOR2X0 U117(.IN1(n132),.IN2(n128),.QN(n63));
  NOR2X0 U118(.IN1(n137),.IN2(n127),.QN(n62));
  NOR2X0 U119(.IN1(n136),.IN2(n127),.QN(n61));
  NOR2X0 U120(.IN1(n135),.IN2(n127),.QN(n60));
  NOR2X0 U121(.IN1(n134),.IN2(n127),.QN(n59));
  NOR2X0 U122(.IN1(n133),.IN2(n127),.QN(n58));
  NOR2X0 U123(.IN1(n132),.IN2(n127),.QN(n57));
  NOR2X0 U124(.IN1(n137),.IN2(n126),.QN(n56));
  NOR2X0 U125(.IN1(n136),.IN2(n126),.QN(n55));
  NOR2X0 U126(.IN1(n135),.IN2(n126),.QN(n54));
  NOR2X0 U127(.IN1(n134),.IN2(n126),.QN(n53));
  NOR2X0 U128(.IN1(n133),.IN2(n126),.QN(n52));
  NOR2X0 U129(.IN1(n132),.IN2(n126),.QN(n51));
endmodule
module mul_24_DW01_add_2_inj (A,B,CI,SUM,CO);
input [47:0] A ;
input [47:0] B ;
output [47:0] SUM ;
input CI ;
output CO ;
wire \A[0]  ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire [47:1] carry ;
// instances
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(n2),.CO(carry[14:14]),.S(SUM[13:13]));
  AND2X1 U1(.IN1(B[35:35]),.IN2(n13),.Q(SUM[36:36]));
  AND2X1 U2(.IN1(A[12:12]),.IN2(B[12:12]),.Q(n2));
  AND2X1 U3(.IN1(B[24:24]),.IN2(carry[24:24]),.Q(n3));
  AND2X1 U4(.IN1(B[25:25]),.IN2(n3),.Q(n4));
  AND2X1 U5(.IN1(B[26:26]),.IN2(n4),.Q(n5));
  AND2X1 U6(.IN1(B[27:27]),.IN2(n5),.Q(n6));
  AND2X1 U7(.IN1(B[28:28]),.IN2(n6),.Q(n7));
  AND2X1 U8(.IN1(B[29:29]),.IN2(n7),.Q(n8));
  AND2X1 U9(.IN1(B[30:30]),.IN2(n8),.Q(n9));
  AND2X1 U10(.IN1(B[31:31]),.IN2(n9),.Q(n10));
  AND2X1 U11(.IN1(B[32:32]),.IN2(n10),.Q(n11));
  AND2X1 U12(.IN1(B[33:33]),.IN2(n11),.Q(n12));
  AND2X1 U13(.IN1(B[34:34]),.IN2(n12),.Q(n13));
  XOR2X1 U14(.IN1(B[35:35]),.IN2(n13),.Q(SUM[35:35]));
  XOR2X1 U15(.IN1(B[34:34]),.IN2(n12),.Q(SUM[34:34]));
  XOR2X1 U16(.IN1(B[33:33]),.IN2(n11),.Q(SUM[33:33]));
  XOR2X1 U17(.IN1(B[32:32]),.IN2(n10),.Q(SUM[32:32]));
  XOR2X1 U18(.IN1(B[31:31]),.IN2(n9),.Q(SUM[31:31]));
  XOR2X1 U19(.IN1(B[30:30]),.IN2(n8),.Q(SUM[30:30]));
  XOR2X1 U20(.IN1(B[29:29]),.IN2(n7),.Q(SUM[29:29]));
  XOR2X1 U21(.IN1(B[28:28]),.IN2(n6),.Q(SUM[28:28]));
  XOR2X1 U22(.IN1(B[27:27]),.IN2(n5),.Q(SUM[27:27]));
  XOR2X1 U23(.IN1(B[26:26]),.IN2(n4),.Q(SUM[26:26]));
  XOR2X1 U24(.IN1(B[25:25]),.IN2(n3),.Q(SUM[25:25]));
  XOR2X1 U25(.IN1(B[24:24]),.IN2(carry[24:24]),.Q(SUM[24:24]));
  XOR2X1 U26(.IN1(A[12:12]),.IN2(B[12:12]),.Q(SUM[12:12]));
assign SUM[11:11]=A[11:11];
assign SUM[10:10]=A[10:10];
assign SUM[9:9]=A[9:9];
assign SUM[8:8]=A[8:8];
assign SUM[7:7]=A[7:7];
assign SUM[6:6]=A[6:6];
assign SUM[5:5]=A[5:5];
assign SUM[4:4]=A[4:4];
assign SUM[3:3]=A[3:3];
assign SUM[2:2]=A[2:2];
assign SUM[1:1]=A[1:1];
assign SUM[0:0]=\A[0] ;
assign \A[0] =A[0:0];
endmodule
module mul_24_DW01_add_1_inj (A,B,CI,SUM,CO);
input [47:0] A ;
input [47:0] B ;
output [47:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire [47:1] carry ;
// instances
  FADDX1 U1_35(.A(A[35:35]),.B(B[35:35]),.CI(carry[35:35]),.CO(carry[36:36]),.S(SUM[35:35]));
  FADDX1 U1_34(.A(A[34:34]),.B(B[34:34]),.CI(carry[34:34]),.CO(carry[35:35]),.S(SUM[34:34]));
  FADDX1 U1_33(.A(A[33:33]),.B(B[33:33]),.CI(carry[33:33]),.CO(carry[34:34]),.S(SUM[33:33]));
  FADDX1 U1_32(.A(A[32:32]),.B(B[32:32]),.CI(carry[32:32]),.CO(carry[33:33]),.S(SUM[32:32]));
  FADDX1 U1_31(.A(A[31:31]),.B(B[31:31]),.CI(carry[31:31]),.CO(carry[32:32]),.S(SUM[31:31]));
  FADDX1 U1_30(.A(A[30:30]),.B(B[30:30]),.CI(carry[30:30]),.CO(carry[31:31]),.S(SUM[30:30]));
  FADDX1 U1_29(.A(A[29:29]),.B(B[29:29]),.CI(carry[29:29]),.CO(carry[30:30]),.S(SUM[29:29]));
  FADDX1 U1_28(.A(A[28:28]),.B(B[28:28]),.CI(carry[28:28]),.CO(carry[29:29]),.S(SUM[28:28]));
  FADDX1 U1_27(.A(A[27:27]),.B(B[27:27]),.CI(carry[27:27]),.CO(carry[28:28]),.S(SUM[27:27]));
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(carry[26:26]),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_25(.A(A[25:25]),.B(B[25:25]),.CI(n2),.CO(carry[26:26]),.S(SUM[25:25]));
  AND2X1 U1(.IN1(B[46:46]),.IN2(n10),.Q(n1));
  AND2X1 U2(.IN1(A[24:24]),.IN2(B[24:24]),.Q(n2));
  AND2X1 U3(.IN1(B[38:38]),.IN2(n12),.Q(n3));
  AND2X1 U4(.IN1(B[39:39]),.IN2(n3),.Q(n4));
  AND2X1 U5(.IN1(B[40:40]),.IN2(n4),.Q(n5));
  AND2X1 U6(.IN1(B[41:41]),.IN2(n5),.Q(n6));
  AND2X1 U7(.IN1(B[42:42]),.IN2(n6),.Q(n7));
  AND2X1 U8(.IN1(B[43:43]),.IN2(n7),.Q(n8));
  AND2X1 U9(.IN1(B[44:44]),.IN2(n8),.Q(n9));
  AND2X1 U10(.IN1(B[45:45]),.IN2(n9),.Q(n10));
  AND2X1 U11(.IN1(B[36:36]),.IN2(carry[36:36]),.Q(n11));
  AND2X1 U12(.IN1(B[37:37]),.IN2(n11),.Q(n12));
  XOR2X1 U13(.IN1(B[47:47]),.IN2(n1),.Q(SUM[47:47]));
  XOR2X1 U14(.IN1(B[46:46]),.IN2(n10),.Q(SUM[46:46]));
  XOR2X1 U15(.IN1(B[45:45]),.IN2(n9),.Q(SUM[45:45]));
  XOR2X1 U16(.IN1(B[44:44]),.IN2(n8),.Q(SUM[44:44]));
  XOR2X1 U17(.IN1(B[43:43]),.IN2(n7),.Q(SUM[43:43]));
  XOR2X1 U18(.IN1(B[42:42]),.IN2(n6),.Q(SUM[42:42]));
  XOR2X1 U19(.IN1(B[41:41]),.IN2(n5),.Q(SUM[41:41]));
  XOR2X1 U20(.IN1(B[40:40]),.IN2(n4),.Q(SUM[40:40]));
  XOR2X1 U21(.IN1(B[39:39]),.IN2(n3),.Q(SUM[39:39]));
  XOR2X1 U22(.IN1(B[38:38]),.IN2(n12),.Q(SUM[38:38]));
  XOR2X1 U23(.IN1(B[37:37]),.IN2(n11),.Q(SUM[37:37]));
  XOR2X1 U24(.IN1(B[36:36]),.IN2(carry[36:36]),.Q(SUM[36:36]));
  XOR2X1 U25(.IN1(A[24:24]),.IN2(B[24:24]),.Q(SUM[24:24]));
assign SUM[23:23]=A[23:23];
assign SUM[22:22]=A[22:22];
assign SUM[21:21]=A[21:21];
assign SUM[20:20]=A[20:20];
assign SUM[19:19]=A[19:19];
assign SUM[18:18]=A[18:18];
assign SUM[17:17]=A[17:17];
assign SUM[16:16]=A[16:16];
assign SUM[15:15]=A[15:15];
assign SUM[14:14]=A[14:14];
assign SUM[13:13]=A[13:13];
assign SUM[12:12]=A[12:12];
endmodule
module mul_24_DW01_add_0_inj (A,B,CI,SUM,CO);
input [47:0] A ;
input [47:0] B ;
output [47:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire [47:1] carry ;
// instances
  FADDX1 U1_36(.A(A[36:36]),.B(B[36:36]),.CI(carry[36:36]),.CO(carry[37:37]),.S(SUM[36:36]));
  FADDX1 U1_35(.A(A[35:35]),.B(B[35:35]),.CI(carry[35:35]),.CO(carry[36:36]),.S(SUM[35:35]));
  FADDX1 U1_34(.A(A[34:34]),.B(B[34:34]),.CI(carry[34:34]),.CO(carry[35:35]),.S(SUM[34:34]));
  FADDX1 U1_33(.A(A[33:33]),.B(B[33:33]),.CI(carry[33:33]),.CO(carry[34:34]),.S(SUM[33:33]));
  FADDX1 U1_32(.A(A[32:32]),.B(B[32:32]),.CI(carry[32:32]),.CO(carry[33:33]),.S(SUM[32:32]));
  FADDX1 U1_31(.A(A[31:31]),.B(B[31:31]),.CI(carry[31:31]),.CO(carry[32:32]),.S(SUM[31:31]));
  FADDX1 U1_30(.A(A[30:30]),.B(B[30:30]),.CI(carry[30:30]),.CO(carry[31:31]),.S(SUM[30:30]));
  FADDX1 U1_29(.A(A[29:29]),.B(B[29:29]),.CI(carry[29:29]),.CO(carry[30:30]),.S(SUM[29:29]));
  FADDX1 U1_28(.A(A[28:28]),.B(B[28:28]),.CI(carry[28:28]),.CO(carry[29:29]),.S(SUM[28:28]));
  FADDX1 U1_27(.A(A[27:27]),.B(B[27:27]),.CI(carry[27:27]),.CO(carry[28:28]),.S(SUM[27:27]));
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(carry[26:26]),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_25(.A(A[25:25]),.B(B[25:25]),.CI(carry[25:25]),.CO(carry[26:26]),.S(SUM[25:25]));
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(carry[24:24]),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(n10),.CO(carry[14:14]),.S(SUM[13:13]));
  AND2X1 U1(.IN1(A[37:37]),.IN2(carry[37:37]),.Q(n1));
  AND2X1 U2(.IN1(A[38:38]),.IN2(n1),.Q(n2));
  AND2X1 U3(.IN1(A[39:39]),.IN2(n2),.Q(n3));
  AND2X1 U4(.IN1(A[41:41]),.IN2(n9),.Q(n4));
  AND2X1 U5(.IN1(A[42:42]),.IN2(n4),.Q(n5));
  AND2X1 U6(.IN1(A[43:43]),.IN2(n5),.Q(n6));
  AND2X1 U7(.IN1(A[44:44]),.IN2(n6),.Q(n7));
  AND2X1 U8(.IN1(A[45:45]),.IN2(n7),.Q(n8));
  AND2X1 U9(.IN1(A[40:40]),.IN2(n3),.Q(n9));
  NAND2X0 U10(.IN1(A[46:46]),.IN2(n8),.QN(n11));
  AND2X1 U11(.IN1(A[12:12]),.IN2(B[12:12]),.Q(n10));
  XNOR2X1 U12(.IN1(A[47:47]),.IN2(n11),.Q(SUM[47:47]));
  XOR2X1 U13(.IN1(A[46:46]),.IN2(n8),.Q(SUM[46:46]));
  XOR2X1 U14(.IN1(A[45:45]),.IN2(n7),.Q(SUM[45:45]));
  XOR2X1 U15(.IN1(A[44:44]),.IN2(n6),.Q(SUM[44:44]));
  XOR2X1 U16(.IN1(A[43:43]),.IN2(n5),.Q(SUM[43:43]));
  XOR2X1 U17(.IN1(A[42:42]),.IN2(n4),.Q(SUM[42:42]));
  XOR2X1 U18(.IN1(A[41:41]),.IN2(n9),.Q(SUM[41:41]));
  XOR2X1 U19(.IN1(A[40:40]),.IN2(n3),.Q(SUM[40:40]));
  XOR2X1 U20(.IN1(A[39:39]),.IN2(n2),.Q(SUM[39:39]));
  XOR2X1 U21(.IN1(A[38:38]),.IN2(n1),.Q(SUM[38:38]));
  XOR2X1 U22(.IN1(A[37:37]),.IN2(carry[37:37]),.Q(SUM[37:37]));
  XOR2X1 U23(.IN1(A[12:12]),.IN2(B[12:12]),.Q(SUM[12:12]));
assign SUM[11:11]=B[11:11];
assign SUM[10:10]=B[10:10];
assign SUM[9:9]=B[9:9];
assign SUM[8:8]=B[8:8];
assign SUM[7:7]=B[7:7];
assign SUM[6:6]=B[6:6];
assign SUM[5:5]=B[5:5];
assign SUM[4:4]=B[4:4];
assign SUM[3:3]=B[3:3];
assign SUM[2:2]=B[2:2];
assign SUM[1:1]=B[1:1];
assign SUM[0:0]=B[0:0];
endmodule
module mul_24_inj (clk_i,fracta_i,fractb_i,signa_i,signb_i,start_i,fract_o,sign_o,ready_o);
input [23:0] fracta_i ;
input [23:0] fractb_i ;
output [47:0] fract_o ;
input clk_i ;
input signa_i ;
input signb_i ;
input start_i ;
output sign_o ;
output ready_o ;
wire N25 ;
wire N26 ;
wire N34 ;
wire s_signa_i ;
wire s_signb_i ;
wire s_start_i ;
wire s_state ;
wire \count[2]  ;
wire N57 ;
wire N58 ;
wire N59 ;
wire N60 ;
wire N61 ;
wire N62 ;
wire N63 ;
wire N64 ;
wire N65 ;
wire N66 ;
wire N67 ;
wire N68 ;
wire \prod2[3][3][11]  ;
wire \prod2[3][3][10]  ;
wire \prod2[3][3][9]  ;
wire \prod2[3][3][8]  ;
wire \prod2[3][3][7]  ;
wire \prod2[3][3][6]  ;
wire \prod2[3][3][5]  ;
wire \prod2[3][3][4]  ;
wire \prod2[3][3][3]  ;
wire \prod2[3][3][2]  ;
wire \prod2[3][3][1]  ;
wire \prod2[3][3][0]  ;
wire \prod2[3][2][17]  ;
wire \prod2[3][2][16]  ;
wire \prod2[3][2][15]  ;
wire \prod2[3][2][14]  ;
wire \prod2[3][2][13]  ;
wire \prod2[3][2][12]  ;
wire \prod2[3][2][11]  ;
wire \prod2[3][2][10]  ;
wire \prod2[3][2][9]  ;
wire \prod2[3][2][8]  ;
wire \prod2[3][2][7]  ;
wire \prod2[3][2][6]  ;
wire \prod2[3][1][17]  ;
wire \prod2[3][1][16]  ;
wire \prod2[3][1][15]  ;
wire \prod2[3][1][14]  ;
wire \prod2[3][1][13]  ;
wire \prod2[3][1][12]  ;
wire \prod2[3][1][11]  ;
wire \prod2[3][1][10]  ;
wire \prod2[3][1][9]  ;
wire \prod2[3][1][8]  ;
wire \prod2[3][1][7]  ;
wire \prod2[3][1][6]  ;
wire \prod2[3][0][23]  ;
wire \prod2[3][0][22]  ;
wire \prod2[3][0][21]  ;
wire \prod2[3][0][20]  ;
wire \prod2[3][0][19]  ;
wire \prod2[3][0][18]  ;
wire \prod2[3][0][17]  ;
wire \prod2[3][0][16]  ;
wire \prod2[3][0][15]  ;
wire \prod2[3][0][14]  ;
wire \prod2[3][0][13]  ;
wire \prod2[3][0][12]  ;
wire \prod2[2][3][11]  ;
wire \prod2[2][3][10]  ;
wire \prod2[2][3][9]  ;
wire \prod2[2][3][8]  ;
wire \prod2[2][3][7]  ;
wire \prod2[2][3][6]  ;
wire \prod2[2][3][5]  ;
wire \prod2[2][3][4]  ;
wire \prod2[2][3][3]  ;
wire \prod2[2][3][2]  ;
wire \prod2[2][3][1]  ;
wire \prod2[2][3][0]  ;
wire \prod2[2][2][17]  ;
wire \prod2[2][2][16]  ;
wire \prod2[2][2][15]  ;
wire \prod2[2][2][14]  ;
wire \prod2[2][2][13]  ;
wire \prod2[2][2][12]  ;
wire \prod2[2][2][11]  ;
wire \prod2[2][2][10]  ;
wire \prod2[2][2][9]  ;
wire \prod2[2][2][8]  ;
wire \prod2[2][2][7]  ;
wire \prod2[2][2][6]  ;
wire \prod2[2][1][17]  ;
wire \prod2[2][1][16]  ;
wire \prod2[2][1][15]  ;
wire \prod2[2][1][14]  ;
wire \prod2[2][1][13]  ;
wire \prod2[2][1][12]  ;
wire \prod2[2][1][11]  ;
wire \prod2[2][1][10]  ;
wire \prod2[2][1][9]  ;
wire \prod2[2][1][8]  ;
wire \prod2[2][1][7]  ;
wire \prod2[2][1][6]  ;
wire \prod2[2][0][23]  ;
wire \prod2[2][0][22]  ;
wire \prod2[2][0][21]  ;
wire \prod2[2][0][20]  ;
wire \prod2[2][0][19]  ;
wire \prod2[2][0][18]  ;
wire \prod2[2][0][17]  ;
wire \prod2[2][0][16]  ;
wire \prod2[2][0][15]  ;
wire \prod2[2][0][14]  ;
wire \prod2[2][0][13]  ;
wire \prod2[2][0][12]  ;
wire \prod2[1][3][11]  ;
wire \prod2[1][3][10]  ;
wire \prod2[1][3][9]  ;
wire \prod2[1][3][8]  ;
wire \prod2[1][3][7]  ;
wire \prod2[1][3][6]  ;
wire \prod2[1][3][5]  ;
wire \prod2[1][3][4]  ;
wire \prod2[1][3][3]  ;
wire \prod2[1][3][2]  ;
wire \prod2[1][3][1]  ;
wire \prod2[1][3][0]  ;
wire \prod2[1][2][17]  ;
wire \prod2[1][2][16]  ;
wire \prod2[1][2][15]  ;
wire \prod2[1][2][14]  ;
wire \prod2[1][2][13]  ;
wire \prod2[1][2][12]  ;
wire \prod2[1][2][11]  ;
wire \prod2[1][2][10]  ;
wire \prod2[1][2][9]  ;
wire \prod2[1][2][8]  ;
wire \prod2[1][2][7]  ;
wire \prod2[1][2][6]  ;
wire \prod2[1][1][17]  ;
wire \prod2[1][1][16]  ;
wire \prod2[1][1][15]  ;
wire \prod2[1][1][14]  ;
wire \prod2[1][1][13]  ;
wire \prod2[1][1][12]  ;
wire \prod2[1][1][11]  ;
wire \prod2[1][1][10]  ;
wire \prod2[1][1][9]  ;
wire \prod2[1][1][8]  ;
wire \prod2[1][1][7]  ;
wire \prod2[1][1][6]  ;
wire \prod2[1][0][23]  ;
wire \prod2[1][0][22]  ;
wire \prod2[1][0][21]  ;
wire \prod2[1][0][20]  ;
wire \prod2[1][0][19]  ;
wire \prod2[1][0][18]  ;
wire \prod2[1][0][17]  ;
wire \prod2[1][0][16]  ;
wire \prod2[1][0][15]  ;
wire \prod2[1][0][14]  ;
wire \prod2[1][0][13]  ;
wire \prod2[1][0][12]  ;
wire \prod2[0][3][11]  ;
wire \prod2[0][3][10]  ;
wire \prod2[0][3][9]  ;
wire \prod2[0][3][8]  ;
wire \prod2[0][3][7]  ;
wire \prod2[0][3][6]  ;
wire \prod2[0][3][5]  ;
wire \prod2[0][3][4]  ;
wire \prod2[0][3][3]  ;
wire \prod2[0][3][2]  ;
wire \prod2[0][3][1]  ;
wire \prod2[0][3][0]  ;
wire \prod2[0][2][17]  ;
wire \prod2[0][2][16]  ;
wire \prod2[0][2][15]  ;
wire \prod2[0][2][14]  ;
wire \prod2[0][2][13]  ;
wire \prod2[0][2][12]  ;
wire \prod2[0][2][11]  ;
wire \prod2[0][2][10]  ;
wire \prod2[0][2][9]  ;
wire \prod2[0][2][8]  ;
wire \prod2[0][2][7]  ;
wire \prod2[0][2][6]  ;
wire \prod2[0][1][17]  ;
wire \prod2[0][1][16]  ;
wire \prod2[0][1][15]  ;
wire \prod2[0][1][14]  ;
wire \prod2[0][1][13]  ;
wire \prod2[0][1][12]  ;
wire \prod2[0][1][11]  ;
wire \prod2[0][1][10]  ;
wire \prod2[0][1][9]  ;
wire \prod2[0][1][8]  ;
wire \prod2[0][1][7]  ;
wire \prod2[0][1][6]  ;
wire \prod2[0][0][23]  ;
wire \prod2[0][0][22]  ;
wire \prod2[0][0][21]  ;
wire \prod2[0][0][20]  ;
wire \prod2[0][0][19]  ;
wire \prod2[0][0][18]  ;
wire \prod2[0][0][17]  ;
wire \prod2[0][0][16]  ;
wire \prod2[0][0][15]  ;
wire \prod2[0][0][14]  ;
wire \prod2[0][0][13]  ;
wire \prod2[0][0][12]  ;
wire N69 ;
wire N70 ;
wire N71 ;
wire N72 ;
wire N73 ;
wire N74 ;
wire N75 ;
wire N76 ;
wire N77 ;
wire N78 ;
wire N79 ;
wire N80 ;
wire N81 ;
wire N82 ;
wire N83 ;
wire N84 ;
wire N85 ;
wire N86 ;
wire N87 ;
wire N88 ;
wire N89 ;
wire N90 ;
wire N91 ;
wire N92 ;
wire N93 ;
wire N94 ;
wire N95 ;
wire N96 ;
wire N97 ;
wire N98 ;
wire N99 ;
wire N100 ;
wire N101 ;
wire N102 ;
wire N103 ;
wire N104 ;
wire N105 ;
wire N106 ;
wire N107 ;
wire N108 ;
wire N109 ;
wire N110 ;
wire N111 ;
wire N112 ;
wire N113 ;
wire N114 ;
wire N115 ;
wire N116 ;
wire N117 ;
wire N118 ;
wire N119 ;
wire N120 ;
wire N121 ;
wire N122 ;
wire N123 ;
wire N124 ;
wire N125 ;
wire N126 ;
wire N127 ;
wire N128 ;
wire N132 ;
wire N144 ;
wire N152 ;
wire N153 ;
wire N154 ;
wire N155 ;
wire N156 ;
wire N157 ;
wire N158 ;
wire N159 ;
wire N160 ;
wire N161 ;
wire N162 ;
wire N163 ;
wire N182 ;
wire N183 ;
wire N184 ;
wire N185 ;
wire N186 ;
wire N187 ;
wire N188 ;
wire N189 ;
wire N190 ;
wire N191 ;
wire N192 ;
wire N193 ;
wire N232 ;
wire N233 ;
wire N234 ;
wire N235 ;
wire N236 ;
wire N237 ;
wire N288 ;
wire N289 ;
wire N290 ;
wire N291 ;
wire N292 ;
wire N293 ;
wire N300 ;
wire N301 ;
wire N302 ;
wire N303 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N308 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N313 ;
wire N314 ;
wire N315 ;
wire N316 ;
wire N317 ;
wire N318 ;
wire N319 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire \sum[3][23]  ;
wire \sum[3][22]  ;
wire \sum[3][21]  ;
wire \sum[3][20]  ;
wire \sum[3][19]  ;
wire \sum[3][18]  ;
wire \sum[3][17]  ;
wire \sum[3][16]  ;
wire \sum[3][15]  ;
wire \sum[3][14]  ;
wire \sum[3][13]  ;
wire \sum[3][12]  ;
wire \sum[3][11]  ;
wire \sum[3][10]  ;
wire \sum[3][9]  ;
wire \sum[3][8]  ;
wire \sum[3][7]  ;
wire \sum[3][6]  ;
wire \sum[3][5]  ;
wire \sum[3][4]  ;
wire \sum[3][3]  ;
wire \sum[3][2]  ;
wire \sum[3][1]  ;
wire \sum[3][0]  ;
wire \sum[2][23]  ;
wire \sum[2][22]  ;
wire \sum[2][21]  ;
wire \sum[2][20]  ;
wire \sum[2][19]  ;
wire \sum[2][18]  ;
wire \sum[2][17]  ;
wire \sum[2][16]  ;
wire \sum[2][15]  ;
wire \sum[2][14]  ;
wire \sum[2][13]  ;
wire \sum[2][12]  ;
wire \sum[2][11]  ;
wire \sum[2][10]  ;
wire \sum[2][9]  ;
wire \sum[2][8]  ;
wire \sum[2][7]  ;
wire \sum[2][6]  ;
wire \sum[2][5]  ;
wire \sum[2][4]  ;
wire \sum[2][3]  ;
wire \sum[2][2]  ;
wire \sum[2][1]  ;
wire \sum[2][0]  ;
wire \sum[1][23]  ;
wire \sum[1][22]  ;
wire \sum[1][21]  ;
wire \sum[1][20]  ;
wire \sum[1][19]  ;
wire \sum[1][18]  ;
wire \sum[1][17]  ;
wire \sum[1][16]  ;
wire \sum[1][15]  ;
wire \sum[1][14]  ;
wire \sum[1][13]  ;
wire \sum[1][12]  ;
wire \sum[1][11]  ;
wire \sum[1][10]  ;
wire \sum[1][9]  ;
wire \sum[1][8]  ;
wire \sum[1][7]  ;
wire \sum[1][6]  ;
wire \sum[1][5]  ;
wire \sum[1][4]  ;
wire \sum[1][3]  ;
wire \sum[1][2]  ;
wire \sum[1][1]  ;
wire \sum[1][0]  ;
wire \sum[0][23]  ;
wire \sum[0][22]  ;
wire \sum[0][21]  ;
wire \sum[0][20]  ;
wire \sum[0][19]  ;
wire \sum[0][18]  ;
wire \sum[0][17]  ;
wire \sum[0][16]  ;
wire \sum[0][15]  ;
wire \sum[0][14]  ;
wire \sum[0][13]  ;
wire \sum[0][12]  ;
wire \sum[0][11]  ;
wire \sum[0][10]  ;
wire \sum[0][9]  ;
wire \sum[0][8]  ;
wire \sum[0][7]  ;
wire \sum[0][6]  ;
wire \sum[0][5]  ;
wire \sum[0][4]  ;
wire \sum[0][3]  ;
wire \sum[0][2]  ;
wire \sum[0][1]  ;
wire \sum[0][0]  ;
wire n25 ;
wire n38 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire N273 ;
wire N272 ;
wire N271 ;
wire N270 ;
wire N269 ;
wire N268 ;
wire N267 ;
wire N266 ;
wire N265 ;
wire N264 ;
wire N263 ;
wire N262 ;
wire N261 ;
wire N260 ;
wire N259 ;
wire N258 ;
wire N257 ;
wire N256 ;
wire N218 ;
wire N217 ;
wire N216 ;
wire N215 ;
wire N214 ;
wire N213 ;
wire N212 ;
wire N211 ;
wire N210 ;
wire N209 ;
wire N208 ;
wire N207 ;
wire N206 ;
wire N205 ;
wire N204 ;
wire N203 ;
wire N202 ;
wire N201 ;
wire N200 ;
wire N412 ;
wire N411 ;
wire N410 ;
wire N409 ;
wire N408 ;
wire N407 ;
wire N406 ;
wire N405 ;
wire N404 ;
wire N403 ;
wire N402 ;
wire N401 ;
wire N400 ;
wire N399 ;
wire N398 ;
wire N397 ;
wire N396 ;
wire N395 ;
wire N394 ;
wire N393 ;
wire N392 ;
wire N391 ;
wire N390 ;
wire N389 ;
wire N388 ;
wire N387 ;
wire N386 ;
wire N385 ;
wire N384 ;
wire N383 ;
wire N382 ;
wire N381 ;
wire N380 ;
wire N379 ;
wire N378 ;
wire N377 ;
wire N376 ;
wire N375 ;
wire N374 ;
wire N373 ;
wire N372 ;
wire N371 ;
wire N370 ;
wire N369 ;
wire N368 ;
wire N367 ;
wire N366 ;
wire N365 ;
wire N364 ;
wire N363 ;
wire N362 ;
wire N361 ;
wire N360 ;
wire N359 ;
wire N358 ;
wire N357 ;
wire N356 ;
wire N355 ;
wire N354 ;
wire N353 ;
wire N352 ;
wire N351 ;
wire N350 ;
wire N349 ;
wire N348 ;
wire N347 ;
wire N346 ;
wire N345 ;
wire N344 ;
wire N343 ;
wire N342 ;
wire N341 ;
wire N340 ;
wire \add_2_root_add_0_root_add_208_3/carry[23]  ;
wire \add_2_root_add_0_root_add_208_3/carry[22]  ;
wire \add_2_root_add_0_root_add_208_3/carry[21]  ;
wire \add_2_root_add_0_root_add_208_3/carry[20]  ;
wire \add_2_root_add_0_root_add_208_3/carry[19]  ;
wire \add_2_root_add_0_root_add_208_3/carry[18]  ;
wire \add_2_root_add_0_root_add_208_3/carry[17]  ;
wire \add_2_root_add_0_root_add_208_3/carry[16]  ;
wire \add_2_root_add_0_root_add_208_3/carry[15]  ;
wire \add_2_root_add_0_root_add_208_3/carry[14]  ;
wire \add_2_root_add_0_root_add_208_3/carry[13]  ;
wire \add_1_root_add_0_root_add_208_3/carry[7]  ;
wire \add_1_root_add_0_root_add_208_3/carry[8]  ;
wire \add_1_root_add_0_root_add_208_3/carry[9]  ;
wire \add_1_root_add_0_root_add_208_3/carry[10]  ;
wire \add_1_root_add_0_root_add_208_3/carry[11]  ;
wire \add_1_root_add_0_root_add_208_3/carry[12]  ;
wire \add_1_root_add_0_root_add_208_3/carry[13]  ;
wire \add_1_root_add_0_root_add_208_3/carry[14]  ;
wire \add_1_root_add_0_root_add_208_3/carry[15]  ;
wire \add_1_root_add_0_root_add_208_3/carry[16]  ;
wire \add_1_root_add_0_root_add_208_3/carry[17]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n39 ;
wire n40 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire [23:0] s_fracta_i ;
wire [23:0] s_fractb_i ;
wire SYNOPSYS_UNCONNECTED__0 ;
wire SYNOPSYS_UNCONNECTED__1 ;
wire SYNOPSYS_UNCONNECTED__2 ;
wire SYNOPSYS_UNCONNECTED__3 ;
wire SYNOPSYS_UNCONNECTED__4 ;
wire SYNOPSYS_UNCONNECTED__5 ;
wire SYNOPSYS_UNCONNECTED__6 ;
wire SYNOPSYS_UNCONNECTED__7 ;
wire SYNOPSYS_UNCONNECTED__8 ;
wire SYNOPSYS_UNCONNECTED__9 ;
wire SYNOPSYS_UNCONNECTED__10 ;
wire SYNOPSYS_UNCONNECTED__11 ;
wire SYNOPSYS_UNCONNECTED__12 ;
wire SYNOPSYS_UNCONNECTED__13 ;
wire SYNOPSYS_UNCONNECTED__14 ;
wire SYNOPSYS_UNCONNECTED__15 ;
wire SYNOPSYS_UNCONNECTED__16 ;
wire SYNOPSYS_UNCONNECTED__17 ;
wire SYNOPSYS_UNCONNECTED__18 ;
wire SYNOPSYS_UNCONNECTED__19 ;
wire SYNOPSYS_UNCONNECTED__20 ;
wire SYNOPSYS_UNCONNECTED__21 ;
wire SYNOPSYS_UNCONNECTED__22 ;
// instances
  DFFX1 desc375(.D(fracta_i[23:23]),.CLK(clk_i),.Q(s_fracta_i[23:23]));
  DFFX1 desc376(.D(fracta_i[22:22]),.CLK(clk_i),.Q(s_fracta_i[22:22]));
  DFFX1 desc377(.D(fracta_i[21:21]),.CLK(clk_i),.Q(s_fracta_i[21:21]));
  DFFX1 desc378(.D(fracta_i[20:20]),.CLK(clk_i),.Q(s_fracta_i[20:20]));
  DFFX1 desc379(.D(fracta_i[19:19]),.CLK(clk_i),.Q(s_fracta_i[19:19]));
  DFFX1 desc380(.D(fracta_i[18:18]),.CLK(clk_i),.Q(s_fracta_i[18:18]));
  DFFX1 desc381(.D(fracta_i[17:17]),.CLK(clk_i),.Q(s_fracta_i[17:17]));
  DFFX1 desc382(.D(fracta_i[16:16]),.CLK(clk_i),.Q(s_fracta_i[16:16]));
  DFFX1 desc383(.D(fracta_i[15:15]),.CLK(clk_i),.Q(s_fracta_i[15:15]));
  DFFX1 desc384(.D(fracta_i[14:14]),.CLK(clk_i),.Q(s_fracta_i[14:14]));
  DFFX1 desc385(.D(fracta_i[13:13]),.CLK(clk_i),.Q(s_fracta_i[13:13]));
  DFFX1 desc386(.D(fracta_i[12:12]),.CLK(clk_i),.Q(s_fracta_i[12:12]));
  DFFX1 desc387(.D(fracta_i[11:11]),.CLK(clk_i),.Q(s_fracta_i[11:11]));
  DFFX1 desc388(.D(fracta_i[10:10]),.CLK(clk_i),.Q(s_fracta_i[10:10]));
  DFFX1 desc389(.D(fracta_i[9:9]),.CLK(clk_i),.Q(s_fracta_i[9:9]));
  DFFX1 desc390(.D(fracta_i[8:8]),.CLK(clk_i),.Q(s_fracta_i[8:8]));
  DFFX1 desc391(.D(fracta_i[7:7]),.CLK(clk_i),.Q(s_fracta_i[7:7]));
  DFFX1 desc392(.D(fracta_i[6:6]),.CLK(clk_i),.Q(s_fracta_i[6:6]));
  DFFX1 desc393(.D(fracta_i[5:5]),.CLK(clk_i),.Q(s_fracta_i[5:5]));
  DFFX1 desc394(.D(fracta_i[4:4]),.CLK(clk_i),.Q(s_fracta_i[4:4]));
  DFFX1 desc395(.D(fracta_i[3:3]),.CLK(clk_i),.Q(s_fracta_i[3:3]));
  DFFX1 desc396(.D(fracta_i[2:2]),.CLK(clk_i),.Q(s_fracta_i[2:2]));
  DFFX1 desc397(.D(fracta_i[1:1]),.CLK(clk_i),.Q(s_fracta_i[1:1]));
  DFFX1 desc398(.D(fracta_i[0:0]),.CLK(clk_i),.Q(s_fracta_i[0:0]));
  DFFX1 desc399(.D(fractb_i[23:23]),.CLK(clk_i),.Q(s_fractb_i[23:23]));
  DFFX1 desc400(.D(fractb_i[22:22]),.CLK(clk_i),.Q(s_fractb_i[22:22]));
  DFFX1 desc401(.D(fractb_i[21:21]),.CLK(clk_i),.Q(s_fractb_i[21:21]));
  DFFX1 desc402(.D(fractb_i[20:20]),.CLK(clk_i),.Q(s_fractb_i[20:20]));
  DFFX1 desc403(.D(fractb_i[19:19]),.CLK(clk_i),.Q(s_fractb_i[19:19]));
  DFFX1 desc404(.D(fractb_i[18:18]),.CLK(clk_i),.Q(s_fractb_i[18:18]));
  DFFX1 desc405(.D(fractb_i[17:17]),.CLK(clk_i),.Q(s_fractb_i[17:17]));
  DFFX1 desc406(.D(fractb_i[16:16]),.CLK(clk_i),.Q(s_fractb_i[16:16]));
  DFFX1 desc407(.D(fractb_i[15:15]),.CLK(clk_i),.Q(s_fractb_i[15:15]));
  DFFX1 desc408(.D(fractb_i[14:14]),.CLK(clk_i),.Q(s_fractb_i[14:14]));
  DFFX1 desc409(.D(fractb_i[13:13]),.CLK(clk_i),.Q(s_fractb_i[13:13]));
  DFFX1 desc410(.D(fractb_i[12:12]),.CLK(clk_i),.Q(s_fractb_i[12:12]));
  DFFX1 desc411(.D(fractb_i[11:11]),.CLK(clk_i),.Q(s_fractb_i[11:11]));
  DFFX1 desc412(.D(fractb_i[10:10]),.CLK(clk_i),.Q(s_fractb_i[10:10]));
  DFFX1 desc413(.D(fractb_i[9:9]),.CLK(clk_i),.Q(s_fractb_i[9:9]));
  DFFX1 desc414(.D(fractb_i[8:8]),.CLK(clk_i),.Q(s_fractb_i[8:8]));
  DFFX1 desc415(.D(fractb_i[7:7]),.CLK(clk_i),.Q(s_fractb_i[7:7]));
  DFFX1 desc416(.D(fractb_i[6:6]),.CLK(clk_i),.Q(s_fractb_i[6:6]));
  DFFX1 desc417(.D(fractb_i[5:5]),.CLK(clk_i),.Q(s_fractb_i[5:5]));
  DFFX1 desc418(.D(fractb_i[4:4]),.CLK(clk_i),.Q(s_fractb_i[4:4]));
  DFFX1 desc419(.D(fractb_i[3:3]),.CLK(clk_i),.Q(s_fractb_i[3:3]));
  DFFX1 desc420(.D(fractb_i[2:2]),.CLK(clk_i),.Q(s_fractb_i[2:2]));
  DFFX1 desc421(.D(fractb_i[1:1]),.CLK(clk_i),.Q(s_fractb_i[1:1]));
  DFFX1 desc422(.D(fractb_i[0:0]),.CLK(clk_i),.Q(s_fractb_i[0:0]));
  DFFX1 s_signa_i_reg(.D(signa_i),.CLK(clk_i),.Q(s_signa_i));
  DFFX1 s_signb_i_reg(.D(signb_i),.CLK(clk_i),.Q(s_signb_i));
  DFFX1 s_start_i_reg(.D(start_i),.CLK(clk_i),.Q(s_start_i),.QN(n25));
  DFFX1 desc423(.D(n352),.CLK(clk_i),.Q(N25),.QN(n41));
  DFFX1 s_state_reg(.D(n350),.CLK(clk_i),.Q(s_state));
  DFFX1 s_ready_o_reg(.D(n349),.CLK(clk_i),.Q(ready_o));
  DFFX1 desc424(.D(n348),.CLK(clk_i),.Q(N26));
  DFFX1 desc425(.D(n351),.CLK(clk_i),.Q(\count[2] ),.QN(n38));
  DFFX1 desc426(.D(n347),.CLK(clk_i),.Q(\prod2[3][3][11] ));
  DFFX1 desc427(.D(n346),.CLK(clk_i),.Q(\prod2[3][3][10] ));
  DFFX1 desc428(.D(n345),.CLK(clk_i),.Q(\prod2[3][3][9] ));
  DFFX1 desc429(.D(n344),.CLK(clk_i),.Q(\prod2[3][3][8] ));
  DFFX1 desc430(.D(n343),.CLK(clk_i),.Q(\prod2[3][3][7] ));
  DFFX1 desc431(.D(n342),.CLK(clk_i),.Q(\prod2[3][3][6] ));
  DFFX1 desc432(.D(n341),.CLK(clk_i),.Q(\prod2[3][3][5] ));
  DFFX1 desc433(.D(n340),.CLK(clk_i),.Q(\prod2[3][3][4] ));
  DFFX1 desc434(.D(n339),.CLK(clk_i),.Q(\prod2[3][3][3] ));
  DFFX1 desc435(.D(n338),.CLK(clk_i),.Q(\prod2[3][3][2] ));
  DFFX1 desc436(.D(n337),.CLK(clk_i),.Q(\prod2[3][3][1] ));
  DFFX1 desc437(.D(n336),.CLK(clk_i),.Q(\prod2[3][3][0] ));
  DFFX1 desc438(.D(n335),.CLK(clk_i),.Q(\prod2[3][2][17] ));
  DFFX1 desc439(.D(n334),.CLK(clk_i),.Q(\prod2[3][2][16] ));
  DFFX1 desc440(.D(n333),.CLK(clk_i),.Q(\prod2[3][2][15] ));
  DFFX1 desc441(.D(n332),.CLK(clk_i),.Q(\prod2[3][2][14] ));
  DFFX1 desc442(.D(n331),.CLK(clk_i),.Q(\prod2[3][2][13] ));
  DFFX1 desc443(.D(n330),.CLK(clk_i),.Q(\prod2[3][2][12] ));
  DFFX1 desc444(.D(n329),.CLK(clk_i),.Q(\prod2[3][2][11] ));
  DFFX1 desc445(.D(n328),.CLK(clk_i),.Q(\prod2[3][2][10] ));
  DFFX1 desc446(.D(n327),.CLK(clk_i),.Q(\prod2[3][2][9] ));
  DFFX1 desc447(.D(n326),.CLK(clk_i),.Q(\prod2[3][2][8] ));
  DFFX1 desc448(.D(n325),.CLK(clk_i),.Q(\prod2[3][2][7] ));
  DFFX1 desc449(.D(n324),.CLK(clk_i),.Q(\prod2[3][2][6] ));
  DFFX1 desc450(.D(n323),.CLK(clk_i),.Q(\prod2[3][1][17] ));
  DFFX1 desc451(.D(n322),.CLK(clk_i),.Q(\prod2[3][1][16] ));
  DFFX1 desc452(.D(n321),.CLK(clk_i),.Q(\prod2[3][1][15] ));
  DFFX1 desc453(.D(n320),.CLK(clk_i),.Q(\prod2[3][1][14] ));
  DFFX1 desc454(.D(n319),.CLK(clk_i),.Q(\prod2[3][1][13] ));
  DFFX1 desc455(.D(n318),.CLK(clk_i),.Q(\prod2[3][1][12] ));
  DFFX1 desc456(.D(n317),.CLK(clk_i),.Q(\prod2[3][1][11] ));
  DFFX1 desc457(.D(n316),.CLK(clk_i),.Q(\prod2[3][1][10] ));
  DFFX1 desc458(.D(n315),.CLK(clk_i),.Q(\prod2[3][1][9] ));
  DFFX1 desc459(.D(n314),.CLK(clk_i),.Q(\prod2[3][1][8] ));
  DFFX1 desc460(.D(n313),.CLK(clk_i),.Q(\prod2[3][1][7] ));
  DFFX1 desc461(.D(n312),.CLK(clk_i),.Q(\prod2[3][1][6] ));
  DFFX1 desc462(.D(n311),.CLK(clk_i),.Q(\prod2[3][0][23] ));
  DFFX1 desc463(.D(n310),.CLK(clk_i),.Q(\prod2[3][0][22] ));
  DFFX1 desc464(.D(n309),.CLK(clk_i),.Q(\prod2[3][0][21] ));
  DFFX1 desc465(.D(n308),.CLK(clk_i),.Q(\prod2[3][0][20] ));
  DFFX1 desc466(.D(n307),.CLK(clk_i),.Q(\prod2[3][0][19] ));
  DFFX1 desc467(.D(n306),.CLK(clk_i),.Q(\prod2[3][0][18] ));
  DFFX1 desc468(.D(n305),.CLK(clk_i),.Q(\prod2[3][0][17] ));
  DFFX1 desc469(.D(n304),.CLK(clk_i),.Q(\prod2[3][0][16] ));
  DFFX1 desc470(.D(n303),.CLK(clk_i),.Q(\prod2[3][0][15] ));
  DFFX1 desc471(.D(n302),.CLK(clk_i),.Q(\prod2[3][0][14] ));
  DFFX1 desc472(.D(n301),.CLK(clk_i),.Q(\prod2[3][0][13] ));
  DFFX1 desc473(.D(n300),.CLK(clk_i),.Q(\prod2[3][0][12] ));
  DFFX1 desc474(.D(n299),.CLK(clk_i),.Q(\prod2[2][3][11] ));
  DFFX1 desc475(.D(n298),.CLK(clk_i),.Q(\prod2[2][3][10] ));
  DFFX1 desc476(.D(n297),.CLK(clk_i),.Q(\prod2[2][3][9] ));
  DFFX1 desc477(.D(n296),.CLK(clk_i),.Q(\prod2[2][3][8] ));
  DFFX1 desc478(.D(n295),.CLK(clk_i),.Q(\prod2[2][3][7] ));
  DFFX1 desc479(.D(n294),.CLK(clk_i),.Q(\prod2[2][3][6] ));
  DFFX1 desc480(.D(n293),.CLK(clk_i),.Q(\prod2[2][3][5] ));
  DFFX1 desc481(.D(n292),.CLK(clk_i),.Q(\prod2[2][3][4] ));
  DFFX1 desc482(.D(n291),.CLK(clk_i),.Q(\prod2[2][3][3] ));
  DFFX1 desc483(.D(n290),.CLK(clk_i),.Q(\prod2[2][3][2] ));
  DFFX1 desc484(.D(n289),.CLK(clk_i),.Q(\prod2[2][3][1] ));
  DFFX1 desc485(.D(n288),.CLK(clk_i),.Q(\prod2[2][3][0] ));
  DFFX1 desc486(.D(n287),.CLK(clk_i),.Q(\prod2[2][2][17] ));
  DFFX1 desc487(.D(n286),.CLK(clk_i),.Q(\prod2[2][2][16] ));
  DFFX1 desc488(.D(n285),.CLK(clk_i),.Q(\prod2[2][2][15] ));
  DFFX1 desc489(.D(n284),.CLK(clk_i),.Q(\prod2[2][2][14] ));
  DFFX1 desc490(.D(n283),.CLK(clk_i),.Q(\prod2[2][2][13] ));
  DFFX1 desc491(.D(n282),.CLK(clk_i),.Q(\prod2[2][2][12] ));
  DFFX1 desc492(.D(n281),.CLK(clk_i),.Q(\prod2[2][2][11] ));
  DFFX1 desc493(.D(n280),.CLK(clk_i),.Q(\prod2[2][2][10] ));
  DFFX1 desc494(.D(n279),.CLK(clk_i),.Q(\prod2[2][2][9] ));
  DFFX1 desc495(.D(n278),.CLK(clk_i),.Q(\prod2[2][2][8] ));
  DFFX1 desc496(.D(n277),.CLK(clk_i),.Q(\prod2[2][2][7] ));
  DFFX1 desc497(.D(n276),.CLK(clk_i),.Q(\prod2[2][2][6] ));
  DFFX1 desc498(.D(n275),.CLK(clk_i),.Q(\prod2[2][1][17] ));
  DFFX1 desc499(.D(n274),.CLK(clk_i),.Q(\prod2[2][1][16] ));
  DFFX1 desc500(.D(n273),.CLK(clk_i),.Q(\prod2[2][1][15] ));
  DFFX1 desc501(.D(n272),.CLK(clk_i),.Q(\prod2[2][1][14] ));
  DFFX1 desc502(.D(n271),.CLK(clk_i),.Q(\prod2[2][1][13] ));
  DFFX1 desc503(.D(n270),.CLK(clk_i),.Q(\prod2[2][1][12] ));
  DFFX1 desc504(.D(n269),.CLK(clk_i),.Q(\prod2[2][1][11] ));
  DFFX1 desc505(.D(n268),.CLK(clk_i),.Q(\prod2[2][1][10] ));
  DFFX1 desc506(.D(n267),.CLK(clk_i),.Q(\prod2[2][1][9] ));
  DFFX1 desc507(.D(n266),.CLK(clk_i),.Q(\prod2[2][1][8] ));
  DFFX1 desc508(.D(n265),.CLK(clk_i),.Q(\prod2[2][1][7] ));
  DFFX1 desc509(.D(n264),.CLK(clk_i),.Q(\prod2[2][1][6] ));
  DFFX1 desc510(.D(n263),.CLK(clk_i),.Q(\prod2[2][0][23] ));
  DFFX1 desc511(.D(n262),.CLK(clk_i),.Q(\prod2[2][0][22] ));
  DFFX1 desc512(.D(n261),.CLK(clk_i),.Q(\prod2[2][0][21] ));
  DFFX1 desc513(.D(n260),.CLK(clk_i),.Q(\prod2[2][0][20] ));
  DFFX1 desc514(.D(n259),.CLK(clk_i),.Q(\prod2[2][0][19] ));
  DFFX1 desc515(.D(n258),.CLK(clk_i),.Q(\prod2[2][0][18] ));
  DFFX1 desc516(.D(n257),.CLK(clk_i),.Q(\prod2[2][0][17] ));
  DFFX1 desc517(.D(n256),.CLK(clk_i),.Q(\prod2[2][0][16] ));
  DFFX1 desc518(.D(n255),.CLK(clk_i),.Q(\prod2[2][0][15] ));
  DFFX1 desc519(.D(n254),.CLK(clk_i),.Q(\prod2[2][0][14] ));
  DFFX1 desc520(.D(n253),.CLK(clk_i),.Q(\prod2[2][0][13] ));
  DFFX1 desc521(.D(n252),.CLK(clk_i),.Q(\prod2[2][0][12] ));
  DFFX1 desc522(.D(n251),.CLK(clk_i),.Q(\prod2[1][3][11] ));
  DFFX1 desc523(.D(n250),.CLK(clk_i),.Q(\prod2[1][3][10] ));
  DFFX1 desc524(.D(n249),.CLK(clk_i),.Q(\prod2[1][3][9] ));
  DFFX1 desc525(.D(n248),.CLK(clk_i),.Q(\prod2[1][3][8] ));
  DFFX1 desc526(.D(n247),.CLK(clk_i),.Q(\prod2[1][3][7] ));
  DFFX1 desc527(.D(n246),.CLK(clk_i),.Q(\prod2[1][3][6] ));
  DFFX1 desc528(.D(n245),.CLK(clk_i),.Q(\prod2[1][3][5] ));
  DFFX1 desc529(.D(n244),.CLK(clk_i),.Q(\prod2[1][3][4] ));
  DFFX1 desc530(.D(n243),.CLK(clk_i),.Q(\prod2[1][3][3] ));
  DFFX1 desc531(.D(n242),.CLK(clk_i),.Q(\prod2[1][3][2] ));
  DFFX1 desc532(.D(n241),.CLK(clk_i),.Q(\prod2[1][3][1] ));
  DFFX1 desc533(.D(n240),.CLK(clk_i),.Q(\prod2[1][3][0] ));
  DFFX1 desc534(.D(n239),.CLK(clk_i),.Q(\prod2[1][2][17] ));
  DFFX1 desc535(.D(n238),.CLK(clk_i),.Q(\prod2[1][2][16] ));
  DFFX1 desc536(.D(n237),.CLK(clk_i),.Q(\prod2[1][2][15] ));
  DFFX1 desc537(.D(n236),.CLK(clk_i),.Q(\prod2[1][2][14] ));
  DFFX1 desc538(.D(n235),.CLK(clk_i),.Q(\prod2[1][2][13] ));
  DFFX1 desc539(.D(n234),.CLK(clk_i),.Q(\prod2[1][2][12] ));
  DFFX1 desc540(.D(n233),.CLK(clk_i),.Q(\prod2[1][2][11] ));
  DFFX1 desc541(.D(n232),.CLK(clk_i),.Q(\prod2[1][2][10] ));
  DFFX1 desc542(.D(n231),.CLK(clk_i),.Q(\prod2[1][2][9] ));
  DFFX1 desc543(.D(n230),.CLK(clk_i),.Q(\prod2[1][2][8] ));
  DFFX1 desc544(.D(n229),.CLK(clk_i),.Q(\prod2[1][2][7] ));
  DFFX1 desc545(.D(n228),.CLK(clk_i),.Q(\prod2[1][2][6] ));
  DFFX1 desc546(.D(n227),.CLK(clk_i),.Q(\prod2[1][1][17] ));
  DFFX1 desc547(.D(n226),.CLK(clk_i),.Q(\prod2[1][1][16] ));
  DFFX1 desc548(.D(n225),.CLK(clk_i),.Q(\prod2[1][1][15] ));
  DFFX1 desc549(.D(n224),.CLK(clk_i),.Q(\prod2[1][1][14] ));
  DFFX1 desc550(.D(n223),.CLK(clk_i),.Q(\prod2[1][1][13] ));
  DFFX1 desc551(.D(n222),.CLK(clk_i),.Q(\prod2[1][1][12] ));
  DFFX1 desc552(.D(n221),.CLK(clk_i),.Q(\prod2[1][1][11] ));
  DFFX1 desc553(.D(n220),.CLK(clk_i),.Q(\prod2[1][1][10] ));
  DFFX1 desc554(.D(n219),.CLK(clk_i),.Q(\prod2[1][1][9] ));
  DFFX1 desc555(.D(n218),.CLK(clk_i),.Q(\prod2[1][1][8] ));
  DFFX1 desc556(.D(n217),.CLK(clk_i),.Q(\prod2[1][1][7] ));
  DFFX1 desc557(.D(n216),.CLK(clk_i),.Q(\prod2[1][1][6] ));
  DFFX1 desc558(.D(n215),.CLK(clk_i),.Q(\prod2[1][0][23] ));
  DFFX1 desc559(.D(n214),.CLK(clk_i),.Q(\prod2[1][0][22] ));
  DFFX1 desc560(.D(n213),.CLK(clk_i),.Q(\prod2[1][0][21] ));
  DFFX1 desc561(.D(n212),.CLK(clk_i),.Q(\prod2[1][0][20] ));
  DFFX1 desc562(.D(n211),.CLK(clk_i),.Q(\prod2[1][0][19] ));
  DFFX1 desc563(.D(n210),.CLK(clk_i),.Q(\prod2[1][0][18] ));
  DFFX1 desc564(.D(n209),.CLK(clk_i),.Q(\prod2[1][0][17] ));
  DFFX1 desc565(.D(n208),.CLK(clk_i),.Q(\prod2[1][0][16] ));
  DFFX1 desc566(.D(n207),.CLK(clk_i),.Q(\prod2[1][0][15] ));
  DFFX1 desc567(.D(n206),.CLK(clk_i),.Q(\prod2[1][0][14] ));
  DFFX1 desc568(.D(n205),.CLK(clk_i),.Q(\prod2[1][0][13] ));
  DFFX1 desc569(.D(n204),.CLK(clk_i),.Q(\prod2[1][0][12] ));
  DFFX1 desc570(.D(n203),.CLK(clk_i),.Q(\prod2[0][3][11] ));
  DFFX1 desc571(.D(n202),.CLK(clk_i),.Q(\prod2[0][3][10] ));
  DFFX1 desc572(.D(n201),.CLK(clk_i),.Q(\prod2[0][3][9] ));
  DFFX1 desc573(.D(n200),.CLK(clk_i),.Q(\prod2[0][3][8] ));
  DFFX1 desc574(.D(n199),.CLK(clk_i),.Q(\prod2[0][3][7] ));
  DFFX1 desc575(.D(n198),.CLK(clk_i),.Q(\prod2[0][3][6] ));
  DFFX1 desc576(.D(n197),.CLK(clk_i),.Q(\prod2[0][3][5] ));
  DFFX1 desc577(.D(n196),.CLK(clk_i),.Q(\prod2[0][3][4] ));
  DFFX1 desc578(.D(n195),.CLK(clk_i),.Q(\prod2[0][3][3] ));
  DFFX1 desc579(.D(n194),.CLK(clk_i),.Q(\prod2[0][3][2] ));
  DFFX1 desc580(.D(n193),.CLK(clk_i),.Q(\prod2[0][3][1] ));
  DFFX1 desc581(.D(n192),.CLK(clk_i),.Q(\prod2[0][3][0] ));
  DFFX1 desc582(.D(n191),.CLK(clk_i),.Q(\prod2[0][2][17] ));
  DFFX1 desc583(.D(n190),.CLK(clk_i),.Q(\prod2[0][2][16] ));
  DFFX1 desc584(.D(n189),.CLK(clk_i),.Q(\prod2[0][2][15] ));
  DFFX1 desc585(.D(n188),.CLK(clk_i),.Q(\prod2[0][2][14] ));
  DFFX1 desc586(.D(n187),.CLK(clk_i),.Q(\prod2[0][2][13] ));
  DFFX1 desc587(.D(n186),.CLK(clk_i),.Q(\prod2[0][2][12] ));
  DFFX1 desc588(.D(n185),.CLK(clk_i),.Q(\prod2[0][2][11] ));
  DFFX1 desc589(.D(n184),.CLK(clk_i),.Q(\prod2[0][2][10] ));
  DFFX1 desc590(.D(n183),.CLK(clk_i),.Q(\prod2[0][2][9] ));
  DFFX1 desc591(.D(n182),.CLK(clk_i),.Q(\prod2[0][2][8] ));
  DFFX1 desc592(.D(n181),.CLK(clk_i),.Q(\prod2[0][2][7] ));
  DFFX1 desc593(.D(n180),.CLK(clk_i),.Q(\prod2[0][2][6] ));
  DFFX1 desc594(.D(n179),.CLK(clk_i),.Q(\prod2[0][1][17] ));
  DFFX1 desc595(.D(n178),.CLK(clk_i),.Q(\prod2[0][1][16] ));
  DFFX1 desc596(.D(n177),.CLK(clk_i),.Q(\prod2[0][1][15] ));
  DFFX1 desc597(.D(n176),.CLK(clk_i),.Q(\prod2[0][1][14] ));
  DFFX1 desc598(.D(n175),.CLK(clk_i),.Q(\prod2[0][1][13] ));
  DFFX1 desc599(.D(n174),.CLK(clk_i),.Q(\prod2[0][1][12] ));
  DFFX1 desc600(.D(n173),.CLK(clk_i),.Q(\prod2[0][1][11] ));
  DFFX1 desc601(.D(n172),.CLK(clk_i),.Q(\prod2[0][1][10] ));
  DFFX1 desc602(.D(n171),.CLK(clk_i),.Q(\prod2[0][1][9] ));
  DFFX1 desc603(.D(n170),.CLK(clk_i),.Q(\prod2[0][1][8] ));
  DFFX1 desc604(.D(n169),.CLK(clk_i),.Q(\prod2[0][1][7] ));
  DFFX1 desc605(.D(n168),.CLK(clk_i),.Q(\prod2[0][1][6] ));
  DFFX1 desc606(.D(n167),.CLK(clk_i),.Q(\prod2[0][0][23] ));
  DFFX1 desc607(.D(n166),.CLK(clk_i),.Q(\prod2[0][0][22] ));
  DFFX1 desc608(.D(n165),.CLK(clk_i),.Q(\prod2[0][0][21] ));
  DFFX1 desc609(.D(n164),.CLK(clk_i),.Q(\prod2[0][0][20] ));
  DFFX1 desc610(.D(n163),.CLK(clk_i),.Q(\prod2[0][0][19] ));
  DFFX1 desc611(.D(n162),.CLK(clk_i),.Q(\prod2[0][0][18] ));
  DFFX1 desc612(.D(n161),.CLK(clk_i),.Q(\prod2[0][0][17] ));
  DFFX1 desc613(.D(n160),.CLK(clk_i),.Q(\prod2[0][0][16] ));
  DFFX1 desc614(.D(n159),.CLK(clk_i),.Q(\prod2[0][0][15] ));
  DFFX1 desc615(.D(n158),.CLK(clk_i),.Q(\prod2[0][0][14] ));
  DFFX1 desc616(.D(n157),.CLK(clk_i),.Q(\prod2[0][0][13] ));
  DFFX1 desc617(.D(n156),.CLK(clk_i),.Q(\prod2[0][0][12] ));
  DFFX1 desc618(.D(n155),.CLK(clk_i),.Q(\sum[3][23] ));
  DFFX1 desc619(.D(n154),.CLK(clk_i),.Q(\sum[3][22] ));
  DFFX1 desc620(.D(n153),.CLK(clk_i),.Q(\sum[3][21] ));
  DFFX1 desc621(.D(n152),.CLK(clk_i),.Q(\sum[3][20] ));
  DFFX1 desc622(.D(n151),.CLK(clk_i),.Q(\sum[3][19] ));
  DFFX1 desc623(.D(n150),.CLK(clk_i),.Q(\sum[3][18] ));
  DFFX1 desc624(.D(n149),.CLK(clk_i),.Q(\sum[3][17] ));
  DFFX1 desc625(.D(n148),.CLK(clk_i),.Q(\sum[3][16] ));
  DFFX1 desc626(.D(n147),.CLK(clk_i),.Q(\sum[3][15] ));
  DFFX1 desc627(.D(n146),.CLK(clk_i),.Q(\sum[3][14] ));
  DFFX1 desc628(.D(n145),.CLK(clk_i),.Q(\sum[3][13] ));
  DFFX1 desc629(.D(n144),.CLK(clk_i),.Q(\sum[3][12] ));
  DFFX1 desc630(.D(n143),.CLK(clk_i),.Q(\sum[3][11] ));
  DFFX1 desc631(.D(n142),.CLK(clk_i),.Q(\sum[3][10] ));
  DFFX1 desc632(.D(n141),.CLK(clk_i),.Q(\sum[3][9] ));
  DFFX1 desc633(.D(n140),.CLK(clk_i),.Q(\sum[3][8] ));
  DFFX1 desc634(.D(n139),.CLK(clk_i),.Q(\sum[3][7] ));
  DFFX1 desc635(.D(n138),.CLK(clk_i),.Q(\sum[3][6] ));
  DFFX1 desc636(.D(n137),.CLK(clk_i),.Q(\sum[3][5] ));
  DFFX1 desc637(.D(n136),.CLK(clk_i),.Q(\sum[3][4] ));
  DFFX1 desc638(.D(n135),.CLK(clk_i),.Q(\sum[3][3] ));
  DFFX1 desc639(.D(n134),.CLK(clk_i),.Q(\sum[3][2] ));
  DFFX1 desc640(.D(n133),.CLK(clk_i),.Q(\sum[3][1] ));
  DFFX1 desc641(.D(n132),.CLK(clk_i),.Q(\sum[3][0] ));
  DFFX1 desc642(.D(n131),.CLK(clk_i),.Q(\sum[2][23] ));
  DFFX1 desc643(.D(n130),.CLK(clk_i),.Q(\sum[2][22] ));
  DFFX1 desc644(.D(n129),.CLK(clk_i),.Q(\sum[2][21] ));
  DFFX1 desc645(.D(n128),.CLK(clk_i),.Q(\sum[2][20] ));
  DFFX1 desc646(.D(n127),.CLK(clk_i),.Q(\sum[2][19] ));
  DFFX1 desc647(.D(n126),.CLK(clk_i),.Q(\sum[2][18] ));
  DFFX1 desc648(.D(n125),.CLK(clk_i),.Q(\sum[2][17] ));
  DFFX1 desc649(.D(n124),.CLK(clk_i),.Q(\sum[2][16] ));
  DFFX1 desc650(.D(n123),.CLK(clk_i),.Q(\sum[2][15] ));
  DFFX1 desc651(.D(n122),.CLK(clk_i),.Q(\sum[2][14] ));
  DFFX1 desc652(.D(n121),.CLK(clk_i),.Q(\sum[2][13] ));
  DFFX1 desc653(.D(n120),.CLK(clk_i),.Q(\sum[2][12] ));
  DFFX1 desc654(.D(n119),.CLK(clk_i),.Q(\sum[2][11] ));
  DFFX1 desc655(.D(n118),.CLK(clk_i),.Q(\sum[2][10] ));
  DFFX1 desc656(.D(n117),.CLK(clk_i),.Q(\sum[2][9] ));
  DFFX1 desc657(.D(n116),.CLK(clk_i),.Q(\sum[2][8] ));
  DFFX1 desc658(.D(n115),.CLK(clk_i),.Q(\sum[2][7] ));
  DFFX1 desc659(.D(n114),.CLK(clk_i),.Q(\sum[2][6] ));
  DFFX1 desc660(.D(n113),.CLK(clk_i),.Q(\sum[2][5] ));
  DFFX1 desc661(.D(n112),.CLK(clk_i),.Q(\sum[2][4] ));
  DFFX1 desc662(.D(n111),.CLK(clk_i),.Q(\sum[2][3] ));
  DFFX1 desc663(.D(n110),.CLK(clk_i),.Q(\sum[2][2] ));
  DFFX1 desc664(.D(n109),.CLK(clk_i),.Q(\sum[2][1] ));
  DFFX1 desc665(.D(n108),.CLK(clk_i),.Q(\sum[2][0] ));
  DFFX1 desc666(.D(n107),.CLK(clk_i),.Q(\sum[1][23] ));
  DFFX1 desc667(.D(n106),.CLK(clk_i),.Q(\sum[1][22] ));
  DFFX1 desc668(.D(n105),.CLK(clk_i),.Q(\sum[1][21] ));
  DFFX1 desc669(.D(n104),.CLK(clk_i),.Q(\sum[1][20] ));
  DFFX1 desc670(.D(n103),.CLK(clk_i),.Q(\sum[1][19] ));
  DFFX1 desc671(.D(n102),.CLK(clk_i),.Q(\sum[1][18] ));
  DFFX1 desc672(.D(n101),.CLK(clk_i),.Q(\sum[1][17] ));
  DFFX1 desc673(.D(n100),.CLK(clk_i),.Q(\sum[1][16] ));
  DFFX1 desc674(.D(n99),.CLK(clk_i),.Q(\sum[1][15] ));
  DFFX1 desc675(.D(n98),.CLK(clk_i),.Q(\sum[1][14] ));
  DFFX1 desc676(.D(n97),.CLK(clk_i),.Q(\sum[1][13] ));
  DFFX1 desc677(.D(n96),.CLK(clk_i),.Q(\sum[1][12] ));
  DFFX1 desc678(.D(n95),.CLK(clk_i),.Q(\sum[1][11] ));
  DFFX1 desc679(.D(n94),.CLK(clk_i),.Q(\sum[1][10] ));
  DFFX1 desc680(.D(n93),.CLK(clk_i),.Q(\sum[1][9] ));
  DFFX1 desc681(.D(n92),.CLK(clk_i),.Q(\sum[1][8] ));
  DFFX1 desc682(.D(n91),.CLK(clk_i),.Q(\sum[1][7] ));
  DFFX1 desc683(.D(n90),.CLK(clk_i),.Q(\sum[1][6] ));
  DFFX1 desc684(.D(n89),.CLK(clk_i),.Q(\sum[1][5] ));
  DFFX1 desc685(.D(n88),.CLK(clk_i),.Q(\sum[1][4] ));
  DFFX1 desc686(.D(n87),.CLK(clk_i),.Q(\sum[1][3] ));
  DFFX1 desc687(.D(n86),.CLK(clk_i),.Q(\sum[1][2] ));
  DFFX1 desc688(.D(n85),.CLK(clk_i),.Q(\sum[1][1] ));
  DFFX1 desc689(.D(n84),.CLK(clk_i),.Q(\sum[1][0] ));
  DFFX1 desc690(.D(n83),.CLK(clk_i),.Q(\sum[0][23] ));
  DFFX1 desc691(.D(n82),.CLK(clk_i),.Q(\sum[0][22] ));
  DFFX1 desc692(.D(n81),.CLK(clk_i),.Q(\sum[0][21] ));
  DFFX1 desc693(.D(n80),.CLK(clk_i),.Q(\sum[0][20] ));
  DFFX1 desc694(.D(n79),.CLK(clk_i),.Q(\sum[0][19] ));
  DFFX1 desc695(.D(n78),.CLK(clk_i),.Q(\sum[0][18] ));
  DFFX1 desc696(.D(n77),.CLK(clk_i),.Q(\sum[0][17] ));
  DFFX1 desc697(.D(n76),.CLK(clk_i),.Q(\sum[0][16] ));
  DFFX1 desc698(.D(n75),.CLK(clk_i),.Q(\sum[0][15] ));
  DFFX1 desc699(.D(n74),.CLK(clk_i),.Q(\sum[0][14] ));
  DFFX1 desc700(.D(n73),.CLK(clk_i),.Q(\sum[0][13] ));
  DFFX1 desc701(.D(n72),.CLK(clk_i),.Q(\sum[0][12] ));
  DFFX1 desc702(.D(n71),.CLK(clk_i),.Q(\sum[0][11] ));
  DFFX1 desc703(.D(n70),.CLK(clk_i),.Q(\sum[0][10] ));
  DFFX1 desc704(.D(n69),.CLK(clk_i),.Q(\sum[0][9] ));
  DFFX1 desc705(.D(n68),.CLK(clk_i),.Q(\sum[0][8] ));
  DFFX1 desc706(.D(n67),.CLK(clk_i),.Q(\sum[0][7] ));
  DFFX1 desc707(.D(n66),.CLK(clk_i),.Q(\sum[0][6] ));
  DFFX1 desc708(.D(n65),.CLK(clk_i),.Q(\sum[0][5] ));
  DFFX1 desc709(.D(n64),.CLK(clk_i),.Q(\sum[0][4] ));
  DFFX1 desc710(.D(n63),.CLK(clk_i),.Q(\sum[0][3] ));
  DFFX1 desc711(.D(n62),.CLK(clk_i),.Q(\sum[0][2] ));
  DFFX1 desc712(.D(n61),.CLK(clk_i),.Q(\sum[0][1] ));
  DFFX1 desc713(.D(n60),.CLK(clk_i),.Q(\sum[0][0] ));
  XOR2X1 U225(.IN1(s_signb_i),.IN2(s_signa_i),.Q(sign_o));
  AO22X1 U226(.IN1(N300),.IN2(n33),.IN3(\sum[0][0] ),.IN4(n42),.Q(n60));
  AO22X1 U227(.IN1(N301),.IN2(n32),.IN3(\sum[0][1] ),.IN4(n42),.Q(n61));
  AO22X1 U228(.IN1(N302),.IN2(n33),.IN3(\sum[0][2] ),.IN4(n42),.Q(n62));
  AO22X1 U229(.IN1(N303),.IN2(n32),.IN3(\sum[0][3] ),.IN4(n42),.Q(n63));
  AO22X1 U230(.IN1(N304),.IN2(n33),.IN3(\sum[0][4] ),.IN4(n42),.Q(n64));
  AO22X1 U231(.IN1(N305),.IN2(n32),.IN3(\sum[0][5] ),.IN4(n42),.Q(n65));
  AO22X1 U232(.IN1(N306),.IN2(n32),.IN3(\sum[0][6] ),.IN4(n42),.Q(n66));
  AO22X1 U233(.IN1(N307),.IN2(n32),.IN3(\sum[0][7] ),.IN4(n42),.Q(n67));
  AO22X1 U234(.IN1(N308),.IN2(n32),.IN3(\sum[0][8] ),.IN4(n42),.Q(n68));
  AO22X1 U235(.IN1(N309),.IN2(n32),.IN3(\sum[0][9] ),.IN4(n42),.Q(n69));
  AO22X1 U236(.IN1(N310),.IN2(n32),.IN3(\sum[0][10] ),.IN4(n42),.Q(n70));
  AO22X1 U237(.IN1(N311),.IN2(n32),.IN3(\sum[0][11] ),.IN4(n42),.Q(n71));
  AO22X1 U238(.IN1(N312),.IN2(n33),.IN3(\sum[0][12] ),.IN4(n31),.Q(n72));
  AO22X1 U239(.IN1(N313),.IN2(n33),.IN3(\sum[0][13] ),.IN4(n31),.Q(n73));
  AO22X1 U240(.IN1(N314),.IN2(n33),.IN3(\sum[0][14] ),.IN4(n31),.Q(n74));
  AO22X1 U241(.IN1(N315),.IN2(n33),.IN3(\sum[0][15] ),.IN4(n31),.Q(n75));
  AO22X1 U242(.IN1(N316),.IN2(n33),.IN3(\sum[0][16] ),.IN4(n31),.Q(n76));
  AO22X1 U243(.IN1(N317),.IN2(n33),.IN3(\sum[0][17] ),.IN4(n31),.Q(n77));
  AO22X1 U244(.IN1(N318),.IN2(n33),.IN3(\sum[0][18] ),.IN4(n31),.Q(n78));
  AO22X1 U245(.IN1(N319),.IN2(n32),.IN3(\sum[0][19] ),.IN4(n31),.Q(n79));
  AO22X1 U246(.IN1(N320),.IN2(n33),.IN3(\sum[0][20] ),.IN4(n31),.Q(n80));
  AO22X1 U247(.IN1(N321),.IN2(n32),.IN3(\sum[0][21] ),.IN4(n31),.Q(n81));
  AO22X1 U248(.IN1(N322),.IN2(n33),.IN3(\sum[0][22] ),.IN4(n31),.Q(n82));
  AO22X1 U249(.IN1(N323),.IN2(n32),.IN3(\sum[0][23] ),.IN4(n31),.Q(n83));
  AO22X1 U250(.IN1(n30),.IN2(N300),.IN3(\sum[1][0] ),.IN4(n44),.Q(n84));
  AO22X1 U251(.IN1(n29),.IN2(N301),.IN3(\sum[1][1] ),.IN4(n44),.Q(n85));
  AO22X1 U252(.IN1(n30),.IN2(N302),.IN3(\sum[1][2] ),.IN4(n44),.Q(n86));
  AO22X1 U253(.IN1(n29),.IN2(N303),.IN3(\sum[1][3] ),.IN4(n44),.Q(n87));
  AO22X1 U254(.IN1(n30),.IN2(N304),.IN3(\sum[1][4] ),.IN4(n44),.Q(n88));
  AO22X1 U255(.IN1(n29),.IN2(N305),.IN3(\sum[1][5] ),.IN4(n44),.Q(n89));
  AO22X1 U256(.IN1(n29),.IN2(N306),.IN3(\sum[1][6] ),.IN4(n44),.Q(n90));
  AO22X1 U257(.IN1(n29),.IN2(N307),.IN3(\sum[1][7] ),.IN4(n44),.Q(n91));
  AO22X1 U258(.IN1(n29),.IN2(N308),.IN3(\sum[1][8] ),.IN4(n44),.Q(n92));
  AO22X1 U259(.IN1(n29),.IN2(N309),.IN3(\sum[1][9] ),.IN4(n44),.Q(n93));
  AO22X1 U260(.IN1(n29),.IN2(N310),.IN3(\sum[1][10] ),.IN4(n44),.Q(n94));
  AO22X1 U261(.IN1(n29),.IN2(N311),.IN3(\sum[1][11] ),.IN4(n44),.Q(n95));
  AO22X1 U262(.IN1(n30),.IN2(N312),.IN3(\sum[1][12] ),.IN4(n28),.Q(n96));
  AO22X1 U263(.IN1(n30),.IN2(N313),.IN3(\sum[1][13] ),.IN4(n28),.Q(n97));
  AO22X1 U264(.IN1(n30),.IN2(N314),.IN3(\sum[1][14] ),.IN4(n28),.Q(n98));
  AO22X1 U265(.IN1(n30),.IN2(N315),.IN3(\sum[1][15] ),.IN4(n28),.Q(n99));
  AO22X1 U266(.IN1(n30),.IN2(N316),.IN3(\sum[1][16] ),.IN4(n28),.Q(n100));
  AO22X1 U267(.IN1(n30),.IN2(N317),.IN3(\sum[1][17] ),.IN4(n28),.Q(n101));
  AO22X1 U268(.IN1(n30),.IN2(N318),.IN3(\sum[1][18] ),.IN4(n28),.Q(n102));
  AO22X1 U269(.IN1(n29),.IN2(N319),.IN3(\sum[1][19] ),.IN4(n28),.Q(n103));
  AO22X1 U270(.IN1(n30),.IN2(N320),.IN3(\sum[1][20] ),.IN4(n28),.Q(n104));
  AO22X1 U271(.IN1(n29),.IN2(N321),.IN3(\sum[1][21] ),.IN4(n28),.Q(n105));
  AO22X1 U272(.IN1(n30),.IN2(N322),.IN3(\sum[1][22] ),.IN4(n28),.Q(n106));
  AO22X1 U273(.IN1(n29),.IN2(N323),.IN3(\sum[1][23] ),.IN4(n28),.Q(n107));
  NAND3X0 U274(.IN1(n375),.IN2(n41),.IN3(N26),.QN(n44));
  AO22X1 U275(.IN1(n24),.IN2(N300),.IN3(\sum[2][0] ),.IN4(n26),.Q(n108));
  AO22X1 U276(.IN1(n24),.IN2(N301),.IN3(\sum[2][1] ),.IN4(n26),.Q(n109));
  AO22X1 U277(.IN1(n24),.IN2(N302),.IN3(\sum[2][2] ),.IN4(n26),.Q(n110));
  AO22X1 U278(.IN1(n24),.IN2(N303),.IN3(\sum[2][3] ),.IN4(n26),.Q(n111));
  AO22X1 U279(.IN1(n24),.IN2(N304),.IN3(\sum[2][4] ),.IN4(n26),.Q(n112));
  AO22X1 U280(.IN1(n23),.IN2(N305),.IN3(\sum[2][5] ),.IN4(n26),.Q(n113));
  AO22X1 U281(.IN1(n23),.IN2(N306),.IN3(\sum[2][6] ),.IN4(n26),.Q(n114));
  AO22X1 U282(.IN1(n23),.IN2(N307),.IN3(\sum[2][7] ),.IN4(n26),.Q(n115));
  AO22X1 U283(.IN1(n23),.IN2(N308),.IN3(\sum[2][8] ),.IN4(n26),.Q(n116));
  AO22X1 U284(.IN1(n23),.IN2(N309),.IN3(\sum[2][9] ),.IN4(n26),.Q(n117));
  AO22X1 U285(.IN1(n23),.IN2(N310),.IN3(\sum[2][10] ),.IN4(n26),.Q(n118));
  AO22X1 U286(.IN1(n23),.IN2(N311),.IN3(\sum[2][11] ),.IN4(n26),.Q(n119));
  AO22X1 U287(.IN1(n22),.IN2(N312),.IN3(\sum[2][12] ),.IN4(n27),.Q(n120));
  AO22X1 U288(.IN1(n22),.IN2(N313),.IN3(\sum[2][13] ),.IN4(n27),.Q(n121));
  AO22X1 U289(.IN1(n22),.IN2(N314),.IN3(\sum[2][14] ),.IN4(n27),.Q(n122));
  AO22X1 U290(.IN1(n22),.IN2(N315),.IN3(\sum[2][15] ),.IN4(n27),.Q(n123));
  AO22X1 U291(.IN1(n22),.IN2(N316),.IN3(\sum[2][16] ),.IN4(n27),.Q(n124));
  AO22X1 U292(.IN1(n22),.IN2(N317),.IN3(\sum[2][17] ),.IN4(n27),.Q(n125));
  AO22X1 U293(.IN1(n22),.IN2(N318),.IN3(\sum[2][18] ),.IN4(n27),.Q(n126));
  AO22X1 U294(.IN1(n21),.IN2(N319),.IN3(\sum[2][19] ),.IN4(n27),.Q(n127));
  AO22X1 U295(.IN1(n21),.IN2(N320),.IN3(\sum[2][20] ),.IN4(n27),.Q(n128));
  AO22X1 U296(.IN1(n21),.IN2(N321),.IN3(\sum[2][21] ),.IN4(n27),.Q(n129));
  AO22X1 U297(.IN1(n21),.IN2(N322),.IN3(\sum[2][22] ),.IN4(n27),.Q(n130));
  AO22X1 U298(.IN1(n21),.IN2(N323),.IN3(\sum[2][23] ),.IN4(n27),.Q(n131));
  AO22X1 U299(.IN1(n20),.IN2(N300),.IN3(\sum[3][0] ),.IN4(n48),.Q(n132));
  AO22X1 U300(.IN1(n19),.IN2(N301),.IN3(\sum[3][1] ),.IN4(n48),.Q(n133));
  AO22X1 U301(.IN1(n20),.IN2(N302),.IN3(\sum[3][2] ),.IN4(n48),.Q(n134));
  AO22X1 U302(.IN1(n19),.IN2(N303),.IN3(\sum[3][3] ),.IN4(n48),.Q(n135));
  AO22X1 U303(.IN1(n20),.IN2(N304),.IN3(\sum[3][4] ),.IN4(n48),.Q(n136));
  AO22X1 U304(.IN1(n19),.IN2(N305),.IN3(\sum[3][5] ),.IN4(n48),.Q(n137));
  AO22X1 U305(.IN1(n19),.IN2(N306),.IN3(\sum[3][6] ),.IN4(n48),.Q(n138));
  AO22X1 U306(.IN1(n19),.IN2(N307),.IN3(\sum[3][7] ),.IN4(n48),.Q(n139));
  AO22X1 U307(.IN1(n19),.IN2(N308),.IN3(\sum[3][8] ),.IN4(n48),.Q(n140));
  AO22X1 U308(.IN1(n19),.IN2(N309),.IN3(\sum[3][9] ),.IN4(n48),.Q(n141));
  AO22X1 U309(.IN1(n19),.IN2(N310),.IN3(\sum[3][10] ),.IN4(n48),.Q(n142));
  AO22X1 U310(.IN1(n19),.IN2(N311),.IN3(\sum[3][11] ),.IN4(n48),.Q(n143));
  AO22X1 U311(.IN1(n20),.IN2(N312),.IN3(\sum[3][12] ),.IN4(n18),.Q(n144));
  AO22X1 U312(.IN1(n20),.IN2(N313),.IN3(\sum[3][13] ),.IN4(n18),.Q(n145));
  AO22X1 U313(.IN1(n20),.IN2(N314),.IN3(\sum[3][14] ),.IN4(n18),.Q(n146));
  AO22X1 U314(.IN1(n20),.IN2(N315),.IN3(\sum[3][15] ),.IN4(n18),.Q(n147));
  AO22X1 U315(.IN1(n20),.IN2(N316),.IN3(\sum[3][16] ),.IN4(n18),.Q(n148));
  AO22X1 U316(.IN1(n20),.IN2(N317),.IN3(\sum[3][17] ),.IN4(n18),.Q(n149));
  AO22X1 U317(.IN1(n20),.IN2(N318),.IN3(\sum[3][18] ),.IN4(n18),.Q(n150));
  AO22X1 U318(.IN1(n19),.IN2(N319),.IN3(\sum[3][19] ),.IN4(n18),.Q(n151));
  AO22X1 U319(.IN1(n20),.IN2(N320),.IN3(\sum[3][20] ),.IN4(n18),.Q(n152));
  AO22X1 U320(.IN1(n19),.IN2(N321),.IN3(\sum[3][21] ),.IN4(n18),.Q(n153));
  AO22X1 U321(.IN1(n20),.IN2(N322),.IN3(\sum[3][22] ),.IN4(n18),.Q(n154));
  AO22X1 U322(.IN1(n19),.IN2(N323),.IN3(\sum[3][23] ),.IN4(n18),.Q(n155));
  AO22X1 U323(.IN1(N57),.IN2(n359),.IN3(\prod2[0][0][12] ),.IN4(n2),.Q(n156));
  AO22X1 U324(.IN1(N58),.IN2(n363),.IN3(\prod2[0][0][13] ),.IN4(n3),.Q(n157));
  AO22X1 U325(.IN1(N59),.IN2(n363),.IN3(\prod2[0][0][14] ),.IN4(n2),.Q(n158));
  AO22X1 U326(.IN1(N60),.IN2(n363),.IN3(\prod2[0][0][15] ),.IN4(n3),.Q(n159));
  AO22X1 U327(.IN1(N61),.IN2(n363),.IN3(\prod2[0][0][16] ),.IN4(n2),.Q(n160));
  AO22X1 U328(.IN1(N62),.IN2(n363),.IN3(\prod2[0][0][17] ),.IN4(n3),.Q(n161));
  AO22X1 U329(.IN1(N63),.IN2(n363),.IN3(\prod2[0][0][18] ),.IN4(n2),.Q(n162));
  AO22X1 U330(.IN1(N64),.IN2(n363),.IN3(\prod2[0][0][19] ),.IN4(n3),.Q(n163));
  AO22X1 U331(.IN1(N65),.IN2(n362),.IN3(\prod2[0][0][20] ),.IN4(n2),.Q(n164));
  AO22X1 U332(.IN1(N66),.IN2(n362),.IN3(\prod2[0][0][21] ),.IN4(n3),.Q(n165));
  AO22X1 U333(.IN1(N67),.IN2(n362),.IN3(\prod2[0][0][22] ),.IN4(n2),.Q(n166));
  AO22X1 U334(.IN1(N68),.IN2(n362),.IN3(\prod2[0][0][23] ),.IN4(n3),.Q(n167));
  AO22X1 U335(.IN1(N75),.IN2(n362),.IN3(\prod2[0][1][6] ),.IN4(n2),.Q(n168));
  AO22X1 U336(.IN1(N76),.IN2(n362),.IN3(\prod2[0][1][7] ),.IN4(n3),.Q(n169));
  AO22X1 U337(.IN1(N77),.IN2(n362),.IN3(\prod2[0][1][8] ),.IN4(n2),.Q(n170));
  AO22X1 U338(.IN1(N78),.IN2(n361),.IN3(\prod2[0][1][9] ),.IN4(n3),.Q(n171));
  AO22X1 U339(.IN1(N79),.IN2(n361),.IN3(\prod2[0][1][10] ),.IN4(n2),.Q(n172));
  AO22X1 U340(.IN1(N80),.IN2(n361),.IN3(\prod2[0][1][11] ),.IN4(n3),.Q(n173));
  AO22X1 U341(.IN1(N81),.IN2(n361),.IN3(\prod2[0][1][12] ),.IN4(n2),.Q(n174));
  AO22X1 U342(.IN1(N82),.IN2(n361),.IN3(\prod2[0][1][13] ),.IN4(n3),.Q(n175));
  AO22X1 U343(.IN1(N83),.IN2(n361),.IN3(\prod2[0][1][14] ),.IN4(n2),.Q(n176));
  AO22X1 U344(.IN1(N84),.IN2(n361),.IN3(\prod2[0][1][15] ),.IN4(n3),.Q(n177));
  AO22X1 U345(.IN1(N85),.IN2(n360),.IN3(\prod2[0][1][16] ),.IN4(n2),.Q(n178));
  AO22X1 U346(.IN1(N86),.IN2(n360),.IN3(\prod2[0][1][17] ),.IN4(n3),.Q(n179));
  AO22X1 U347(.IN1(N93),.IN2(n360),.IN3(\prod2[0][2][6] ),.IN4(n2),.Q(n180));
  AO22X1 U348(.IN1(N94),.IN2(n360),.IN3(\prod2[0][2][7] ),.IN4(n3),.Q(n181));
  AO22X1 U349(.IN1(N95),.IN2(n360),.IN3(\prod2[0][2][8] ),.IN4(n2),.Q(n182));
  AO22X1 U350(.IN1(N96),.IN2(n360),.IN3(\prod2[0][2][9] ),.IN4(n3),.Q(n183));
  AO22X1 U351(.IN1(N97),.IN2(n360),.IN3(\prod2[0][2][10] ),.IN4(n2),.Q(n184));
  AO22X1 U352(.IN1(N98),.IN2(n359),.IN3(\prod2[0][2][11] ),.IN4(n3),.Q(n185));
  AO22X1 U353(.IN1(N99),.IN2(n359),.IN3(\prod2[0][2][12] ),.IN4(n2),.Q(n186));
  AO22X1 U354(.IN1(N100),.IN2(n359),.IN3(\prod2[0][2][13] ),.IN4(n3),.Q(n187));
  AO22X1 U355(.IN1(N101),.IN2(n359),.IN3(\prod2[0][2][14] ),.IN4(n364),.Q(n188));
  AO22X1 U356(.IN1(N102),.IN2(n359),.IN3(\prod2[0][2][15] ),.IN4(n364),.Q(n189));
  AO22X1 U357(.IN1(N103),.IN2(n359),.IN3(\prod2[0][2][16] ),.IN4(n364),.Q(n190));
  AO22X1 U358(.IN1(N104),.IN2(n359),.IN3(\prod2[0][2][17] ),.IN4(n364),.Q(n191));
  AO22X1 U359(.IN1(N117),.IN2(n358),.IN3(\prod2[0][3][0] ),.IN4(n364),.Q(n192));
  AO22X1 U360(.IN1(N118),.IN2(n358),.IN3(\prod2[0][3][1] ),.IN4(n364),.Q(n193));
  AO22X1 U361(.IN1(N119),.IN2(n358),.IN3(\prod2[0][3][2] ),.IN4(n364),.Q(n194));
  AO22X1 U362(.IN1(N120),.IN2(n358),.IN3(\prod2[0][3][3] ),.IN4(n364),.Q(n195));
  AO22X1 U363(.IN1(N121),.IN2(n358),.IN3(\prod2[0][3][4] ),.IN4(n364),.Q(n196));
  AO22X1 U364(.IN1(N122),.IN2(n358),.IN3(\prod2[0][3][5] ),.IN4(n364),.Q(n197));
  AO22X1 U365(.IN1(N123),.IN2(n358),.IN3(\prod2[0][3][6] ),.IN4(n364),.Q(n198));
  AO22X1 U366(.IN1(N124),.IN2(n357),.IN3(\prod2[0][3][7] ),.IN4(n364),.Q(n199));
  AO22X1 U367(.IN1(N125),.IN2(n357),.IN3(\prod2[0][3][8] ),.IN4(n364),.Q(n200));
  AO22X1 U368(.IN1(N126),.IN2(n357),.IN3(\prod2[0][3][9] ),.IN4(n364),.Q(n201));
  AO22X1 U369(.IN1(N127),.IN2(n357),.IN3(\prod2[0][3][10] ),.IN4(n364),.Q(n202));
  AO22X1 U370(.IN1(N128),.IN2(n357),.IN3(\prod2[0][3][11] ),.IN4(n364),.Q(n203));
  AO22X1 U371(.IN1(n17),.IN2(N57),.IN3(\prod2[1][0][12] ),.IN4(n14),.Q(n204));
  AO22X1 U372(.IN1(n16),.IN2(N58),.IN3(\prod2[1][0][13] ),.IN4(n14),.Q(n205));
  AO22X1 U373(.IN1(n16),.IN2(N59),.IN3(\prod2[1][0][14] ),.IN4(n14),.Q(n206));
  AO22X1 U374(.IN1(n15),.IN2(N60),.IN3(\prod2[1][0][15] ),.IN4(n14),.Q(n207));
  AO22X1 U375(.IN1(n17),.IN2(N61),.IN3(\prod2[1][0][16] ),.IN4(n14),.Q(n208));
  AO22X1 U376(.IN1(n17),.IN2(N62),.IN3(\prod2[1][0][17] ),.IN4(n14),.Q(n209));
  AO22X1 U377(.IN1(n16),.IN2(N63),.IN3(\prod2[1][0][18] ),.IN4(n14),.Q(n210));
  AO22X1 U378(.IN1(n15),.IN2(N64),.IN3(\prod2[1][0][19] ),.IN4(n14),.Q(n211));
  AO22X1 U379(.IN1(n17),.IN2(N65),.IN3(\prod2[1][0][20] ),.IN4(n14),.Q(n212));
  AO22X1 U380(.IN1(n15),.IN2(N66),.IN3(\prod2[1][0][21] ),.IN4(n14),.Q(n213));
  AO22X1 U381(.IN1(n15),.IN2(N67),.IN3(\prod2[1][0][22] ),.IN4(n14),.Q(n214));
  AO22X1 U382(.IN1(n15),.IN2(N68),.IN3(\prod2[1][0][23] ),.IN4(n14),.Q(n215));
  AO22X1 U383(.IN1(n15),.IN2(N75),.IN3(\prod2[1][1][6] ),.IN4(n13),.Q(n216));
  AO22X1 U384(.IN1(n15),.IN2(N76),.IN3(\prod2[1][1][7] ),.IN4(n13),.Q(n217));
  AO22X1 U385(.IN1(n15),.IN2(N77),.IN3(\prod2[1][1][8] ),.IN4(n13),.Q(n218));
  AO22X1 U386(.IN1(n15),.IN2(N78),.IN3(\prod2[1][1][9] ),.IN4(n13),.Q(n219));
  AO22X1 U387(.IN1(n16),.IN2(N79),.IN3(\prod2[1][1][10] ),.IN4(n13),.Q(n220));
  AO22X1 U388(.IN1(n16),.IN2(N80),.IN3(\prod2[1][1][11] ),.IN4(n13),.Q(n221));
  AO22X1 U389(.IN1(n16),.IN2(N81),.IN3(\prod2[1][1][12] ),.IN4(n13),.Q(n222));
  AO22X1 U390(.IN1(n16),.IN2(N82),.IN3(\prod2[1][1][13] ),.IN4(n13),.Q(n223));
  AO22X1 U391(.IN1(n16),.IN2(N83),.IN3(\prod2[1][1][14] ),.IN4(n13),.Q(n224));
  AO22X1 U392(.IN1(n16),.IN2(N84),.IN3(\prod2[1][1][15] ),.IN4(n13),.Q(n225));
  AO22X1 U393(.IN1(n16),.IN2(N85),.IN3(\prod2[1][1][16] ),.IN4(n13),.Q(n226));
  AO22X1 U394(.IN1(n17),.IN2(N86),.IN3(\prod2[1][1][17] ),.IN4(n13),.Q(n227));
  AO22X1 U395(.IN1(n16),.IN2(N93),.IN3(\prod2[1][2][6] ),.IN4(n12),.Q(n228));
  AO22X1 U396(.IN1(n15),.IN2(N94),.IN3(\prod2[1][2][7] ),.IN4(n12),.Q(n229));
  AO22X1 U397(.IN1(n17),.IN2(N95),.IN3(\prod2[1][2][8] ),.IN4(n12),.Q(n230));
  AO22X1 U398(.IN1(n16),.IN2(N96),.IN3(\prod2[1][2][9] ),.IN4(n12),.Q(n231));
  AO22X1 U399(.IN1(n15),.IN2(N97),.IN3(\prod2[1][2][10] ),.IN4(n12),.Q(n232));
  AO22X1 U400(.IN1(n17),.IN2(N98),.IN3(\prod2[1][2][11] ),.IN4(n12),.Q(n233));
  AO22X1 U401(.IN1(n17),.IN2(N99),.IN3(\prod2[1][2][12] ),.IN4(n12),.Q(n234));
  AO22X1 U402(.IN1(n15),.IN2(N100),.IN3(\prod2[1][2][13] ),.IN4(n12),.Q(n235));
  AO22X1 U403(.IN1(n16),.IN2(N101),.IN3(\prod2[1][2][14] ),.IN4(n12),.Q(n236));
  AO22X1 U404(.IN1(n15),.IN2(N102),.IN3(\prod2[1][2][15] ),.IN4(n12),.Q(n237));
  AO22X1 U405(.IN1(n15),.IN2(N103),.IN3(\prod2[1][2][16] ),.IN4(n12),.Q(n238));
  AO22X1 U406(.IN1(n17),.IN2(N104),.IN3(\prod2[1][2][17] ),.IN4(n12),.Q(n239));
  AO22X1 U407(.IN1(n17),.IN2(N117),.IN3(\prod2[1][3][0] ),.IN4(n11),.Q(n240));
  AO22X1 U408(.IN1(n17),.IN2(N118),.IN3(\prod2[1][3][1] ),.IN4(n11),.Q(n241));
  AO22X1 U409(.IN1(n17),.IN2(N119),.IN3(\prod2[1][3][2] ),.IN4(n11),.Q(n242));
  AO22X1 U410(.IN1(n17),.IN2(N120),.IN3(\prod2[1][3][3] ),.IN4(n11),.Q(n243));
  AO22X1 U411(.IN1(n17),.IN2(N121),.IN3(\prod2[1][3][4] ),.IN4(n11),.Q(n244));
  AO22X1 U412(.IN1(n17),.IN2(N122),.IN3(\prod2[1][3][5] ),.IN4(n11),.Q(n245));
  AO22X1 U413(.IN1(n17),.IN2(N123),.IN3(\prod2[1][3][6] ),.IN4(n11),.Q(n246));
  AO22X1 U414(.IN1(n17),.IN2(N124),.IN3(\prod2[1][3][7] ),.IN4(n11),.Q(n247));
  AO22X1 U415(.IN1(n16),.IN2(N125),.IN3(\prod2[1][3][8] ),.IN4(n11),.Q(n248));
  AO22X1 U416(.IN1(n16),.IN2(N126),.IN3(\prod2[1][3][9] ),.IN4(n11),.Q(n249));
  AO22X1 U417(.IN1(n15),.IN2(N127),.IN3(\prod2[1][3][10] ),.IN4(n11),.Q(n250));
  AO22X1 U418(.IN1(n16),.IN2(N128),.IN3(\prod2[1][3][11] ),.IN4(n11),.Q(n251));
  AO22X1 U419(.IN1(n9),.IN2(N57),.IN3(\prod2[2][0][12] ),.IN4(n51),.Q(n252));
  AO22X1 U420(.IN1(n10),.IN2(N58),.IN3(\prod2[2][0][13] ),.IN4(n51),.Q(n253));
  AO22X1 U421(.IN1(n8),.IN2(N59),.IN3(\prod2[2][0][14] ),.IN4(n51),.Q(n254));
  AO22X1 U422(.IN1(n7),.IN2(N60),.IN3(\prod2[2][0][15] ),.IN4(n51),.Q(n255));
  AO22X1 U423(.IN1(n10),.IN2(N61),.IN3(\prod2[2][0][16] ),.IN4(n51),.Q(n256));
  AO22X1 U424(.IN1(n9),.IN2(N62),.IN3(\prod2[2][0][17] ),.IN4(n51),.Q(n257));
  AO22X1 U425(.IN1(n8),.IN2(N63),.IN3(\prod2[2][0][18] ),.IN4(n51),.Q(n258));
  AO22X1 U426(.IN1(n7),.IN2(N64),.IN3(\prod2[2][0][19] ),.IN4(n51),.Q(n259));
  AO22X1 U427(.IN1(n9),.IN2(N65),.IN3(\prod2[2][0][20] ),.IN4(n51),.Q(n260));
  AO22X1 U428(.IN1(n7),.IN2(N66),.IN3(\prod2[2][0][21] ),.IN4(n51),.Q(n261));
  AO22X1 U429(.IN1(n7),.IN2(N67),.IN3(\prod2[2][0][22] ),.IN4(n51),.Q(n262));
  AO22X1 U430(.IN1(n7),.IN2(N68),.IN3(\prod2[2][0][23] ),.IN4(n51),.Q(n263));
  AO22X1 U431(.IN1(n7),.IN2(N75),.IN3(\prod2[2][1][6] ),.IN4(n6),.Q(n264));
  AO22X1 U432(.IN1(n7),.IN2(N76),.IN3(\prod2[2][1][7] ),.IN4(n6),.Q(n265));
  AO22X1 U433(.IN1(n7),.IN2(N77),.IN3(\prod2[2][1][8] ),.IN4(n6),.Q(n266));
  AO22X1 U434(.IN1(n7),.IN2(N78),.IN3(\prod2[2][1][9] ),.IN4(n6),.Q(n267));
  AO22X1 U435(.IN1(n8),.IN2(N79),.IN3(\prod2[2][1][10] ),.IN4(n6),.Q(n268));
  AO22X1 U436(.IN1(n8),.IN2(N80),.IN3(\prod2[2][1][11] ),.IN4(n6),.Q(n269));
  AO22X1 U437(.IN1(n8),.IN2(N81),.IN3(\prod2[2][1][12] ),.IN4(n6),.Q(n270));
  AO22X1 U438(.IN1(n8),.IN2(N82),.IN3(\prod2[2][1][13] ),.IN4(n6),.Q(n271));
  AO22X1 U439(.IN1(n8),.IN2(N83),.IN3(\prod2[2][1][14] ),.IN4(n6),.Q(n272));
  AO22X1 U440(.IN1(n8),.IN2(N84),.IN3(\prod2[2][1][15] ),.IN4(n6),.Q(n273));
  AO22X1 U441(.IN1(n8),.IN2(N85),.IN3(\prod2[2][1][16] ),.IN4(n6),.Q(n274));
  AO22X1 U442(.IN1(n9),.IN2(N86),.IN3(\prod2[2][1][17] ),.IN4(n6),.Q(n275));
  AO22X1 U443(.IN1(n9),.IN2(N93),.IN3(\prod2[2][2][6] ),.IN4(n5),.Q(n276));
  AO22X1 U444(.IN1(n9),.IN2(N94),.IN3(\prod2[2][2][7] ),.IN4(n5),.Q(n277));
  AO22X1 U445(.IN1(n9),.IN2(N95),.IN3(\prod2[2][2][8] ),.IN4(n5),.Q(n278));
  AO22X1 U446(.IN1(n9),.IN2(N96),.IN3(\prod2[2][2][9] ),.IN4(n5),.Q(n279));
  AO22X1 U447(.IN1(n9),.IN2(N97),.IN3(\prod2[2][2][10] ),.IN4(n5),.Q(n280));
  AO22X1 U448(.IN1(n9),.IN2(N98),.IN3(\prod2[2][2][11] ),.IN4(n5),.Q(n281));
  AO22X1 U449(.IN1(n10),.IN2(N99),.IN3(\prod2[2][2][12] ),.IN4(n5),.Q(n282));
  AO22X1 U450(.IN1(n9),.IN2(N100),.IN3(\prod2[2][2][13] ),.IN4(n5),.Q(n283));
  AO22X1 U451(.IN1(n8),.IN2(N101),.IN3(\prod2[2][2][14] ),.IN4(n5),.Q(n284));
  AO22X1 U452(.IN1(n7),.IN2(N102),.IN3(\prod2[2][2][15] ),.IN4(n5),.Q(n285));
  AO22X1 U453(.IN1(n7),.IN2(N103),.IN3(\prod2[2][2][16] ),.IN4(n5),.Q(n286));
  AO22X1 U454(.IN1(n10),.IN2(N104),.IN3(\prod2[2][2][17] ),.IN4(n5),.Q(n287));
  AO22X1 U455(.IN1(n10),.IN2(N117),.IN3(\prod2[2][3][0] ),.IN4(n4),.Q(n288));
  AO22X1 U456(.IN1(n10),.IN2(N118),.IN3(\prod2[2][3][1] ),.IN4(n4),.Q(n289));
  AO22X1 U457(.IN1(n10),.IN2(N119),.IN3(\prod2[2][3][2] ),.IN4(n4),.Q(n290));
  AO22X1 U458(.IN1(n10),.IN2(N120),.IN3(\prod2[2][3][3] ),.IN4(n4),.Q(n291));
  AO22X1 U459(.IN1(n10),.IN2(N121),.IN3(\prod2[2][3][4] ),.IN4(n4),.Q(n292));
  AO22X1 U460(.IN1(n10),.IN2(N122),.IN3(\prod2[2][3][5] ),.IN4(n4),.Q(n293));
  AO22X1 U461(.IN1(n10),.IN2(N123),.IN3(\prod2[2][3][6] ),.IN4(n4),.Q(n294));
  AO22X1 U462(.IN1(n10),.IN2(N124),.IN3(\prod2[2][3][7] ),.IN4(n4),.Q(n295));
  AO22X1 U463(.IN1(n9),.IN2(N125),.IN3(\prod2[2][3][8] ),.IN4(n4),.Q(n296));
  AO22X1 U464(.IN1(n8),.IN2(N126),.IN3(\prod2[2][3][9] ),.IN4(n4),.Q(n297));
  AO22X1 U465(.IN1(n7),.IN2(N127),.IN3(\prod2[2][3][10] ),.IN4(n4),.Q(n298));
  AO22X1 U466(.IN1(n8),.IN2(N128),.IN3(\prod2[2][3][11] ),.IN4(n4),.Q(n299));
  AO22X1 U467(.IN1(n34),.IN2(N57),.IN3(\prod2[3][0][12] ),.IN4(n356),.Q(n300));
  AO22X1 U468(.IN1(n353),.IN2(N58),.IN3(\prod2[3][0][13] ),.IN4(n355),.Q(n301));
  AO22X1 U469(.IN1(n353),.IN2(N59),.IN3(\prod2[3][0][14] ),.IN4(n354),.Q(n302));
  AO22X1 U470(.IN1(n353),.IN2(N60),.IN3(\prod2[3][0][15] ),.IN4(n356),.Q(n303));
  AO22X1 U471(.IN1(n353),.IN2(N61),.IN3(\prod2[3][0][16] ),.IN4(n355),.Q(n304));
  AO22X1 U472(.IN1(n353),.IN2(N62),.IN3(\prod2[3][0][17] ),.IN4(n354),.Q(n305));
  AO22X1 U473(.IN1(n353),.IN2(N63),.IN3(\prod2[3][0][18] ),.IN4(n356),.Q(n306));
  AO22X1 U474(.IN1(n40),.IN2(N64),.IN3(\prod2[3][0][19] ),.IN4(n355),.Q(n307));
  AO22X1 U475(.IN1(n40),.IN2(N65),.IN3(\prod2[3][0][20] ),.IN4(n354),.Q(n308));
  AO22X1 U476(.IN1(n40),.IN2(N66),.IN3(\prod2[3][0][21] ),.IN4(n356),.Q(n309));
  AO22X1 U477(.IN1(n40),.IN2(N67),.IN3(\prod2[3][0][22] ),.IN4(n355),.Q(n310));
  AO22X1 U478(.IN1(n40),.IN2(N68),.IN3(\prod2[3][0][23] ),.IN4(n354),.Q(n311));
  AO22X1 U479(.IN1(n40),.IN2(N75),.IN3(\prod2[3][1][6] ),.IN4(n354),.Q(n312));
  AO22X1 U480(.IN1(n40),.IN2(N76),.IN3(\prod2[3][1][7] ),.IN4(n354),.Q(n313));
  AO22X1 U481(.IN1(n40),.IN2(N77),.IN3(\prod2[3][1][8] ),.IN4(n354),.Q(n314));
  AO22X1 U482(.IN1(n39),.IN2(N78),.IN3(\prod2[3][1][9] ),.IN4(n354),.Q(n315));
  AO22X1 U483(.IN1(n39),.IN2(N79),.IN3(\prod2[3][1][10] ),.IN4(n354),.Q(n316));
  AO22X1 U484(.IN1(n39),.IN2(N80),.IN3(\prod2[3][1][11] ),.IN4(n354),.Q(n317));
  AO22X1 U485(.IN1(n39),.IN2(N81),.IN3(\prod2[3][1][12] ),.IN4(n354),.Q(n318));
  AO22X1 U486(.IN1(n39),.IN2(N82),.IN3(\prod2[3][1][13] ),.IN4(n354),.Q(n319));
  AO22X1 U487(.IN1(n39),.IN2(N83),.IN3(\prod2[3][1][14] ),.IN4(n354),.Q(n320));
  AO22X1 U488(.IN1(n39),.IN2(N84),.IN3(\prod2[3][1][15] ),.IN4(n354),.Q(n321));
  AO22X1 U489(.IN1(n39),.IN2(N85),.IN3(\prod2[3][1][16] ),.IN4(n354),.Q(n322));
  AO22X1 U490(.IN1(n37),.IN2(N86),.IN3(\prod2[3][1][17] ),.IN4(n354),.Q(n323));
  AO22X1 U491(.IN1(n37),.IN2(N93),.IN3(\prod2[3][2][6] ),.IN4(n355),.Q(n324));
  AO22X1 U492(.IN1(n37),.IN2(N94),.IN3(\prod2[3][2][7] ),.IN4(n355),.Q(n325));
  AO22X1 U493(.IN1(n37),.IN2(N95),.IN3(\prod2[3][2][8] ),.IN4(n355),.Q(n326));
  AO22X1 U494(.IN1(n37),.IN2(N96),.IN3(\prod2[3][2][9] ),.IN4(n355),.Q(n327));
  AO22X1 U495(.IN1(n37),.IN2(N97),.IN3(\prod2[3][2][10] ),.IN4(n355),.Q(n328));
  AO22X1 U496(.IN1(n37),.IN2(N98),.IN3(\prod2[3][2][11] ),.IN4(n355),.Q(n329));
  AO22X1 U497(.IN1(n36),.IN2(N99),.IN3(\prod2[3][2][12] ),.IN4(n355),.Q(n330));
  AO22X1 U498(.IN1(n36),.IN2(N100),.IN3(\prod2[3][2][13] ),.IN4(n355),.Q(n331));
  AO22X1 U499(.IN1(n36),.IN2(N101),.IN3(\prod2[3][2][14] ),.IN4(n355),.Q(n332));
  AO22X1 U500(.IN1(n36),.IN2(N102),.IN3(\prod2[3][2][15] ),.IN4(n355),.Q(n333));
  AO22X1 U501(.IN1(n36),.IN2(N103),.IN3(\prod2[3][2][16] ),.IN4(n355),.Q(n334));
  AO22X1 U502(.IN1(n36),.IN2(N104),.IN3(\prod2[3][2][17] ),.IN4(n355),.Q(n335));
  AO22X1 U503(.IN1(n36),.IN2(N117),.IN3(\prod2[3][3][0] ),.IN4(n356),.Q(n336));
  AO22X1 U504(.IN1(n36),.IN2(N118),.IN3(\prod2[3][3][1] ),.IN4(n356),.Q(n337));
  AO22X1 U505(.IN1(n35),.IN2(N119),.IN3(\prod2[3][3][2] ),.IN4(n356),.Q(n338));
  AO22X1 U506(.IN1(n35),.IN2(N120),.IN3(\prod2[3][3][3] ),.IN4(n356),.Q(n339));
  AO22X1 U507(.IN1(n37),.IN2(N121),.IN3(\prod2[3][3][4] ),.IN4(n356),.Q(n340));
  AO22X1 U508(.IN1(n35),.IN2(N122),.IN3(\prod2[3][3][5] ),.IN4(n356),.Q(n341));
  AO22X1 U509(.IN1(n35),.IN2(N123),.IN3(\prod2[3][3][6] ),.IN4(n356),.Q(n342));
  AO22X1 U510(.IN1(n35),.IN2(N124),.IN3(\prod2[3][3][7] ),.IN4(n356),.Q(n343));
  AO22X1 U511(.IN1(n35),.IN2(N125),.IN3(\prod2[3][3][8] ),.IN4(n356),.Q(n344));
  AO22X1 U512(.IN1(n35),.IN2(N126),.IN3(\prod2[3][3][9] ),.IN4(n356),.Q(n345));
  AO22X1 U513(.IN1(n35),.IN2(N127),.IN3(\prod2[3][3][10] ),.IN4(n356),.Q(n346));
  AO22X1 U514(.IN1(n34),.IN2(N128),.IN3(\prod2[3][3][11] ),.IN4(n356),.Q(n347));
  AO22X1 U515(.IN1(N26),.IN2(n372),.IN3(n52),.IN4(n53),.Q(n348));
  AND2X1 U516(.IN1(n373),.IN2(n43),.Q(n52));
  AO22X1 U517(.IN1(n377),.IN2(n25),.IN3(ready_o),.IN4(n373),.Q(n349));
  AO21X1 U518(.IN1(s_state),.IN2(n55),.IN3(s_start_i),.Q(n350));
  OAI21X1 U519(.IN1(n56),.IN2(n38),.IN3(n57),.QN(n351));
  NAND3X0 U520(.IN1(n34),.IN2(n373),.IN3(n53),.QN(n57));
  AO22X1 U521(.IN1(n58),.IN2(N25),.IN3(n59),.IN4(n53),.Q(n352));
  NAND3X0 U522(.IN1(s_state),.IN2(n49),.IN3(\count[2] ),.QN(n55));
  NAND3X0 U523(.IN1(n41),.IN2(n38),.IN3(N26),.QN(n51));
  mul_24_DW01_add_3_inj add_0_root_add_0_root_add_208_3(.A({N273,N272,N271,N270,N269,N268,N267,N266,N265,N264,N263,N262,N261,N260,N259,N258,N257,N256,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.B({1'b0,1'b0,1'b0,1'b0,1'b0,N218,N217,N216,N215,N214,N213,N212,N211,N210,N209,N208,N207,N206,N205,N204,N203,N202,N201,N200}),.CI(1'b0),.SUM({N323,N322,N321,N320,N319,N318,N317,N316,N315,N314,N313,N312,N311,N310,N309,N308,N307,N306,N305,N304,N303,N302,N301,N300}));
  mul_24_DW_mult_uns_3_inj mult_194(.a({N69,N70,N71,N72,N73,N74}),.b({N87,N88,N89,N90,N91,N92}),.product({N68,N67,N66,N65,N64,N63,N62,N61,N60,N59,N58,N57}));
  mul_24_DW_mult_uns_2_inj mult_195(.a({N69,N70,N71,N72,N73,N74}),.b({N111,N112,N113,N114,N115,N116}),.product({N86,N85,N84,N83,N82,N81,N80,N79,N78,N77,N76,N75}));
  mul_24_DW_mult_uns_1_inj mult_196(.a({N105,N106,N107,N108,N109,N110}),.b({N87,N88,N89,N90,N91,N92}),.product({N104,N103,N102,N101,N100,N99,N98,N97,N96,N95,N94,N93}));
  mul_24_DW_mult_uns_0_inj mult_197(.a({N105,N106,N107,N108,N109,N110}),.b({N111,N112,N113,N114,N115,N116}),.product({N128,N127,N126,N125,N124,N123,N122,N121,N120,N119,N118,N117}));
  mul_24_DW01_add_2_inj add_2_root_add_0_root_add_223_3(.A({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\sum[3][23] ,\sum[3][22] ,\sum[3][21] ,\sum[3][20] ,\sum[3][19] ,\sum[3][18] ,\sum[3][17] ,\sum[3][16] ,\sum[3][15] ,\sum[3][14] ,\sum[3][13] ,\sum[3][12] ,\sum[3][11] ,\sum[3][10] ,\sum[3][9] ,\sum[3][8] ,\sum[3][7] ,\sum[3][6] ,\sum[3][5] ,\sum[3][4] ,\sum[3][3] ,\sum[3][2] ,\sum[3][1] ,\sum[3][0] }),.B({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\sum[2][23] ,\sum[2][22] ,\sum[2][21] ,\sum[2][20] ,\sum[2][19] ,\sum[2][18] ,\sum[2][17] ,\sum[2][16] ,\sum[2][15] ,\sum[2][14] ,\sum[2][13] ,\sum[2][12] ,\sum[2][11] ,\sum[2][10] ,\sum[2][9] ,\sum[2][8] ,\sum[2][7] ,\sum[2][6] ,\sum[2][5] ,\sum[2][4] ,\sum[2][3] ,\sum[2][2] ,\sum[2][1] ,\sum[2][0] ,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.CI(1'b0),.SUM({SYNOPSYS_UNCONNECTED__0,SYNOPSYS_UNCONNECTED__1,SYNOPSYS_UNCONNECTED__2,SYNOPSYS_UNCONNECTED__3,SYNOPSYS_UNCONNECTED__4,SYNOPSYS_UNCONNECTED__5,SYNOPSYS_UNCONNECTED__6,SYNOPSYS_UNCONNECTED__7,SYNOPSYS_UNCONNECTED__8,SYNOPSYS_UNCONNECTED__9,SYNOPSYS_UNCONNECTED__10,N412,N411,N410,N409,N408,N407,N406,N405,N404,N403,N402,N401,N400,N399,N398,N397,N396,N395,N394,N393,N392,N391,N390,N389,N388,N387,N386,N385,N384,N383,N382,N381,N380,N379,N378,N377,N376}));
  mul_24_DW01_add_1_inj add_1_root_add_0_root_add_223_3(.A({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,\sum[1][23] ,\sum[1][22] ,\sum[1][21] ,\sum[1][20] ,\sum[1][19] ,\sum[1][18] ,\sum[1][17] ,\sum[1][16] ,\sum[1][15] ,\sum[1][14] ,\sum[1][13] ,\sum[1][12] ,\sum[1][11] ,\sum[1][10] ,\sum[1][9] ,\sum[1][8] ,\sum[1][7] ,\sum[1][6] ,\sum[1][5] ,\sum[1][4] ,\sum[1][3] ,\sum[1][2] ,\sum[1][1] ,\sum[1][0] ,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.B({\sum[0][23] ,\sum[0][22] ,\sum[0][21] ,\sum[0][20] ,\sum[0][19] ,\sum[0][18] ,\sum[0][17] ,\sum[0][16] ,\sum[0][15] ,\sum[0][14] ,\sum[0][13] ,\sum[0][12] ,\sum[0][11] ,\sum[0][10] ,\sum[0][9] ,\sum[0][8] ,\sum[0][7] ,\sum[0][6] ,\sum[0][5] ,\sum[0][4] ,\sum[0][3] ,\sum[0][2] ,\sum[0][1] ,\sum[0][0] ,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.CI(1'b0),.SUM({N375,N374,N373,N372,N371,N370,N369,N368,N367,N366,N365,N364,N363,N362,N361,N360,N359,N358,N357,N356,N355,N354,N353,N352,N351,N350,N349,N348,N347,N346,N345,N344,N343,N342,N341,N340,SYNOPSYS_UNCONNECTED__11,SYNOPSYS_UNCONNECTED__12,SYNOPSYS_UNCONNECTED__13,SYNOPSYS_UNCONNECTED__14,SYNOPSYS_UNCONNECTED__15,SYNOPSYS_UNCONNECTED__16,SYNOPSYS_UNCONNECTED__17,SYNOPSYS_UNCONNECTED__18,SYNOPSYS_UNCONNECTED__19,SYNOPSYS_UNCONNECTED__20,SYNOPSYS_UNCONNECTED__21,SYNOPSYS_UNCONNECTED__22}));
  mul_24_DW01_add_0_inj add_0_root_add_0_root_add_223_3(.A({N375,N374,N373,N372,N371,N370,N369,N368,N367,N366,N365,N364,N363,N362,N361,N360,N359,N358,N357,N356,N355,N354,N353,N352,N351,N350,N349,N348,N347,N346,N345,N344,N343,N342,N341,N340,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.B({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,N412,N411,N410,N409,N408,N407,N406,N405,N404,N403,N402,N401,N400,N399,N398,N397,N396,N395,N394,N393,N392,N391,N390,N389,N388,N387,N386,N385,N384,N383,N382,N381,N380,N379,N378,N377,N376}),.CI(1'b0),.SUM(fract_o));
  FADDX1 desc714(.A(N162),.B(N236),.CI(\add_2_root_add_0_root_add_208_3/carry[13] ),.CO(\add_2_root_add_0_root_add_208_3/carry[14] ),.S(N263));
  FADDX1 desc715(.A(N161),.B(N235),.CI(\add_2_root_add_0_root_add_208_3/carry[14] ),.CO(\add_2_root_add_0_root_add_208_3/carry[15] ),.S(N264));
  FADDX1 desc716(.A(N160),.B(N234),.CI(\add_2_root_add_0_root_add_208_3/carry[15] ),.CO(\add_2_root_add_0_root_add_208_3/carry[16] ),.S(N265));
  FADDX1 desc717(.A(N159),.B(N233),.CI(\add_2_root_add_0_root_add_208_3/carry[16] ),.CO(\add_2_root_add_0_root_add_208_3/carry[17] ),.S(N266));
  FADDX1 desc718(.A(N158),.B(N232),.CI(\add_2_root_add_0_root_add_208_3/carry[17] ),.CO(\add_2_root_add_0_root_add_208_3/carry[18] ),.S(N267));
  FADDX1 desc719(.A(N192),.B(N292),.CI(\add_1_root_add_0_root_add_208_3/carry[7] ),.CO(\add_1_root_add_0_root_add_208_3/carry[8] ),.S(N207));
  FADDX1 desc720(.A(N191),.B(N291),.CI(\add_1_root_add_0_root_add_208_3/carry[8] ),.CO(\add_1_root_add_0_root_add_208_3/carry[9] ),.S(N208));
  FADDX1 desc721(.A(N190),.B(N290),.CI(\add_1_root_add_0_root_add_208_3/carry[9] ),.CO(\add_1_root_add_0_root_add_208_3/carry[10] ),.S(N209));
  FADDX1 desc722(.A(N189),.B(N289),.CI(\add_1_root_add_0_root_add_208_3/carry[10] ),.CO(\add_1_root_add_0_root_add_208_3/carry[11] ),.S(N210));
  FADDX1 desc723(.A(N188),.B(N288),.CI(\add_1_root_add_0_root_add_208_3/carry[11] ),.CO(\add_1_root_add_0_root_add_208_3/carry[12] ),.S(N211));
  NBUFFX2 U3(.INP(n364),.Z(n2));
  NBUFFX2 U4(.INP(n364),.Z(n3));
  NBUFFX2 U5(.INP(N34),.Z(n367));
  NBUFFX2 U6(.INP(N34),.Z(n366));
  NBUFFX2 U7(.INP(N34),.Z(n365));
  NBUFFX2 U8(.INP(N34),.Z(n368));
  NBUFFX2 U9(.INP(n45),.Z(n21));
  NBUFFX2 U10(.INP(n45),.Z(n23));
  NBUFFX2 U11(.INP(n45),.Z(n22));
  NBUFFX2 U12(.INP(n45),.Z(n24));
  INVX0 U13(.INP(n42),.ZN(n32));
  INVX0 U14(.INP(n42),.ZN(n33));
  INVX0 U15(.INP(n48),.ZN(n19));
  INVX0 U16(.INP(n48),.ZN(n20));
  INVX0 U17(.INP(n49),.ZN(n376));
  NAND2X1 U18(.IN1(n376),.IN2(n46),.QN(N34));
  INVX0 U19(.INP(n44),.ZN(n29));
  INVX0 U20(.INP(n44),.ZN(n30));
  NAND2X1 U21(.IN1(n375),.IN2(n43),.QN(n42));
  NAND2X1 U22(.IN1(n375),.IN2(n49),.QN(n48));
  NBUFFX2 U23(.INP(N132),.Z(n357));
  INVX0 U24(.INP(n47),.ZN(n375));
  NOR2X0 U25(.IN1(n46),.IN2(n47),.QN(n45));
  NBUFFX2 U26(.INP(N144),.Z(n40));
  NBUFFX2 U27(.INP(N144),.Z(n39));
  NBUFFX2 U28(.INP(N144),.Z(n36));
  NBUFFX2 U29(.INP(N144),.Z(n37));
  NBUFFX2 U30(.INP(N144),.Z(n35));
  NBUFFX2 U31(.INP(N144),.Z(n34));
  NBUFFX2 U32(.INP(N132),.Z(n363));
  NBUFFX2 U33(.INP(N132),.Z(n362));
  NBUFFX2 U34(.INP(N132),.Z(n361));
  NBUFFX2 U35(.INP(N132),.Z(n360));
  NBUFFX2 U36(.INP(N132),.Z(n359));
  NBUFFX2 U37(.INP(N132),.Z(n358));
  NBUFFX2 U38(.INP(N144),.Z(n353));
  INVX0 U39(.INP(n55),.ZN(n377));
  OA21X1 U40(.IN1(n374),.IN2(N25),.IN3(n373),.Q(n54));
  NOR2X0 U41(.IN1(N25),.IN2(n58),.QN(n59));
  INVX0 U42(.INP(n53),.ZN(n374));
  INVX0 U43(.INP(n50),.ZN(n15));
  INVX0 U44(.INP(n50),.ZN(n16));
  INVX0 U45(.INP(n50),.ZN(n17));
  INVX0 U46(.INP(n51),.ZN(n7));
  INVX0 U47(.INP(n51),.ZN(n8));
  INVX0 U48(.INP(n51),.ZN(n9));
  INVX0 U49(.INP(n51),.ZN(n10));
  INVX0 U50(.INP(n58),.ZN(n373));
  NOR2X0 U51(.IN1(N25),.IN2(N26),.QN(n49));
  NAND2X1 U52(.IN1(N26),.IN2(N25),.QN(n46));
  NBUFFX2 U53(.INP(N26),.Z(n1));
  NOR2X0 U54(.IN1(n376),.IN2(\count[2] ),.QN(N132));
  NAND2X1 U55(.IN1(s_state),.IN2(n364),.QN(n47));
  NOR2X0 U56(.IN1(n46),.IN2(\count[2] ),.QN(N144));
  NOR2X0 U57(.IN1(n377),.IN2(s_start_i),.QN(n53));
  INVX0 U58(.INP(n54),.ZN(n372));
  OA21X1 U59(.IN1(N26),.IN2(n374),.IN3(n54),.Q(n56));
  NAND2X1 U60(.IN1(n43),.IN2(n38),.QN(n50));
  NOR2X0 U61(.IN1(n41),.IN2(N26),.QN(n43));
  NOR2X0 U62(.IN1(s_state),.IN2(s_start_i),.QN(n58));
  MUX21X1 U63(.IN1(s_fracta_i[12:12]),.IN2(s_fracta_i[0:0]),.S(n1),.Q(N110));
  MUX21X1 U64(.IN1(s_fracta_i[13:13]),.IN2(s_fracta_i[1:1]),.S(n1),.Q(N109));
  MUX21X1 U65(.IN1(s_fracta_i[14:14]),.IN2(s_fracta_i[2:2]),.S(n1),.Q(N108));
  MUX21X1 U66(.IN1(s_fracta_i[15:15]),.IN2(s_fracta_i[3:3]),.S(n1),.Q(N107));
  MUX21X1 U67(.IN1(s_fracta_i[16:16]),.IN2(s_fracta_i[4:4]),.S(n1),.Q(N106));
  MUX21X1 U68(.IN1(s_fracta_i[17:17]),.IN2(s_fracta_i[5:5]),.S(n1),.Q(N105));
  MUX21X1 U69(.IN1(s_fractb_i[12:12]),.IN2(s_fractb_i[0:0]),.S(N25),.Q(N116));
  MUX21X1 U70(.IN1(s_fractb_i[13:13]),.IN2(s_fractb_i[1:1]),.S(N25),.Q(N115));
  MUX21X1 U71(.IN1(s_fractb_i[14:14]),.IN2(s_fractb_i[2:2]),.S(N25),.Q(N114));
  MUX21X1 U72(.IN1(s_fractb_i[15:15]),.IN2(s_fractb_i[3:3]),.S(N25),.Q(N113));
  MUX21X1 U73(.IN1(s_fractb_i[16:16]),.IN2(s_fractb_i[4:4]),.S(N25),.Q(N112));
  MUX21X1 U74(.IN1(s_fractb_i[17:17]),.IN2(s_fractb_i[5:5]),.S(N25),.Q(N111));
  MUX21X1 U75(.IN1(s_fractb_i[18:18]),.IN2(s_fractb_i[6:6]),.S(N25),.Q(N92));
  MUX21X1 U76(.IN1(s_fractb_i[19:19]),.IN2(s_fractb_i[7:7]),.S(N25),.Q(N91));
  MUX21X1 U77(.IN1(s_fractb_i[20:20]),.IN2(s_fractb_i[8:8]),.S(N25),.Q(N90));
  MUX21X1 U78(.IN1(s_fractb_i[21:21]),.IN2(s_fractb_i[9:9]),.S(N25),.Q(N89));
  MUX21X1 U79(.IN1(s_fractb_i[22:22]),.IN2(s_fractb_i[10:10]),.S(N25),.Q(N88));
  MUX21X1 U80(.IN1(s_fractb_i[23:23]),.IN2(s_fractb_i[11:11]),.S(N25),.Q(N87));
  MUX21X1 U81(.IN1(s_fracta_i[18:18]),.IN2(s_fracta_i[6:6]),.S(n1),.Q(N74));
  MUX21X1 U82(.IN1(s_fracta_i[19:19]),.IN2(s_fracta_i[7:7]),.S(n1),.Q(N73));
  MUX21X1 U83(.IN1(s_fracta_i[20:20]),.IN2(s_fracta_i[8:8]),.S(n1),.Q(N72));
  MUX21X1 U84(.IN1(s_fracta_i[21:21]),.IN2(s_fracta_i[9:9]),.S(n1),.Q(N71));
  MUX21X1 U85(.IN1(s_fracta_i[22:22]),.IN2(s_fracta_i[10:10]),.S(n1),.Q(N70));
  MUX21X1 U86(.IN1(s_fracta_i[23:23]),.IN2(s_fracta_i[11:11]),.S(n1),.Q(N69));
  INVX0 U87(.INP(n10),.ZN(n4));
  INVX0 U88(.INP(n9),.ZN(n5));
  INVX0 U89(.INP(n7),.ZN(n6));
  INVX0 U90(.INP(n15),.ZN(n11));
  INVX0 U91(.INP(n16),.ZN(n12));
  INVX0 U92(.INP(n17),.ZN(n13));
  INVX0 U93(.INP(n15),.ZN(n14));
  INVX0 U94(.INP(n20),.ZN(n18));
  INVX0 U95(.INP(n21),.ZN(n26));
  INVX0 U96(.INP(n21),.ZN(n27));
  INVX0 U97(.INP(n30),.ZN(n28));
  INVX0 U98(.INP(n33),.ZN(n31));
  INVX0 U99(.INP(n34),.ZN(n354));
  INVX0 U100(.INP(n34),.ZN(n355));
  INVX0 U101(.INP(n34),.ZN(n356));
  INVX0 U102(.INP(n357),.ZN(n364));
  INVX0 U103(.INP(N25),.ZN(n369));
  INVX0 U104(.INP(N25),.ZN(n370));
  INVX0 U105(.INP(N25),.ZN(n371));
  AND2X1 U106(.IN1(\add_1_root_add_0_root_add_208_3/carry[17] ),.IN2(N182),.Q(N218));
  XOR2X1 U107(.IN1(N182),.IN2(\add_1_root_add_0_root_add_208_3/carry[17] ),.Q(N217));
  AND2X1 U108(.IN1(\add_1_root_add_0_root_add_208_3/carry[16] ),.IN2(N183),.Q(\add_1_root_add_0_root_add_208_3/carry[17] ));
  XOR2X1 U109(.IN1(N183),.IN2(\add_1_root_add_0_root_add_208_3/carry[16] ),.Q(N216));
  AND2X1 U110(.IN1(\add_1_root_add_0_root_add_208_3/carry[15] ),.IN2(N184),.Q(\add_1_root_add_0_root_add_208_3/carry[16] ));
  XOR2X1 U111(.IN1(N184),.IN2(\add_1_root_add_0_root_add_208_3/carry[15] ),.Q(N215));
  AND2X1 U112(.IN1(\add_1_root_add_0_root_add_208_3/carry[14] ),.IN2(N185),.Q(\add_1_root_add_0_root_add_208_3/carry[15] ));
  XOR2X1 U113(.IN1(N185),.IN2(\add_1_root_add_0_root_add_208_3/carry[14] ),.Q(N214));
  AND2X1 U114(.IN1(\add_1_root_add_0_root_add_208_3/carry[13] ),.IN2(N186),.Q(\add_1_root_add_0_root_add_208_3/carry[14] ));
  XOR2X1 U115(.IN1(N186),.IN2(\add_1_root_add_0_root_add_208_3/carry[13] ),.Q(N213));
  AND2X1 U116(.IN1(\add_1_root_add_0_root_add_208_3/carry[12] ),.IN2(N187),.Q(\add_1_root_add_0_root_add_208_3/carry[13] ));
  XOR2X1 U117(.IN1(N187),.IN2(\add_1_root_add_0_root_add_208_3/carry[12] ),.Q(N212));
  AND2X1 U118(.IN1(N293),.IN2(N193),.Q(\add_1_root_add_0_root_add_208_3/carry[7] ));
  XOR2X1 U119(.IN1(N193),.IN2(N293),.Q(N206));
  XOR2X1 U120(.IN1(N152),.IN2(\add_2_root_add_0_root_add_208_3/carry[23] ),.Q(N273));
  AND2X1 U121(.IN1(\add_2_root_add_0_root_add_208_3/carry[22] ),.IN2(N153),.Q(\add_2_root_add_0_root_add_208_3/carry[23] ));
  XOR2X1 U122(.IN1(N153),.IN2(\add_2_root_add_0_root_add_208_3/carry[22] ),.Q(N272));
  AND2X1 U123(.IN1(\add_2_root_add_0_root_add_208_3/carry[21] ),.IN2(N154),.Q(\add_2_root_add_0_root_add_208_3/carry[22] ));
  XOR2X1 U124(.IN1(N154),.IN2(\add_2_root_add_0_root_add_208_3/carry[21] ),.Q(N271));
  AND2X1 U125(.IN1(\add_2_root_add_0_root_add_208_3/carry[20] ),.IN2(N155),.Q(\add_2_root_add_0_root_add_208_3/carry[21] ));
  XOR2X1 U126(.IN1(N155),.IN2(\add_2_root_add_0_root_add_208_3/carry[20] ),.Q(N270));
  AND2X1 U127(.IN1(\add_2_root_add_0_root_add_208_3/carry[19] ),.IN2(N156),.Q(\add_2_root_add_0_root_add_208_3/carry[20] ));
  XOR2X1 U128(.IN1(N156),.IN2(\add_2_root_add_0_root_add_208_3/carry[19] ),.Q(N269));
  AND2X1 U129(.IN1(\add_2_root_add_0_root_add_208_3/carry[18] ),.IN2(N157),.Q(\add_2_root_add_0_root_add_208_3/carry[19] ));
  XOR2X1 U130(.IN1(N157),.IN2(\add_2_root_add_0_root_add_208_3/carry[18] ),.Q(N268));
  AND2X1 U131(.IN1(N237),.IN2(N163),.Q(\add_2_root_add_0_root_add_208_3/carry[13] ));
  XOR2X1 U132(.IN1(N163),.IN2(N237),.Q(N262));
  MUX41X1 U133(.IN1(\prod2[0][0][12] ),.IN3(\prod2[2][0][12] ),.IN2(\prod2[1][0][12] ),.IN4(\prod2[3][0][12] ),.S0(n368),.S1(n41),.Q(N163));
  MUX41X1 U134(.IN1(\prod2[0][0][13] ),.IN3(\prod2[2][0][13] ),.IN2(\prod2[1][0][13] ),.IN4(\prod2[3][0][13] ),.S0(n368),.S1(n41),.Q(N162));
  MUX41X1 U135(.IN1(\prod2[0][0][14] ),.IN3(\prod2[2][0][14] ),.IN2(\prod2[1][0][14] ),.IN4(\prod2[3][0][14] ),.S0(n368),.S1(n41),.Q(N161));
  MUX41X1 U136(.IN1(\prod2[0][0][15] ),.IN3(\prod2[2][0][15] ),.IN2(\prod2[1][0][15] ),.IN4(\prod2[3][0][15] ),.S0(n368),.S1(n41),.Q(N160));
  MUX41X1 U137(.IN1(\prod2[0][0][16] ),.IN3(\prod2[2][0][16] ),.IN2(\prod2[1][0][16] ),.IN4(\prod2[3][0][16] ),.S0(n368),.S1(n41),.Q(N159));
  MUX41X1 U138(.IN1(\prod2[0][0][17] ),.IN3(\prod2[2][0][17] ),.IN2(\prod2[1][0][17] ),.IN4(\prod2[3][0][17] ),.S0(n368),.S1(n41),.Q(N158));
  MUX41X1 U139(.IN1(\prod2[0][0][18] ),.IN3(\prod2[2][0][18] ),.IN2(\prod2[1][0][18] ),.IN4(\prod2[3][0][18] ),.S0(n368),.S1(n41),.Q(N157));
  MUX41X1 U140(.IN1(\prod2[0][0][19] ),.IN3(\prod2[2][0][19] ),.IN2(\prod2[1][0][19] ),.IN4(\prod2[3][0][19] ),.S0(n368),.S1(n41),.Q(N156));
  MUX41X1 U141(.IN1(\prod2[0][0][20] ),.IN3(\prod2[2][0][20] ),.IN2(\prod2[1][0][20] ),.IN4(\prod2[3][0][20] ),.S0(n368),.S1(n41),.Q(N155));
  MUX41X1 U142(.IN1(\prod2[0][0][21] ),.IN3(\prod2[2][0][21] ),.IN2(\prod2[1][0][21] ),.IN4(\prod2[3][0][21] ),.S0(n368),.S1(n41),.Q(N154));
  MUX41X1 U143(.IN1(\prod2[0][0][22] ),.IN3(\prod2[2][0][22] ),.IN2(\prod2[1][0][22] ),.IN4(\prod2[3][0][22] ),.S0(n368),.S1(n41),.Q(N153));
  MUX41X1 U144(.IN1(\prod2[0][0][23] ),.IN3(\prod2[2][0][23] ),.IN2(\prod2[1][0][23] ),.IN4(\prod2[3][0][23] ),.S0(n368),.S1(n41),.Q(N152));
  MUX41X1 U145(.IN1(\prod2[0][1][6] ),.IN3(\prod2[2][1][6] ),.IN2(\prod2[1][1][6] ),.IN4(\prod2[3][1][6] ),.S0(n367),.S1(n369),.Q(N193));
  MUX41X1 U146(.IN1(\prod2[0][1][7] ),.IN3(\prod2[2][1][7] ),.IN2(\prod2[1][1][7] ),.IN4(\prod2[3][1][7] ),.S0(n367),.S1(n369),.Q(N192));
  MUX41X1 U147(.IN1(\prod2[0][1][8] ),.IN3(\prod2[2][1][8] ),.IN2(\prod2[1][1][8] ),.IN4(\prod2[3][1][8] ),.S0(n367),.S1(n369),.Q(N191));
  MUX41X1 U148(.IN1(\prod2[0][1][9] ),.IN3(\prod2[2][1][9] ),.IN2(\prod2[1][1][9] ),.IN4(\prod2[3][1][9] ),.S0(n367),.S1(n369),.Q(N190));
  MUX41X1 U149(.IN1(\prod2[0][1][10] ),.IN3(\prod2[2][1][10] ),.IN2(\prod2[1][1][10] ),.IN4(\prod2[3][1][10] ),.S0(n367),.S1(n369),.Q(N189));
  MUX41X1 U150(.IN1(\prod2[0][1][11] ),.IN3(\prod2[2][1][11] ),.IN2(\prod2[1][1][11] ),.IN4(\prod2[3][1][11] ),.S0(n367),.S1(n369),.Q(N188));
  MUX41X1 U151(.IN1(\prod2[0][1][12] ),.IN3(\prod2[2][1][12] ),.IN2(\prod2[1][1][12] ),.IN4(\prod2[3][1][12] ),.S0(n367),.S1(n369),.Q(N187));
  MUX41X1 U152(.IN1(\prod2[0][1][13] ),.IN3(\prod2[2][1][13] ),.IN2(\prod2[1][1][13] ),.IN4(\prod2[3][1][13] ),.S0(n367),.S1(n369),.Q(N186));
  MUX41X1 U153(.IN1(\prod2[0][1][14] ),.IN3(\prod2[2][1][14] ),.IN2(\prod2[1][1][14] ),.IN4(\prod2[3][1][14] ),.S0(n367),.S1(n369),.Q(N185));
  MUX41X1 U154(.IN1(\prod2[0][1][15] ),.IN3(\prod2[2][1][15] ),.IN2(\prod2[1][1][15] ),.IN4(\prod2[3][1][15] ),.S0(n367),.S1(n369),.Q(N184));
  MUX41X1 U155(.IN1(\prod2[0][1][16] ),.IN3(\prod2[2][1][16] ),.IN2(\prod2[1][1][16] ),.IN4(\prod2[3][1][16] ),.S0(n367),.S1(n369),.Q(N183));
  MUX41X1 U156(.IN1(\prod2[0][1][17] ),.IN3(\prod2[2][1][17] ),.IN2(\prod2[1][1][17] ),.IN4(\prod2[3][1][17] ),.S0(n367),.S1(n369),.Q(N182));
  MUX41X1 U157(.IN1(\prod2[0][2][6] ),.IN3(\prod2[2][2][6] ),.IN2(\prod2[1][2][6] ),.IN4(\prod2[3][2][6] ),.S0(n366),.S1(n370),.Q(N256));
  MUX41X1 U158(.IN1(\prod2[0][2][7] ),.IN3(\prod2[2][2][7] ),.IN2(\prod2[1][2][7] ),.IN4(\prod2[3][2][7] ),.S0(n366),.S1(n370),.Q(N257));
  MUX41X1 U159(.IN1(\prod2[0][2][8] ),.IN3(\prod2[2][2][8] ),.IN2(\prod2[1][2][8] ),.IN4(\prod2[3][2][8] ),.S0(n366),.S1(n370),.Q(N258));
  MUX41X1 U160(.IN1(\prod2[0][2][9] ),.IN3(\prod2[2][2][9] ),.IN2(\prod2[1][2][9] ),.IN4(\prod2[3][2][9] ),.S0(n366),.S1(n370),.Q(N259));
  MUX41X1 U161(.IN1(\prod2[0][2][10] ),.IN3(\prod2[2][2][10] ),.IN2(\prod2[1][2][10] ),.IN4(\prod2[3][2][10] ),.S0(n366),.S1(n370),.Q(N260));
  MUX41X1 U162(.IN1(\prod2[0][2][11] ),.IN3(\prod2[2][2][11] ),.IN2(\prod2[1][2][11] ),.IN4(\prod2[3][2][11] ),.S0(n366),.S1(n370),.Q(N261));
  MUX41X1 U163(.IN1(\prod2[0][2][12] ),.IN3(\prod2[2][2][12] ),.IN2(\prod2[1][2][12] ),.IN4(\prod2[3][2][12] ),.S0(n366),.S1(n370),.Q(N237));
  MUX41X1 U164(.IN1(\prod2[0][2][13] ),.IN3(\prod2[2][2][13] ),.IN2(\prod2[1][2][13] ),.IN4(\prod2[3][2][13] ),.S0(n366),.S1(n370),.Q(N236));
  MUX41X1 U165(.IN1(\prod2[0][2][14] ),.IN3(\prod2[2][2][14] ),.IN2(\prod2[1][2][14] ),.IN4(\prod2[3][2][14] ),.S0(n366),.S1(n370),.Q(N235));
  MUX41X1 U166(.IN1(\prod2[0][2][15] ),.IN3(\prod2[2][2][15] ),.IN2(\prod2[1][2][15] ),.IN4(\prod2[3][2][15] ),.S0(n366),.S1(n370),.Q(N234));
  MUX41X1 U167(.IN1(\prod2[0][2][16] ),.IN3(\prod2[2][2][16] ),.IN2(\prod2[1][2][16] ),.IN4(\prod2[3][2][16] ),.S0(n366),.S1(n370),.Q(N233));
  MUX41X1 U168(.IN1(\prod2[0][2][17] ),.IN3(\prod2[2][2][17] ),.IN2(\prod2[1][2][17] ),.IN4(\prod2[3][2][17] ),.S0(n366),.S1(n370),.Q(N232));
  MUX41X1 U169(.IN1(\prod2[0][3][0] ),.IN3(\prod2[2][3][0] ),.IN2(\prod2[1][3][0] ),.IN4(\prod2[3][3][0] ),.S0(n365),.S1(n371),.Q(N200));
  MUX41X1 U170(.IN1(\prod2[0][3][1] ),.IN3(\prod2[2][3][1] ),.IN2(\prod2[1][3][1] ),.IN4(\prod2[3][3][1] ),.S0(n365),.S1(n371),.Q(N201));
  MUX41X1 U171(.IN1(\prod2[0][3][2] ),.IN3(\prod2[2][3][2] ),.IN2(\prod2[1][3][2] ),.IN4(\prod2[3][3][2] ),.S0(n365),.S1(n371),.Q(N202));
  MUX41X1 U172(.IN1(\prod2[0][3][3] ),.IN3(\prod2[2][3][3] ),.IN2(\prod2[1][3][3] ),.IN4(\prod2[3][3][3] ),.S0(n365),.S1(n371),.Q(N203));
  MUX41X1 U173(.IN1(\prod2[0][3][4] ),.IN3(\prod2[2][3][4] ),.IN2(\prod2[1][3][4] ),.IN4(\prod2[3][3][4] ),.S0(n365),.S1(n371),.Q(N204));
  MUX41X1 U174(.IN1(\prod2[0][3][5] ),.IN3(\prod2[2][3][5] ),.IN2(\prod2[1][3][5] ),.IN4(\prod2[3][3][5] ),.S0(n365),.S1(n371),.Q(N205));
  MUX41X1 U175(.IN1(\prod2[0][3][6] ),.IN3(\prod2[2][3][6] ),.IN2(\prod2[1][3][6] ),.IN4(\prod2[3][3][6] ),.S0(n365),.S1(n371),.Q(N293));
  MUX41X1 U176(.IN1(\prod2[0][3][7] ),.IN3(\prod2[2][3][7] ),.IN2(\prod2[1][3][7] ),.IN4(\prod2[3][3][7] ),.S0(n365),.S1(n371),.Q(N292));
  MUX41X1 U177(.IN1(\prod2[0][3][8] ),.IN3(\prod2[2][3][8] ),.IN2(\prod2[1][3][8] ),.IN4(\prod2[3][3][8] ),.S0(n365),.S1(n371),.Q(N291));
  MUX41X1 U178(.IN1(\prod2[0][3][9] ),.IN3(\prod2[2][3][9] ),.IN2(\prod2[1][3][9] ),.IN4(\prod2[3][3][9] ),.S0(n365),.S1(n371),.Q(N290));
  MUX41X1 U179(.IN1(\prod2[0][3][10] ),.IN3(\prod2[2][3][10] ),.IN2(\prod2[1][3][10] ),.IN4(\prod2[3][3][10] ),.S0(n365),.S1(n371),.Q(N289));
  MUX41X1 U180(.IN1(\prod2[0][3][11] ),.IN3(\prod2[2][3][11] ),.IN2(\prod2[1][3][11] ),.IN4(\prod2[3][3][11] ),.S0(n365),.S1(n371),.Q(N288));
endmodule
module serial_mul_DW_mult_uns_0_inj (a,b,product);
input [47:0] a ;
output [48:0] product ;
input b ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
// instances
  NBUFFX2 U103(.INP(b),.Z(n154));
  NBUFFX2 U104(.INP(b),.Z(n155));
  NBUFFX2 U105(.INP(b),.Z(n156));
  NBUFFX2 U106(.INP(b),.Z(n157));
  AND2X1 U107(.IN1(n157),.IN2(a[9:9]),.Q(product[9:9]));
  AND2X1 U108(.IN1(a[8:8]),.IN2(n157),.Q(product[8:8]));
  AND2X1 U109(.IN1(a[7:7]),.IN2(n157),.Q(product[7:7]));
  AND2X1 U110(.IN1(a[6:6]),.IN2(n157),.Q(product[6:6]));
  AND2X1 U111(.IN1(a[5:5]),.IN2(n157),.Q(product[5:5]));
  AND2X1 U112(.IN1(a[4:4]),.IN2(n157),.Q(product[4:4]));
  AND2X1 U113(.IN1(a[47:47]),.IN2(n157),.Q(product[47:47]));
  AND2X1 U114(.IN1(a[46:46]),.IN2(n157),.Q(product[46:46]));
  AND2X1 U115(.IN1(a[45:45]),.IN2(n157),.Q(product[45:45]));
  AND2X1 U116(.IN1(a[44:44]),.IN2(n157),.Q(product[44:44]));
  AND2X1 U117(.IN1(a[43:43]),.IN2(n157),.Q(product[43:43]));
  AND2X1 U118(.IN1(a[42:42]),.IN2(n157),.Q(product[42:42]));
  AND2X1 U119(.IN1(a[41:41]),.IN2(n156),.Q(product[41:41]));
  AND2X1 U120(.IN1(a[40:40]),.IN2(n156),.Q(product[40:40]));
  AND2X1 U121(.IN1(a[3:3]),.IN2(n156),.Q(product[3:3]));
  AND2X1 U122(.IN1(a[39:39]),.IN2(n156),.Q(product[39:39]));
  AND2X1 U123(.IN1(a[38:38]),.IN2(n156),.Q(product[38:38]));
  AND2X1 U124(.IN1(a[37:37]),.IN2(n156),.Q(product[37:37]));
  AND2X1 U125(.IN1(a[36:36]),.IN2(n156),.Q(product[36:36]));
  AND2X1 U126(.IN1(a[35:35]),.IN2(n156),.Q(product[35:35]));
  AND2X1 U127(.IN1(a[34:34]),.IN2(n156),.Q(product[34:34]));
  AND2X1 U128(.IN1(a[33:33]),.IN2(n156),.Q(product[33:33]));
  AND2X1 U129(.IN1(a[32:32]),.IN2(n156),.Q(product[32:32]));
  AND2X1 U130(.IN1(a[31:31]),.IN2(n156),.Q(product[31:31]));
  AND2X1 U131(.IN1(a[30:30]),.IN2(n155),.Q(product[30:30]));
  AND2X1 U132(.IN1(a[2:2]),.IN2(n155),.Q(product[2:2]));
  AND2X1 U133(.IN1(a[29:29]),.IN2(n155),.Q(product[29:29]));
  AND2X1 U134(.IN1(a[28:28]),.IN2(n155),.Q(product[28:28]));
  AND2X1 U135(.IN1(a[27:27]),.IN2(n155),.Q(product[27:27]));
  AND2X1 U136(.IN1(a[26:26]),.IN2(n155),.Q(product[26:26]));
  AND2X1 U137(.IN1(a[25:25]),.IN2(n155),.Q(product[25:25]));
  AND2X1 U138(.IN1(a[24:24]),.IN2(n155),.Q(product[24:24]));
  AND2X1 U139(.IN1(a[23:23]),.IN2(n155),.Q(product[23:23]));
  AND2X1 U140(.IN1(a[22:22]),.IN2(n155),.Q(product[22:22]));
  AND2X1 U141(.IN1(a[21:21]),.IN2(n155),.Q(product[21:21]));
  AND2X1 U142(.IN1(a[20:20]),.IN2(n155),.Q(product[20:20]));
  AND2X1 U143(.IN1(a[1:1]),.IN2(n154),.Q(product[1:1]));
  AND2X1 U144(.IN1(a[19:19]),.IN2(n154),.Q(product[19:19]));
  AND2X1 U145(.IN1(a[18:18]),.IN2(n154),.Q(product[18:18]));
  AND2X1 U146(.IN1(a[17:17]),.IN2(n154),.Q(product[17:17]));
  AND2X1 U147(.IN1(a[16:16]),.IN2(n154),.Q(product[16:16]));
  AND2X1 U148(.IN1(a[15:15]),.IN2(n154),.Q(product[15:15]));
  AND2X1 U149(.IN1(a[14:14]),.IN2(n154),.Q(product[14:14]));
  AND2X1 U150(.IN1(a[13:13]),.IN2(n154),.Q(product[13:13]));
  AND2X1 U151(.IN1(a[12:12]),.IN2(n154),.Q(product[12:12]));
  AND2X1 U152(.IN1(a[11:11]),.IN2(n154),.Q(product[11:11]));
  AND2X1 U153(.IN1(a[10:10]),.IN2(n154),.Q(product[10:10]));
  AND2X1 U154(.IN1(a[0:0]),.IN2(n154),.Q(product[0:0]));
endmodule
module serial_mul_DW01_add_0_inj (A,B,CI,SUM,CO);
input [47:0] A ;
input [47:0] B ;
output [47:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire [47:1] carry ;
// instances
  FADDX1 U1_46(.A(A[46:46]),.B(B[46:46]),.CI(carry[46:46]),.CO(carry[47:47]),.S(SUM[46:46]));
  FADDX1 U1_45(.A(A[45:45]),.B(B[45:45]),.CI(carry[45:45]),.CO(carry[46:46]),.S(SUM[45:45]));
  FADDX1 U1_44(.A(A[44:44]),.B(B[44:44]),.CI(carry[44:44]),.CO(carry[45:45]),.S(SUM[44:44]));
  FADDX1 U1_43(.A(A[43:43]),.B(B[43:43]),.CI(carry[43:43]),.CO(carry[44:44]),.S(SUM[43:43]));
  FADDX1 U1_42(.A(A[42:42]),.B(B[42:42]),.CI(carry[42:42]),.CO(carry[43:43]),.S(SUM[42:42]));
  FADDX1 U1_41(.A(A[41:41]),.B(B[41:41]),.CI(carry[41:41]),.CO(carry[42:42]),.S(SUM[41:41]));
  FADDX1 U1_40(.A(A[40:40]),.B(B[40:40]),.CI(carry[40:40]),.CO(carry[41:41]),.S(SUM[40:40]));
  FADDX1 U1_39(.A(A[39:39]),.B(B[39:39]),.CI(carry[39:39]),.CO(carry[40:40]),.S(SUM[39:39]));
  FADDX1 U1_38(.A(A[38:38]),.B(B[38:38]),.CI(carry[38:38]),.CO(carry[39:39]),.S(SUM[38:38]));
  FADDX1 U1_37(.A(A[37:37]),.B(B[37:37]),.CI(carry[37:37]),.CO(carry[38:38]),.S(SUM[37:37]));
  FADDX1 U1_36(.A(A[36:36]),.B(B[36:36]),.CI(carry[36:36]),.CO(carry[37:37]),.S(SUM[36:36]));
  FADDX1 U1_35(.A(A[35:35]),.B(B[35:35]),.CI(carry[35:35]),.CO(carry[36:36]),.S(SUM[35:35]));
  FADDX1 U1_34(.A(A[34:34]),.B(B[34:34]),.CI(carry[34:34]),.CO(carry[35:35]),.S(SUM[34:34]));
  FADDX1 U1_33(.A(A[33:33]),.B(B[33:33]),.CI(carry[33:33]),.CO(carry[34:34]),.S(SUM[33:33]));
  FADDX1 U1_32(.A(A[32:32]),.B(B[32:32]),.CI(carry[32:32]),.CO(carry[33:33]),.S(SUM[32:32]));
  FADDX1 U1_31(.A(A[31:31]),.B(B[31:31]),.CI(carry[31:31]),.CO(carry[32:32]),.S(SUM[31:31]));
  FADDX1 U1_30(.A(A[30:30]),.B(B[30:30]),.CI(carry[30:30]),.CO(carry[31:31]),.S(SUM[30:30]));
  FADDX1 U1_29(.A(A[29:29]),.B(B[29:29]),.CI(carry[29:29]),.CO(carry[30:30]),.S(SUM[29:29]));
  FADDX1 U1_28(.A(A[28:28]),.B(B[28:28]),.CI(carry[28:28]),.CO(carry[29:29]),.S(SUM[28:28]));
  FADDX1 U1_27(.A(A[27:27]),.B(B[27:27]),.CI(carry[27:27]),.CO(carry[28:28]),.S(SUM[27:27]));
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(carry[26:26]),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_25(.A(A[25:25]),.B(B[25:25]),.CI(carry[25:25]),.CO(carry[26:26]),.S(SUM[25:25]));
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(carry[24:24]),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(carry[13:13]),.CO(carry[14:14]),.S(SUM[13:13]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(carry[12:12]),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_11(.A(A[11:11]),.B(B[11:11]),.CI(carry[11:11]),.CO(carry[12:12]),.S(SUM[11:11]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(carry[10:10]),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_9(.A(A[9:9]),.B(B[9:9]),.CI(carry[9:9]),.CO(carry[10:10]),.S(SUM[9:9]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(carry[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  XOR3X1 U1_47(.IN1(A[47:47]),.IN2(B[47:47]),.IN3(carry[47:47]),.Q(SUM[47:47]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  XOR2X1 U2(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module serial_mul_inj (clk_i,fracta_i,fractb_i,signa_i,signb_i,start_i,fract_o,sign_o,ready_o);
input [23:0] fracta_i ;
input [23:0] fractb_i ;
output [47:0] fract_o ;
input clk_i ;
input signa_i ;
input signb_i ;
input start_i ;
output sign_o ;
output ready_o ;
wire s_start_i ;
wire s_sign_o ;
wire s_ready_o ;
wire s_state ;
wire \s_count[4]  ;
wire N1833 ;
wire N1834 ;
wire N1835 ;
wire N1836 ;
wire N2451 ;
wire N2453 ;
wire N2454 ;
wire N2455 ;
wire N2456 ;
wire N2457 ;
wire N2458 ;
wire N2459 ;
wire N2460 ;
wire N2461 ;
wire N2462 ;
wire N2463 ;
wire N2464 ;
wire N2465 ;
wire N2466 ;
wire N2467 ;
wire N2468 ;
wire N2469 ;
wire N2470 ;
wire N2471 ;
wire N2472 ;
wire N2473 ;
wire N2474 ;
wire N2475 ;
wire N2476 ;
wire N2484 ;
wire N2485 ;
wire N2486 ;
wire N2487 ;
wire N2488 ;
wire N2489 ;
wire N2490 ;
wire N2491 ;
wire N2492 ;
wire N2493 ;
wire N2494 ;
wire N2495 ;
wire N2496 ;
wire N2497 ;
wire N2498 ;
wire N2499 ;
wire N2500 ;
wire N2503 ;
wire N2504 ;
wire N2505 ;
wire N2506 ;
wire N2507 ;
wire N2508 ;
wire N2509 ;
wire N2510 ;
wire N2511 ;
wire N2512 ;
wire N2513 ;
wire N2514 ;
wire N2515 ;
wire N2516 ;
wire N2517 ;
wire N2518 ;
wire N2519 ;
wire N2520 ;
wire N2521 ;
wire N2522 ;
wire N2523 ;
wire N2524 ;
wire N2525 ;
wire N2526 ;
wire N2527 ;
wire N2528 ;
wire N2529 ;
wire N2530 ;
wire N2531 ;
wire N2532 ;
wire N2533 ;
wire N2534 ;
wire N2535 ;
wire N2536 ;
wire N2537 ;
wire N2538 ;
wire N2539 ;
wire N2540 ;
wire N2541 ;
wire N2542 ;
wire N2543 ;
wire N2544 ;
wire N2545 ;
wire N2546 ;
wire N2547 ;
wire N2548 ;
wire N2549 ;
wire N2550 ;
wire N2554 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire N2611 ;
wire N2610 ;
wire N2609 ;
wire N2608 ;
wire N2607 ;
wire N2606 ;
wire N2605 ;
wire N2604 ;
wire N2603 ;
wire N2602 ;
wire N2601 ;
wire N2600 ;
wire N2599 ;
wire N2598 ;
wire N2597 ;
wire N2596 ;
wire N2595 ;
wire N2594 ;
wire N2593 ;
wire N2592 ;
wire N2591 ;
wire N2590 ;
wire N2589 ;
wire N2588 ;
wire N2587 ;
wire N2586 ;
wire N2585 ;
wire N2584 ;
wire N2583 ;
wire N2582 ;
wire N2581 ;
wire N2580 ;
wire N2579 ;
wire N2578 ;
wire N2577 ;
wire N2576 ;
wire N2575 ;
wire N2574 ;
wire N2573 ;
wire N2572 ;
wire N2571 ;
wire N2570 ;
wire N2569 ;
wire N2568 ;
wire N2567 ;
wire N2566 ;
wire N2565 ;
wire N2564 ;
wire \add_118/carry[4]  ;
wire \add_118/carry[3]  ;
wire \add_118/carry[2]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n11 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire [23:0] s_fractb_i ;
wire [47:0] s_fract_o ;
wire [23:0] s_tem_prod ;
wire SYNOPSYS_UNCONNECTED__0 ;
// instances
  DFFX1 desc724(.D(fracta_i[23:23]),.CLK(clk_i),.QN(n28));
  DFFX1 desc725(.D(fracta_i[22:22]),.CLK(clk_i),.QN(n27));
  DFFX1 desc726(.D(fracta_i[21:21]),.CLK(clk_i),.QN(n26));
  DFFX1 desc727(.D(fracta_i[20:20]),.CLK(clk_i),.QN(n25));
  DFFX1 desc728(.D(fracta_i[19:19]),.CLK(clk_i),.QN(n23));
  DFFX1 desc729(.D(fracta_i[18:18]),.CLK(clk_i),.QN(n22));
  DFFX1 desc730(.D(fracta_i[17:17]),.CLK(clk_i),.QN(n21));
  DFFX1 desc731(.D(fracta_i[16:16]),.CLK(clk_i),.QN(n20));
  DFFX1 desc732(.D(fracta_i[15:15]),.CLK(clk_i),.QN(n19));
  DFFX1 desc733(.D(fracta_i[14:14]),.CLK(clk_i),.QN(n18));
  DFFX1 desc734(.D(fracta_i[13:13]),.CLK(clk_i),.QN(n17));
  DFFX1 desc735(.D(fracta_i[12:12]),.CLK(clk_i),.QN(n16));
  DFFX1 desc736(.D(fracta_i[11:11]),.CLK(clk_i),.QN(n15));
  DFFX1 desc737(.D(fracta_i[10:10]),.CLK(clk_i),.QN(n14));
  DFFX1 desc738(.D(fracta_i[9:9]),.CLK(clk_i),.QN(n36));
  DFFX1 desc739(.D(fracta_i[8:8]),.CLK(clk_i),.QN(n35));
  DFFX1 desc740(.D(fracta_i[7:7]),.CLK(clk_i),.QN(n34));
  DFFX1 desc741(.D(fracta_i[6:6]),.CLK(clk_i),.QN(n33));
  DFFX1 desc742(.D(fracta_i[5:5]),.CLK(clk_i),.QN(n32));
  DFFX1 desc743(.D(fracta_i[4:4]),.CLK(clk_i),.QN(n31));
  DFFX1 desc744(.D(fracta_i[3:3]),.CLK(clk_i),.QN(n30));
  DFFX1 desc745(.D(fracta_i[2:2]),.CLK(clk_i),.QN(n29));
  DFFX1 desc746(.D(fracta_i[1:1]),.CLK(clk_i),.QN(n24));
  DFFX1 desc747(.D(fracta_i[0:0]),.CLK(clk_i),.QN(n13));
  DFFX1 desc748(.D(fractb_i[23:23]),.CLK(clk_i),.Q(s_fractb_i[23:23]));
  DFFX1 desc749(.D(fractb_i[22:22]),.CLK(clk_i),.Q(s_fractb_i[22:22]));
  DFFX1 desc750(.D(fractb_i[21:21]),.CLK(clk_i),.Q(s_fractb_i[21:21]));
  DFFX1 desc751(.D(fractb_i[20:20]),.CLK(clk_i),.Q(s_fractb_i[20:20]));
  DFFX1 desc752(.D(fractb_i[19:19]),.CLK(clk_i),.Q(s_fractb_i[19:19]));
  DFFX1 desc753(.D(fractb_i[18:18]),.CLK(clk_i),.Q(s_fractb_i[18:18]));
  DFFX1 desc754(.D(fractb_i[17:17]),.CLK(clk_i),.Q(s_fractb_i[17:17]));
  DFFX1 desc755(.D(fractb_i[16:16]),.CLK(clk_i),.Q(s_fractb_i[16:16]));
  DFFX1 desc756(.D(fractb_i[15:15]),.CLK(clk_i),.Q(s_fractb_i[15:15]));
  DFFX1 desc757(.D(fractb_i[14:14]),.CLK(clk_i),.Q(s_fractb_i[14:14]));
  DFFX1 desc758(.D(fractb_i[13:13]),.CLK(clk_i),.Q(s_fractb_i[13:13]));
  DFFX1 desc759(.D(fractb_i[12:12]),.CLK(clk_i),.Q(s_fractb_i[12:12]));
  DFFX1 desc760(.D(fractb_i[11:11]),.CLK(clk_i),.Q(s_fractb_i[11:11]));
  DFFX1 desc761(.D(fractb_i[10:10]),.CLK(clk_i),.Q(s_fractb_i[10:10]));
  DFFX1 desc762(.D(fractb_i[9:9]),.CLK(clk_i),.Q(s_fractb_i[9:9]));
  DFFX1 desc763(.D(fractb_i[8:8]),.CLK(clk_i),.Q(s_fractb_i[8:8]));
  DFFX1 desc764(.D(fractb_i[7:7]),.CLK(clk_i),.Q(s_fractb_i[7:7]));
  DFFX1 desc765(.D(fractb_i[6:6]),.CLK(clk_i),.Q(s_fractb_i[6:6]));
  DFFX1 desc766(.D(fractb_i[5:5]),.CLK(clk_i),.Q(s_fractb_i[5:5]));
  DFFX1 desc767(.D(fractb_i[4:4]),.CLK(clk_i),.Q(s_fractb_i[4:4]));
  DFFX1 desc768(.D(fractb_i[3:3]),.CLK(clk_i),.Q(s_fractb_i[3:3]));
  DFFX1 desc769(.D(fractb_i[2:2]),.CLK(clk_i),.Q(s_fractb_i[2:2]));
  DFFX1 desc770(.D(fractb_i[1:1]),.CLK(clk_i),.Q(s_fractb_i[1:1]));
  DFFX1 desc771(.D(fractb_i[0:0]),.CLK(clk_i),.Q(s_fractb_i[0:0]));
  DFFX1 s_start_i_reg(.D(start_i),.CLK(clk_i),.Q(s_start_i),.QN(n93));
  DFFX1 sign_o_reg(.D(s_sign_o),.CLK(clk_i),.Q(sign_o));
  DFFX1 desc772(.D(n91),.CLK(clk_i),.QN(n4));
  DFFX1 s_state_reg(.D(n90),.CLK(clk_i),.Q(s_state),.QN(n2));
  DFFX1 s_ready_o_reg(.D(n85),.CLK(clk_i),.Q(s_ready_o));
  DFFX1 ready_o_reg(.D(s_ready_o),.CLK(clk_i),.Q(ready_o));
  DFFX1 desc773(.D(n89),.CLK(clk_i),.Q(n1),.QN(n5));
  DFFX1 desc774(.D(n88),.CLK(clk_i),.QN(n3));
  DFFX1 desc775(.D(n87),.CLK(clk_i),.QN(n92));
  DFFX1 desc776(.D(n86),.CLK(clk_i),.Q(\s_count[4] ),.QN(n11));
  DFFX1 desc777(.D(n84),.CLK(clk_i),.Q(s_fract_o[47:47]));
  DFFX1 desc778(.D(s_fract_o[47:47]),.CLK(clk_i),.Q(fract_o[47:47]));
  DFFX1 desc779(.D(n83),.CLK(clk_i),.Q(s_fract_o[46:46]));
  DFFX1 desc780(.D(s_fract_o[46:46]),.CLK(clk_i),.Q(fract_o[46:46]));
  DFFX1 desc781(.D(n82),.CLK(clk_i),.Q(s_fract_o[45:45]));
  DFFX1 desc782(.D(s_fract_o[45:45]),.CLK(clk_i),.Q(fract_o[45:45]));
  DFFX1 desc783(.D(n81),.CLK(clk_i),.Q(s_fract_o[44:44]));
  DFFX1 desc784(.D(s_fract_o[44:44]),.CLK(clk_i),.Q(fract_o[44:44]));
  DFFX1 desc785(.D(n80),.CLK(clk_i),.Q(s_fract_o[43:43]));
  DFFX1 desc786(.D(s_fract_o[43:43]),.CLK(clk_i),.Q(fract_o[43:43]));
  DFFX1 desc787(.D(n79),.CLK(clk_i),.Q(s_fract_o[42:42]));
  DFFX1 desc788(.D(s_fract_o[42:42]),.CLK(clk_i),.Q(fract_o[42:42]));
  DFFX1 desc789(.D(n78),.CLK(clk_i),.Q(s_fract_o[41:41]));
  DFFX1 desc790(.D(s_fract_o[41:41]),.CLK(clk_i),.Q(fract_o[41:41]));
  DFFX1 desc791(.D(n77),.CLK(clk_i),.Q(s_fract_o[40:40]));
  DFFX1 desc792(.D(s_fract_o[40:40]),.CLK(clk_i),.Q(fract_o[40:40]));
  DFFX1 desc793(.D(n76),.CLK(clk_i),.Q(s_fract_o[39:39]));
  DFFX1 desc794(.D(s_fract_o[39:39]),.CLK(clk_i),.Q(fract_o[39:39]));
  DFFX1 desc795(.D(n75),.CLK(clk_i),.Q(s_fract_o[38:38]));
  DFFX1 desc796(.D(s_fract_o[38:38]),.CLK(clk_i),.Q(fract_o[38:38]));
  DFFX1 desc797(.D(n74),.CLK(clk_i),.Q(s_fract_o[37:37]));
  DFFX1 desc798(.D(s_fract_o[37:37]),.CLK(clk_i),.Q(fract_o[37:37]));
  DFFX1 desc799(.D(n73),.CLK(clk_i),.Q(s_fract_o[36:36]));
  DFFX1 desc800(.D(s_fract_o[36:36]),.CLK(clk_i),.Q(fract_o[36:36]));
  DFFX1 desc801(.D(n72),.CLK(clk_i),.Q(s_fract_o[35:35]));
  DFFX1 desc802(.D(s_fract_o[35:35]),.CLK(clk_i),.Q(fract_o[35:35]));
  DFFX1 desc803(.D(n71),.CLK(clk_i),.Q(s_fract_o[34:34]));
  DFFX1 desc804(.D(s_fract_o[34:34]),.CLK(clk_i),.Q(fract_o[34:34]));
  DFFX1 desc805(.D(n70),.CLK(clk_i),.Q(s_fract_o[33:33]));
  DFFX1 desc806(.D(s_fract_o[33:33]),.CLK(clk_i),.Q(fract_o[33:33]));
  DFFX1 desc807(.D(n69),.CLK(clk_i),.Q(s_fract_o[32:32]));
  DFFX1 desc808(.D(s_fract_o[32:32]),.CLK(clk_i),.Q(fract_o[32:32]));
  DFFX1 desc809(.D(n68),.CLK(clk_i),.Q(s_fract_o[31:31]));
  DFFX1 desc810(.D(s_fract_o[31:31]),.CLK(clk_i),.Q(fract_o[31:31]));
  DFFX1 desc811(.D(n67),.CLK(clk_i),.Q(s_fract_o[30:30]));
  DFFX1 desc812(.D(s_fract_o[30:30]),.CLK(clk_i),.Q(fract_o[30:30]));
  DFFX1 desc813(.D(n66),.CLK(clk_i),.Q(s_fract_o[29:29]));
  DFFX1 desc814(.D(s_fract_o[29:29]),.CLK(clk_i),.Q(fract_o[29:29]));
  DFFX1 desc815(.D(n65),.CLK(clk_i),.Q(s_fract_o[28:28]));
  DFFX1 desc816(.D(s_fract_o[28:28]),.CLK(clk_i),.Q(fract_o[28:28]));
  DFFX1 desc817(.D(n64),.CLK(clk_i),.Q(s_fract_o[27:27]));
  DFFX1 desc818(.D(s_fract_o[27:27]),.CLK(clk_i),.Q(fract_o[27:27]));
  DFFX1 desc819(.D(n63),.CLK(clk_i),.Q(s_fract_o[26:26]));
  DFFX1 desc820(.D(s_fract_o[26:26]),.CLK(clk_i),.Q(fract_o[26:26]));
  DFFX1 desc821(.D(n62),.CLK(clk_i),.Q(s_fract_o[25:25]));
  DFFX1 desc822(.D(s_fract_o[25:25]),.CLK(clk_i),.Q(fract_o[25:25]));
  DFFX1 desc823(.D(n61),.CLK(clk_i),.Q(s_fract_o[24:24]));
  DFFX1 desc824(.D(s_fract_o[24:24]),.CLK(clk_i),.Q(fract_o[24:24]));
  DFFX1 desc825(.D(n60),.CLK(clk_i),.Q(s_fract_o[23:23]));
  DFFX1 desc826(.D(s_fract_o[23:23]),.CLK(clk_i),.Q(fract_o[23:23]));
  DFFX1 desc827(.D(n59),.CLK(clk_i),.Q(s_fract_o[22:22]));
  DFFX1 desc828(.D(s_fract_o[22:22]),.CLK(clk_i),.Q(fract_o[22:22]));
  DFFX1 desc829(.D(n58),.CLK(clk_i),.Q(s_fract_o[21:21]));
  DFFX1 desc830(.D(s_fract_o[21:21]),.CLK(clk_i),.Q(fract_o[21:21]));
  DFFX1 desc831(.D(n57),.CLK(clk_i),.Q(s_fract_o[20:20]));
  DFFX1 desc832(.D(s_fract_o[20:20]),.CLK(clk_i),.Q(fract_o[20:20]));
  DFFX1 desc833(.D(n56),.CLK(clk_i),.Q(s_fract_o[19:19]));
  DFFX1 desc834(.D(s_fract_o[19:19]),.CLK(clk_i),.Q(fract_o[19:19]));
  DFFX1 desc835(.D(n55),.CLK(clk_i),.Q(s_fract_o[18:18]));
  DFFX1 desc836(.D(s_fract_o[18:18]),.CLK(clk_i),.Q(fract_o[18:18]));
  DFFX1 desc837(.D(n54),.CLK(clk_i),.Q(s_fract_o[17:17]));
  DFFX1 desc838(.D(s_fract_o[17:17]),.CLK(clk_i),.Q(fract_o[17:17]));
  DFFX1 desc839(.D(n53),.CLK(clk_i),.Q(s_fract_o[16:16]));
  DFFX1 desc840(.D(s_fract_o[16:16]),.CLK(clk_i),.Q(fract_o[16:16]));
  DFFX1 desc841(.D(n52),.CLK(clk_i),.Q(s_fract_o[15:15]));
  DFFX1 desc842(.D(s_fract_o[15:15]),.CLK(clk_i),.Q(fract_o[15:15]));
  DFFX1 desc843(.D(n51),.CLK(clk_i),.Q(s_fract_o[14:14]));
  DFFX1 desc844(.D(s_fract_o[14:14]),.CLK(clk_i),.Q(fract_o[14:14]));
  DFFX1 desc845(.D(n50),.CLK(clk_i),.Q(s_fract_o[13:13]));
  DFFX1 desc846(.D(s_fract_o[13:13]),.CLK(clk_i),.Q(fract_o[13:13]));
  DFFX1 desc847(.D(n49),.CLK(clk_i),.Q(s_fract_o[12:12]));
  DFFX1 desc848(.D(s_fract_o[12:12]),.CLK(clk_i),.Q(fract_o[12:12]));
  DFFX1 desc849(.D(n48),.CLK(clk_i),.Q(s_fract_o[11:11]));
  DFFX1 desc850(.D(s_fract_o[11:11]),.CLK(clk_i),.Q(fract_o[11:11]));
  DFFX1 desc851(.D(n47),.CLK(clk_i),.Q(s_fract_o[10:10]));
  DFFX1 desc852(.D(s_fract_o[10:10]),.CLK(clk_i),.Q(fract_o[10:10]));
  DFFX1 desc853(.D(n46),.CLK(clk_i),.Q(s_fract_o[9:9]));
  DFFX1 desc854(.D(s_fract_o[9:9]),.CLK(clk_i),.Q(fract_o[9:9]));
  DFFX1 desc855(.D(n45),.CLK(clk_i),.Q(s_fract_o[8:8]));
  DFFX1 desc856(.D(s_fract_o[8:8]),.CLK(clk_i),.Q(fract_o[8:8]));
  DFFX1 desc857(.D(n44),.CLK(clk_i),.Q(s_fract_o[7:7]));
  DFFX1 desc858(.D(s_fract_o[7:7]),.CLK(clk_i),.Q(fract_o[7:7]));
  DFFX1 desc859(.D(n43),.CLK(clk_i),.Q(s_fract_o[6:6]));
  DFFX1 desc860(.D(s_fract_o[6:6]),.CLK(clk_i),.Q(fract_o[6:6]));
  DFFX1 desc861(.D(n42),.CLK(clk_i),.Q(s_fract_o[5:5]));
  DFFX1 desc862(.D(s_fract_o[5:5]),.CLK(clk_i),.Q(fract_o[5:5]));
  DFFX1 desc863(.D(n41),.CLK(clk_i),.Q(s_fract_o[4:4]));
  DFFX1 desc864(.D(s_fract_o[4:4]),.CLK(clk_i),.Q(fract_o[4:4]));
  DFFX1 desc865(.D(n40),.CLK(clk_i),.Q(s_fract_o[3:3]));
  DFFX1 desc866(.D(s_fract_o[3:3]),.CLK(clk_i),.Q(fract_o[3:3]));
  DFFX1 desc867(.D(n39),.CLK(clk_i),.Q(s_fract_o[2:2]));
  DFFX1 desc868(.D(s_fract_o[2:2]),.CLK(clk_i),.Q(fract_o[2:2]));
  DFFX1 desc869(.D(n38),.CLK(clk_i),.Q(s_fract_o[1:1]));
  DFFX1 desc870(.D(s_fract_o[1:1]),.CLK(clk_i),.Q(fract_o[1:1]));
  DFFX1 desc871(.D(n37),.CLK(clk_i),.Q(s_fract_o[0:0]));
  DFFX1 desc872(.D(s_fract_o[0:0]),.CLK(clk_i),.Q(fract_o[0:0]));
  XOR2X1 U29(.IN1(signb_i),.IN2(signa_i),.Q(s_sign_o));
  AO22X1 U30(.IN1(s_fract_o[0:0]),.IN2(n114),.IN3(n110),.IN4(N2503),.Q(n37));
  AO22X1 U31(.IN1(s_fract_o[1:1]),.IN2(n2),.IN3(N2504),.IN4(n112),.Q(n38));
  AO22X1 U32(.IN1(s_fract_o[2:2]),.IN2(n113),.IN3(N2505),.IN4(n112),.Q(n39));
  AO22X1 U33(.IN1(s_fract_o[3:3]),.IN2(n114),.IN3(N2506),.IN4(n112),.Q(n40));
  AO22X1 U34(.IN1(s_fract_o[4:4]),.IN2(n2),.IN3(N2507),.IN4(n112),.Q(n41));
  AO22X1 U35(.IN1(s_fract_o[5:5]),.IN2(n2),.IN3(N2508),.IN4(n112),.Q(n42));
  AO22X1 U36(.IN1(s_fract_o[6:6]),.IN2(n114),.IN3(N2509),.IN4(n112),.Q(n43));
  AO22X1 U37(.IN1(s_fract_o[7:7]),.IN2(n113),.IN3(N2510),.IN4(n112),.Q(n44));
  AO22X1 U38(.IN1(s_fract_o[8:8]),.IN2(n113),.IN3(N2511),.IN4(n112),.Q(n45));
  AO22X1 U39(.IN1(s_fract_o[9:9]),.IN2(n2),.IN3(N2512),.IN4(n112),.Q(n46));
  AO22X1 U40(.IN1(s_fract_o[10:10]),.IN2(n114),.IN3(N2513),.IN4(n112),.Q(n47));
  AO22X1 U41(.IN1(s_fract_o[11:11]),.IN2(n2),.IN3(N2514),.IN4(n112),.Q(n48));
  AO22X1 U42(.IN1(s_fract_o[12:12]),.IN2(n114),.IN3(N2515),.IN4(n111),.Q(n49));
  AO22X1 U43(.IN1(s_fract_o[13:13]),.IN2(n113),.IN3(N2516),.IN4(n111),.Q(n50));
  AO22X1 U44(.IN1(s_fract_o[14:14]),.IN2(n2),.IN3(N2517),.IN4(n111),.Q(n51));
  AO22X1 U45(.IN1(s_fract_o[15:15]),.IN2(n2),.IN3(N2518),.IN4(n111),.Q(n52));
  AO22X1 U46(.IN1(s_fract_o[16:16]),.IN2(n114),.IN3(N2519),.IN4(n111),.Q(n53));
  AO22X1 U47(.IN1(s_fract_o[17:17]),.IN2(n113),.IN3(N2520),.IN4(n111),.Q(n54));
  AO22X1 U48(.IN1(s_fract_o[18:18]),.IN2(n2),.IN3(N2521),.IN4(n111),.Q(n55));
  AO22X1 U49(.IN1(s_fract_o[19:19]),.IN2(n114),.IN3(N2522),.IN4(n111),.Q(n56));
  AO22X1 U50(.IN1(s_fract_o[20:20]),.IN2(n2),.IN3(N2523),.IN4(n111),.Q(n57));
  AO22X1 U51(.IN1(s_fract_o[21:21]),.IN2(n114),.IN3(N2524),.IN4(n111),.Q(n58));
  AO22X1 U52(.IN1(s_fract_o[22:22]),.IN2(n113),.IN3(N2525),.IN4(n111),.Q(n59));
  AO22X1 U53(.IN1(s_fract_o[23:23]),.IN2(n113),.IN3(N2526),.IN4(n111),.Q(n60));
  AO22X1 U54(.IN1(s_fract_o[24:24]),.IN2(n113),.IN3(N2527),.IN4(n110),.Q(n61));
  AO22X1 U55(.IN1(s_fract_o[25:25]),.IN2(n114),.IN3(N2528),.IN4(n110),.Q(n62));
  AO22X1 U56(.IN1(s_fract_o[26:26]),.IN2(n113),.IN3(N2529),.IN4(n110),.Q(n63));
  AO22X1 U57(.IN1(s_fract_o[27:27]),.IN2(n2),.IN3(N2530),.IN4(n110),.Q(n64));
  AO22X1 U58(.IN1(s_fract_o[28:28]),.IN2(n113),.IN3(N2531),.IN4(n110),.Q(n65));
  AO22X1 U59(.IN1(s_fract_o[29:29]),.IN2(n113),.IN3(N2532),.IN4(n110),.Q(n66));
  AO22X1 U60(.IN1(s_fract_o[30:30]),.IN2(n113),.IN3(N2533),.IN4(n110),.Q(n67));
  AO22X1 U61(.IN1(s_fract_o[31:31]),.IN2(n113),.IN3(N2534),.IN4(n110),.Q(n68));
  AO22X1 U62(.IN1(s_fract_o[32:32]),.IN2(n113),.IN3(N2535),.IN4(n110),.Q(n69));
  AO22X1 U63(.IN1(s_fract_o[33:33]),.IN2(n113),.IN3(N2536),.IN4(n110),.Q(n70));
  AO22X1 U64(.IN1(s_fract_o[34:34]),.IN2(n113),.IN3(N2537),.IN4(n110),.Q(n71));
  AO22X1 U65(.IN1(s_fract_o[35:35]),.IN2(n113),.IN3(N2538),.IN4(n109),.Q(n72));
  AO22X1 U66(.IN1(s_fract_o[36:36]),.IN2(n113),.IN3(N2539),.IN4(n110),.Q(n73));
  AO22X1 U67(.IN1(s_fract_o[37:37]),.IN2(n114),.IN3(N2540),.IN4(n109),.Q(n74));
  AO22X1 U68(.IN1(s_fract_o[38:38]),.IN2(n114),.IN3(N2541),.IN4(n109),.Q(n75));
  AO22X1 U69(.IN1(s_fract_o[39:39]),.IN2(n114),.IN3(N2542),.IN4(n109),.Q(n76));
  AO22X1 U70(.IN1(s_fract_o[40:40]),.IN2(n114),.IN3(N2543),.IN4(n109),.Q(n77));
  AO22X1 U71(.IN1(s_fract_o[41:41]),.IN2(n114),.IN3(N2544),.IN4(n109),.Q(n78));
  AO22X1 U72(.IN1(s_fract_o[42:42]),.IN2(n114),.IN3(N2545),.IN4(n109),.Q(n79));
  AO22X1 U73(.IN1(s_fract_o[43:43]),.IN2(n114),.IN3(N2546),.IN4(n109),.Q(n80));
  AO22X1 U74(.IN1(s_fract_o[44:44]),.IN2(n114),.IN3(N2547),.IN4(n109),.Q(n81));
  AO22X1 U75(.IN1(s_fract_o[45:45]),.IN2(n114),.IN3(N2548),.IN4(n109),.Q(n82));
  AO22X1 U76(.IN1(s_fract_o[46:46]),.IN2(n115),.IN3(N2549),.IN4(n109),.Q(n83));
  AO22X1 U77(.IN1(s_fract_o[47:47]),.IN2(n115),.IN3(N2550),.IN4(n109),.Q(n84));
  AO22X1 U78(.IN1(n162),.IN2(n93),.IN3(s_ready_o),.IN4(n6),.Q(n85));
  AO22X1 U80(.IN1(n7),.IN2(n106),.IN3(N1836),.IN4(n8),.Q(n86));
  AO22X1 U81(.IN1(n103),.IN2(n7),.IN3(N1835),.IN4(n8),.Q(n87));
  AO22X1 U82(.IN1(n7),.IN2(n101),.IN3(N1834),.IN4(n8),.Q(n88));
  AO22X1 U83(.IN1(n7),.IN2(n1),.IN3(N1833),.IN4(n8),.Q(n89));
  AO21X1 U84(.IN1(n112),.IN2(n9),.IN3(s_start_i),.Q(n90));
  AO22X1 U85(.IN1(n7),.IN2(n97),.IN3(n4),.IN4(n8),.Q(n91));
  NOR3X0 U86(.IN1(n7),.IN2(s_start_i),.IN3(n162),.QN(n8));
  AND3X1 U88(.IN1(n93),.IN2(n115),.IN3(n9),.Q(n7));
  NAND4X0 U89(.IN1(n106),.IN2(n101),.IN3(n10),.IN4(n1),.QN(n9));
  OR4X1 U94(.IN1(n97),.IN2(n1),.IN3(n12),.IN4(n101),.Q(N2554));
  OR2X1 U95(.IN1(n106),.IN2(n102),.Q(n12));
  serial_mul_DW_mult_uns_0_inj mult_add_137_aco(.a(s_fract_o),.b(N2554),.product({SYNOPSYS_UNCONNECTED__0,N2611,N2610,N2609,N2608,N2607,N2606,N2605,N2604,N2603,N2602,N2601,N2600,N2599,N2598,N2597,N2596,N2595,N2594,N2593,N2592,N2591,N2590,N2589,N2588,N2587,N2586,N2585,N2584,N2583,N2582,N2581,N2580,N2579,N2578,N2577,N2576,N2575,N2574,N2573,N2572,N2571,N2570,N2569,N2568,N2567,N2566,N2565,N2564}));
  serial_mul_DW01_add_0_inj add_137_aco(.A({N2500,N2499,N2498,N2497,N2496,N2495,N2494,N2493,N2492,N2491,N2490,N2489,N2488,N2487,N2486,N2485,N2484,n133,n128,n130,n126,n131,n127,n129,N2476,N2475,N2474,N2473,N2472,N2471,N2470,N2469,N2468,N2467,N2466,N2465,N2464,N2463,N2462,N2461,N2460,N2459,N2458,N2457,N2456,N2455,N2454,N2453}),.B({N2611,N2610,N2609,N2608,N2607,N2606,N2605,N2604,N2603,N2602,N2601,N2600,N2599,N2598,N2597,N2596,N2595,N2594,N2593,N2592,N2591,N2590,N2589,N2588,N2587,N2586,N2585,N2584,N2583,N2582,N2581,N2580,N2579,N2578,N2577,N2576,N2575,N2574,N2573,N2572,N2571,N2570,N2569,N2568,N2567,N2566,N2565,N2564}),.CI(1'b0),.SUM({N2550,N2549,N2548,N2547,N2546,N2545,N2544,N2543,N2542,N2541,N2540,N2539,N2538,N2537,N2536,N2535,N2534,N2533,N2532,N2531,N2530,N2529,N2528,N2527,N2526,N2525,N2524,N2523,N2522,N2521,N2520,N2519,N2518,N2517,N2516,N2515,N2514,N2513,N2512,N2511,N2510,N2509,N2508,N2507,N2506,N2505,N2504,N2503}));
  HADDX1 desc873(.A0(n1),.B0(n97),.C1(\add_118/carry[2] ),.SO(N1833));
  HADDX1 desc874(.A0(n100),.B0(\add_118/carry[2] ),.C1(\add_118/carry[3] ),.SO(N1834));
  HADDX1 desc875(.A0(n102),.B0(\add_118/carry[3] ),.C1(\add_118/carry[4] ),.SO(N1835));
  NAND2X0 U3(.IN1(n98),.IN2(n234),.QN(n252));
  NAND2X0 U4(.IN1(n257),.IN2(n99),.QN(n275));
  NAND2X0 U5(.IN1(n99),.IN2(n244),.QN(n268));
  NAND2X0 U6(.IN1(s_tem_prod[0:0]),.IN2(n4),.QN(n169));
  NBUFFX2 U7(.INP(n161),.Z(n94));
  NBUFFX2 U8(.INP(n161),.Z(n95));
  NOR2X0 U9(.IN1(n231),.IN2(n103),.QN(n196));
  NOR2X0 U10(.IN1(n236),.IN2(n103),.QN(n210));
  NOR2X0 U11(.IN1(n205),.IN2(n103),.QN(n256));
  NOR2X0 U12(.IN1(n209),.IN2(n103),.QN(n278));
  NOR2X0 U13(.IN1(n215),.IN2(n103),.QN(n287));
  NOR2X0 U14(.IN1(n220),.IN2(n103),.QN(n288));
  INVX0 U15(.INP(n179),.ZN(n158));
  NOR2X0 U16(.IN1(n225),.IN2(n103),.QN(n289));
  NOR2X0 U17(.IN1(n156),.IN2(n103),.QN(n290));
  INVX0 U18(.INP(n190),.ZN(n156));
  INVX0 U19(.INP(n176),.ZN(n154));
  INVX0 U20(.INP(n208),.ZN(n152));
  INVX0 U21(.INP(n173),.ZN(n150));
  INVX0 U22(.INP(n198),.ZN(n144));
  INVX0 U23(.INP(n187),.ZN(n148));
  INVX0 U24(.INP(n195),.ZN(n145));
  INVX0 U25(.INP(n199),.ZN(n143));
  INVX0 U26(.INP(n217),.ZN(n137));
  INVX0 U27(.INP(n228),.ZN(n125));
  INVX0 U28(.INP(n204),.ZN(n141));
  INVX0 U79(.INP(n214),.ZN(n138));
  INVX0 U87(.INP(n224),.ZN(n134));
  INVX0 U90(.INP(n219),.ZN(n136));
  INVX0 U91(.INP(n245),.ZN(n140));
  INVX0 U92(.INP(n257),.ZN(n132));
  INVX0 U93(.INP(n9),.ZN(n162));
  INVX0 U96(.INP(n92),.ZN(n102));
  INVX0 U97(.INP(n11),.ZN(n105));
  INVX0 U98(.INP(n5),.ZN(n98));
  INVX0 U99(.INP(n3),.ZN(n99));
  NAND2X0 U100(.IN1(n180),.IN2(n5),.QN(n200));
  INVX0 U101(.INP(N2451),.ZN(n161));
  INVX0 U102(.INP(n168),.ZN(n160));
  INVX0 U103(.INP(n4),.ZN(n96));
  NAND2X0 U104(.IN1(n188),.IN2(n3),.QN(n209));
  INVX0 U105(.INP(n167),.ZN(n159));
  INVX0 U106(.INP(n3),.ZN(n100));
  INVX0 U107(.INP(n166),.ZN(n157));
  INVX0 U108(.INP(n165),.ZN(n155));
  INVX0 U109(.INP(n164),.ZN(n153));
  INVX0 U110(.INP(n170),.ZN(n151));
  INVX0 U111(.INP(n107),.ZN(n104));
  INVX0 U112(.INP(n181),.ZN(n149));
  INVX0 U113(.INP(n191),.ZN(n146));
  NAND2X0 U114(.IN1(s_tem_prod[23:23]),.IN2(n96),.QN(n239));
  INVX0 U115(.INP(n201),.ZN(n142));
  INVX0 U116(.INP(n211),.ZN(n139));
  INVX0 U117(.INP(n221),.ZN(n135));
  NOR2X0 U118(.IN1(n239),.IN2(n5),.QN(n257));
  NOR2X0 U119(.IN1(n92),.IN2(n125),.QN(n286));
  NOR2X0 U120(.IN1(n103),.IN2(n4),.QN(n10));
  NOR2X0 U121(.IN1(n94),.IN2(n13),.QN(s_tem_prod[0:0]));
  NOR2X0 U122(.IN1(n94),.IN2(n24),.QN(s_tem_prod[1:1]));
  NOR2X0 U123(.IN1(n95),.IN2(n29),.QN(s_tem_prod[2:2]));
  NOR2X0 U124(.IN1(n104),.IN2(n291),.QN(N2461));
  NOR2X0 U125(.IN1(n104),.IN2(n292),.QN(N2462));
  NOR2X0 U126(.IN1(n104),.IN2(n242),.QN(N2463));
  NOR2X0 U127(.IN1(n104),.IN2(n246),.QN(N2464));
  NOR2X0 U128(.IN1(n104),.IN2(n250),.QN(N2465));
  NOR2X0 U129(.IN1(n104),.IN2(n254),.QN(N2466));
  NOR2X0 U130(.IN1(n104),.IN2(n259),.QN(N2467));
  NOR2X0 U131(.IN1(n104),.IN2(n261),.QN(N2468));
  INVX0 U132(.INP(n260),.ZN(n133));
  INVX0 U133(.INP(n255),.ZN(n128));
  INVX0 U134(.INP(n251),.ZN(n130));
  INVX0 U135(.INP(n247),.ZN(n126));
  INVX0 U136(.INP(n233),.ZN(n129));
  INVX0 U137(.INP(n238),.ZN(n127));
  INVX0 U138(.INP(n243),.ZN(n131));
  NOR2X0 U139(.IN1(n285),.IN2(n108),.QN(N2499));
  NOR2X0 U140(.IN1(n284),.IN2(n11),.QN(N2498));
  NOR2X0 U141(.IN1(n283),.IN2(n11),.QN(N2497));
  NOR2X0 U142(.IN1(n282),.IN2(n11),.QN(N2496));
  NOR2X0 U143(.IN1(n281),.IN2(n11),.QN(N2495));
  NOR2X0 U144(.IN1(n280),.IN2(n108),.QN(N2494));
  NOR2X0 U145(.IN1(n279),.IN2(n107),.QN(N2493));
  NOR2X0 U146(.IN1(n277),.IN2(n107),.QN(N2492));
  NOR2X0 U147(.IN1(n266),.IN2(n92),.QN(n267));
  INVX0 U148(.INP(n261),.ZN(n147));
  INVX0 U149(.INP(n277),.ZN(n124));
  NOR2X0 U150(.IN1(n92),.IN2(n275),.QN(n276));
  NOR2X0 U151(.IN1(n92),.IN2(n273),.QN(n274));
  NOR2X0 U152(.IN1(n92),.IN2(n271),.QN(n272));
  NOR2X0 U153(.IN1(n92),.IN2(n268),.QN(n270));
  NOR2X0 U154(.IN1(n264),.IN2(n92),.QN(n265));
  NOR2X0 U155(.IN1(n262),.IN2(n92),.QN(n263));
  INVX0 U156(.INP(\s_count[4] ),.ZN(n107));
  NOR2X0 U157(.IN1(n95),.IN2(n30),.QN(s_tem_prod[3:3]));
  NOR2X0 U158(.IN1(n95),.IN2(n31),.QN(s_tem_prod[4:4]));
  NOR2X0 U159(.IN1(n95),.IN2(n32),.QN(s_tem_prod[5:5]));
  NOR2X0 U160(.IN1(n95),.IN2(n33),.QN(s_tem_prod[6:6]));
  NOR2X0 U161(.IN1(n95),.IN2(n34),.QN(s_tem_prod[7:7]));
  NOR2X0 U162(.IN1(n95),.IN2(n35),.QN(s_tem_prod[8:8]));
  NOR2X0 U163(.IN1(n95),.IN2(n36),.QN(s_tem_prod[9:9]));
  INVX0 U164(.INP(\s_count[4] ),.ZN(n108));
  NOR2X0 U165(.IN1(n94),.IN2(n14),.QN(s_tem_prod[10:10]));
  NOR2X0 U166(.IN1(n94),.IN2(n15),.QN(s_tem_prod[11:11]));
  NOR2X0 U167(.IN1(n94),.IN2(n16),.QN(s_tem_prod[12:12]));
  NOR2X0 U168(.IN1(n94),.IN2(n17),.QN(s_tem_prod[13:13]));
  NOR2X0 U169(.IN1(n94),.IN2(n18),.QN(s_tem_prod[14:14]));
  NOR2X0 U170(.IN1(n94),.IN2(n19),.QN(s_tem_prod[15:15]));
  NOR2X0 U171(.IN1(n94),.IN2(n20),.QN(s_tem_prod[16:16]));
  NOR2X0 U172(.IN1(n94),.IN2(n21),.QN(s_tem_prod[17:17]));
  NOR2X0 U173(.IN1(n95),.IN2(n28),.QN(s_tem_prod[23:23]));
  NOR2X0 U174(.IN1(n94),.IN2(n22),.QN(s_tem_prod[18:18]));
  NOR2X0 U175(.IN1(n94),.IN2(n23),.QN(s_tem_prod[19:19]));
  NOR2X0 U176(.IN1(n95),.IN2(n26),.QN(s_tem_prod[21:21]));
  NOR2X0 U177(.IN1(n95),.IN2(n25),.QN(s_tem_prod[20:20]));
  NOR2X0 U178(.IN1(n95),.IN2(n27),.QN(s_tem_prod[22:22]));
  NAND2X1 U179(.IN1(n2),.IN2(n93),.QN(n6));
  INVX0 U180(.INP(s_state),.ZN(n113));
  INVX0 U181(.INP(s_state),.ZN(n114));
  INVX0 U182(.INP(s_state),.ZN(n115));
  INVX0 U183(.INP(n4),.ZN(n97));
  INVX0 U184(.INP(n3),.ZN(n101));
  INVX0 U185(.INP(n92),.ZN(n103));
  INVX0 U186(.INP(n107),.ZN(n106));
  INVX0 U187(.INP(n2),.ZN(n109));
  INVX0 U188(.INP(n2),.ZN(n110));
  INVX0 U189(.INP(n2),.ZN(n111));
  INVX0 U190(.INP(n2),.ZN(n112));
  XOR2X1 U191(.IN1(\add_118/carry[4] ),.IN2(n106),.Q(N1836));
  MUX41X1 U192(.IN1(s_fractb_i[18:18]),.IN3(s_fractb_i[19:19]),.IN2(s_fractb_i[22:22]),.IN4(s_fractb_i[23:23]),.S0(n97),.S1(n99),.Q(n116));
  MUX41X1 U193(.IN1(s_fractb_i[16:16]),.IN3(s_fractb_i[17:17]),.IN2(s_fractb_i[20:20]),.IN4(s_fractb_i[21:21]),.S0(n97),.S1(n99),.Q(n117));
  MUX21X1 U194(.IN1(n117),.IN2(n116),.S(n1),.Q(n118));
  MUX41X1 U195(.IN1(s_fractb_i[10:10]),.IN3(s_fractb_i[11:11]),.IN2(s_fractb_i[14:14]),.IN4(s_fractb_i[15:15]),.S0(n97),.S1(n99),.Q(n119));
  MUX41X1 U196(.IN1(s_fractb_i[8:8]),.IN3(s_fractb_i[9:9]),.IN2(s_fractb_i[12:12]),.IN4(s_fractb_i[13:13]),.S0(n97),.S1(n99),.Q(n120));
  MUX41X1 U197(.IN1(s_fractb_i[2:2]),.IN3(s_fractb_i[3:3]),.IN2(s_fractb_i[6:6]),.IN4(s_fractb_i[7:7]),.S0(n97),.S1(n99),.Q(n121));
  MUX41X1 U198(.IN1(s_fractb_i[0:0]),.IN3(s_fractb_i[1:1]),.IN2(s_fractb_i[4:4]),.IN4(s_fractb_i[5:5]),.S0(n97),.S1(n99),.Q(n122));
  MUX41X1 U199(.IN1(n122),.IN3(n120),.IN2(n121),.IN4(n119),.S0(n102),.S1(n98),.Q(n123));
  MUX21X1 U200(.IN1(n123),.IN2(n118),.S(n105),.Q(N2451));
  OR2X1 U202(.IN1(n169),.IN2(n1),.Q(n171));
  OR2X1 U203(.IN1(n171),.IN2(n101),.Q(n231));
  AND2X1 U204(.IN1(n108),.IN2(n196),.Q(N2453));
  MUX21X1 U205(.IN1(s_tem_prod[10:10]),.IN2(s_tem_prod[9:9]),.S(n97),.Q(n164));
  MUX21X1 U206(.IN1(s_tem_prod[8:8]),.IN2(s_tem_prod[7:7]),.S(n97),.Q(n165));
  MUX21X1 U207(.IN1(n153),.IN2(n155),.S(n1),.Q(n182));
  MUX21X1 U208(.IN1(s_tem_prod[6:6]),.IN2(s_tem_prod[5:5]),.S(n97),.Q(n166));
  MUX21X1 U209(.IN1(s_tem_prod[4:4]),.IN2(s_tem_prod[3:3]),.S(n97),.Q(n167));
  MUX21X1 U210(.IN1(n157),.IN2(n159),.S(n1),.Q(n184));
  MUX21X1 U211(.IN1(n182),.IN2(n184),.S(n100),.Q(n203));
  MUX21X1 U212(.IN1(s_tem_prod[2:2]),.IN2(s_tem_prod[1:1]),.S(n97),.Q(n168));
  MUX21X1 U213(.IN1(n160),.IN2(n169),.S(n1),.Q(n183));
  OR2X1 U214(.IN1(n183),.IN2(n101),.Q(n205));
  MUX21X1 U215(.IN1(n203),.IN2(n205),.S(n102),.Q(n242));
  MUX21X1 U216(.IN1(s_tem_prod[11:11]),.IN2(s_tem_prod[10:10]),.S(n97),.Q(n172));
  MUX21X1 U217(.IN1(s_tem_prod[9:9]),.IN2(s_tem_prod[8:8]),.S(n97),.Q(n175));
  MUX21X1 U218(.IN1(n172),.IN2(n175),.S(n1),.Q(n186));
  MUX21X1 U219(.IN1(s_tem_prod[7:7]),.IN2(s_tem_prod[6:6]),.S(n96),.Q(n174));
  MUX21X1 U220(.IN1(s_tem_prod[5:5]),.IN2(s_tem_prod[4:4]),.S(n96),.Q(n178));
  MUX21X1 U221(.IN1(n174),.IN2(n178),.S(n1),.Q(n189));
  MUX21X1 U222(.IN1(n186),.IN2(n189),.S(n100),.Q(n208));
  MUX21X1 U223(.IN1(s_tem_prod[3:3]),.IN2(s_tem_prod[2:2]),.S(n96),.Q(n177));
  MUX21X1 U224(.IN1(s_tem_prod[1:1]),.IN2(s_tem_prod[0:0]),.S(n96),.Q(n180));
  MUX21X1 U225(.IN1(n177),.IN2(n180),.S(n1),.Q(n188));
  MUX21X1 U226(.IN1(n152),.IN2(n209),.S(n102),.Q(n246));
  MUX21X1 U227(.IN1(s_tem_prod[12:12]),.IN2(s_tem_prod[11:11]),.S(n96),.Q(n170));
  MUX21X1 U228(.IN1(n151),.IN2(n153),.S(n1),.Q(n192));
  MUX21X1 U229(.IN1(n155),.IN2(n157),.S(n1),.Q(n194));
  MUX21X1 U230(.IN1(n192),.IN2(n194),.S(n100),.Q(n213));
  MUX21X1 U231(.IN1(n159),.IN2(n160),.S(n98),.Q(n193));
  MUX21X1 U232(.IN1(n193),.IN2(n171),.S(n100),.Q(n215));
  MUX21X1 U233(.IN1(n213),.IN2(n215),.S(n102),.Q(n250));
  MUX21X1 U234(.IN1(s_tem_prod[13:13]),.IN2(s_tem_prod[12:12]),.S(n96),.Q(n185));
  MUX21X1 U235(.IN1(n185),.IN2(n172),.S(n98),.Q(n173));
  MUX21X1 U236(.IN1(n175),.IN2(n174),.S(n98),.Q(n176));
  MUX21X1 U237(.IN1(n150),.IN2(n154),.S(n100),.Q(n218));
  MUX21X1 U238(.IN1(n178),.IN2(n177),.S(n98),.Q(n179));
  MUX21X1 U239(.IN1(n158),.IN2(n200),.S(n100),.Q(n220));
  MUX21X1 U240(.IN1(n218),.IN2(n220),.S(n102),.Q(n254));
  MUX21X1 U241(.IN1(s_tem_prod[14:14]),.IN2(s_tem_prod[13:13]),.S(n96),.Q(n181));
  MUX21X1 U242(.IN1(n149),.IN2(n151),.S(n98),.Q(n202));
  MUX21X1 U243(.IN1(n202),.IN2(n182),.S(n100),.Q(n223));
  MUX21X1 U244(.IN1(n184),.IN2(n183),.S(n100),.Q(n225));
  MUX21X1 U245(.IN1(n223),.IN2(n225),.S(n102),.Q(n259));
  MUX21X1 U246(.IN1(s_tem_prod[15:15]),.IN2(s_tem_prod[14:14]),.S(n96),.Q(n197));
  MUX21X1 U247(.IN1(n197),.IN2(n185),.S(n98),.Q(n207));
  MUX21X1 U248(.IN1(n207),.IN2(n186),.S(n100),.Q(n187));
  MUX21X1 U249(.IN1(n189),.IN2(n188),.S(n100),.Q(n190));
  MUX21X1 U250(.IN1(n148),.IN2(n156),.S(n102),.Q(n261));
  MUX21X1 U251(.IN1(s_tem_prod[16:16]),.IN2(s_tem_prod[15:15]),.S(n96),.Q(n191));
  MUX21X1 U252(.IN1(n146),.IN2(n149),.S(n98),.Q(n212));
  MUX21X1 U253(.IN1(n212),.IN2(n192),.S(n100),.Q(n230));
  MUX21X1 U254(.IN1(n194),.IN2(n193),.S(n100),.Q(n232));
  MUX21X1 U255(.IN1(n230),.IN2(n232),.S(n102),.Q(n195));
  MUX21X1 U256(.IN1(n145),.IN2(n196),.S(n105),.Q(N2469));
  MUX21X1 U257(.IN1(s_tem_prod[17:17]),.IN2(s_tem_prod[16:16]),.S(n96),.Q(n206));
  MUX21X1 U258(.IN1(n206),.IN2(n197),.S(n98),.Q(n198));
  MUX21X1 U259(.IN1(n144),.IN2(n150),.S(n100),.Q(n235));
  MUX21X1 U260(.IN1(n154),.IN2(n158),.S(n100),.Q(n237));
  MUX21X1 U261(.IN1(n235),.IN2(n237),.S(n102),.Q(n199));
  OR2X1 U262(.IN1(n200),.IN2(n101),.Q(n236));
  MUX21X1 U263(.IN1(n143),.IN2(n210),.S(n105),.Q(N2470));
  MUX21X1 U264(.IN1(s_tem_prod[18:18]),.IN2(s_tem_prod[17:17]),.S(n96),.Q(n201));
  MUX21X1 U265(.IN1(n142),.IN2(n146),.S(n98),.Q(n222));
  MUX21X1 U266(.IN1(n222),.IN2(n202),.S(n100),.Q(n241));
  MUX21X1 U267(.IN1(n241),.IN2(n203),.S(n102),.Q(n204));
  MUX21X1 U268(.IN1(n141),.IN2(n256),.S(n105),.Q(N2471));
  MUX21X1 U269(.IN1(s_tem_prod[19:19]),.IN2(s_tem_prod[18:18]),.S(n96),.Q(n216));
  MUX21X1 U270(.IN1(n216),.IN2(n206),.S(n98),.Q(n227));
  MUX21X1 U271(.IN1(n227),.IN2(n207),.S(n100),.Q(n245));
  MUX21X1 U272(.IN1(n208),.IN2(n245),.S(n92),.Q(n269));
  MUX21X1 U273(.IN1(n269),.IN2(n278),.S(n105),.Q(N2472));
  AND2X1 U274(.IN1(n108),.IN2(n210),.Q(N2454));
  MUX21X1 U275(.IN1(s_tem_prod[20:20]),.IN2(s_tem_prod[19:19]),.S(n96),.Q(n211));
  MUX21X1 U276(.IN1(n139),.IN2(n142),.S(n98),.Q(n229));
  MUX21X1 U277(.IN1(n229),.IN2(n212),.S(n99),.Q(n249));
  MUX21X1 U278(.IN1(n249),.IN2(n213),.S(n102),.Q(n214));
  MUX21X1 U279(.IN1(n138),.IN2(n287),.S(n105),.Q(N2473));
  MUX21X1 U280(.IN1(s_tem_prod[21:21]),.IN2(s_tem_prod[20:20]),.S(n96),.Q(n226));
  MUX21X1 U281(.IN1(n226),.IN2(n216),.S(n98),.Q(n217));
  MUX21X1 U282(.IN1(n137),.IN2(n144),.S(n100),.Q(n253));
  MUX21X1 U283(.IN1(n253),.IN2(n218),.S(n102),.Q(n219));
  MUX21X1 U284(.IN1(n136),.IN2(n288),.S(n105),.Q(N2474));
  MUX21X1 U285(.IN1(s_tem_prod[22:22]),.IN2(s_tem_prod[21:21]),.S(n96),.Q(n221));
  MUX21X1 U286(.IN1(n135),.IN2(n139),.S(n98),.Q(n240));
  MUX21X1 U287(.IN1(n240),.IN2(n222),.S(n99),.Q(n258));
  MUX21X1 U288(.IN1(n258),.IN2(n223),.S(n102),.Q(n224));
  MUX21X1 U289(.IN1(n134),.IN2(n289),.S(n105),.Q(N2475));
  MUX21X1 U290(.IN1(s_tem_prod[23:23]),.IN2(s_tem_prod[22:22]),.S(n96),.Q(n234));
  MUX21X1 U291(.IN1(n234),.IN2(n226),.S(n98),.Q(n244));
  MUX21X1 U292(.IN1(n244),.IN2(n227),.S(n99),.Q(n228));
  MUX21X1 U293(.IN1(n125),.IN2(n148),.S(n102),.Q(n277));
  MUX21X1 U294(.IN1(n124),.IN2(n290),.S(n105),.Q(N2476));
  MUX21X1 U295(.IN1(n239),.IN2(n135),.S(n98),.Q(n248));
  MUX21X1 U296(.IN1(n248),.IN2(n229),.S(n99),.Q(n262));
  MUX21X1 U297(.IN1(n262),.IN2(n230),.S(n102),.Q(n279));
  MUX21X1 U298(.IN1(n232),.IN2(n231),.S(n102),.Q(n291));
  MUX21X1 U299(.IN1(n279),.IN2(n291),.S(n105),.Q(n233));
  MUX21X1 U300(.IN1(n252),.IN2(n137),.S(n99),.Q(n264));
  MUX21X1 U301(.IN1(n264),.IN2(n235),.S(n102),.Q(n280));
  MUX21X1 U302(.IN1(n237),.IN2(n236),.S(n102),.Q(n292));
  MUX21X1 U303(.IN1(n280),.IN2(n292),.S(n105),.Q(n238));
  MUX21X1 U304(.IN1(n132),.IN2(n240),.S(n99),.Q(n266));
  MUX21X1 U305(.IN1(n266),.IN2(n241),.S(n103),.Q(n281));
  MUX21X1 U306(.IN1(n281),.IN2(n242),.S(n105),.Q(n243));
  MUX21X1 U307(.IN1(n268),.IN2(n140),.S(n103),.Q(n282));
  MUX21X1 U308(.IN1(n282),.IN2(n246),.S(n105),.Q(n247));
  OR2X1 U309(.IN1(n3),.IN2(n248),.Q(n271));
  MUX21X1 U310(.IN1(n271),.IN2(n249),.S(n103),.Q(n283));
  MUX21X1 U311(.IN1(n283),.IN2(n250),.S(n105),.Q(n251));
  OR2X1 U312(.IN1(n252),.IN2(n3),.Q(n273));
  MUX21X1 U313(.IN1(n273),.IN2(n253),.S(n103),.Q(n284));
  MUX21X1 U314(.IN1(n284),.IN2(n254),.S(n105),.Q(n255));
  AND2X1 U315(.IN1(n108),.IN2(n256),.Q(N2455));
  MUX21X1 U316(.IN1(n275),.IN2(n258),.S(n103),.Q(n285));
  MUX21X1 U317(.IN1(n285),.IN2(n259),.S(n105),.Q(n260));
  MUX21X1 U318(.IN1(n286),.IN2(n147),.S(n105),.Q(N2484));
  MUX21X1 U319(.IN1(n263),.IN2(n145),.S(n104),.Q(N2485));
  MUX21X1 U320(.IN1(n265),.IN2(n143),.S(n104),.Q(N2486));
  MUX21X1 U321(.IN1(n267),.IN2(n141),.S(n105),.Q(N2487));
  MUX21X1 U322(.IN1(n270),.IN2(n269),.S(n104),.Q(N2488));
  MUX21X1 U323(.IN1(n272),.IN2(n138),.S(n104),.Q(N2489));
  MUX21X1 U324(.IN1(n274),.IN2(n136),.S(n104),.Q(N2490));
  MUX21X1 U325(.IN1(n276),.IN2(n134),.S(n104),.Q(N2491));
  AND2X1 U326(.IN1(n11),.IN2(n278),.Q(N2456));
  AND2X1 U327(.IN1(n286),.IN2(n106),.Q(N2500));
  AND2X1 U328(.IN1(n11),.IN2(n287),.Q(N2457));
  AND2X1 U329(.IN1(n11),.IN2(n288),.Q(N2458));
  AND2X1 U330(.IN1(n11),.IN2(n289),.Q(N2459));
  AND2X1 U331(.IN1(n108),.IN2(n290),.Q(N2460));
endmodule
module post_norm_mul_DW01_inc_0_inj (A,SUM);
input [8:0] A ;
output [8:0] SUM ;
wire [8:2] carry ;
// instances
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[8:8]),.IN2(A[8:8]),.Q(SUM[8:8]));
endmodule
module post_norm_mul_DW01_inc_1_inj (A,SUM);
input [24:0] A ;
output [24:0] SUM ;
wire [24:2] carry ;
// instances
  HADDX1 U1_1_23(.A0(A[23:23]),.B0(carry[23:23]),.C1(carry[24:24]),.SO(SUM[23:23]));
  HADDX1 U1_1_22(.A0(A[22:22]),.B0(carry[22:22]),.C1(carry[23:23]),.SO(SUM[22:22]));
  HADDX1 U1_1_21(.A0(A[21:21]),.B0(carry[21:21]),.C1(carry[22:22]),.SO(SUM[21:21]));
  HADDX1 U1_1_20(.A0(A[20:20]),.B0(carry[20:20]),.C1(carry[21:21]),.SO(SUM[20:20]));
  HADDX1 U1_1_19(.A0(A[19:19]),.B0(carry[19:19]),.C1(carry[20:20]),.SO(SUM[19:19]));
  HADDX1 U1_1_18(.A0(A[18:18]),.B0(carry[18:18]),.C1(carry[19:19]),.SO(SUM[18:18]));
  HADDX1 U1_1_17(.A0(A[17:17]),.B0(carry[17:17]),.C1(carry[18:18]),.SO(SUM[17:17]));
  HADDX1 U1_1_16(.A0(A[16:16]),.B0(carry[16:16]),.C1(carry[17:17]),.SO(SUM[16:16]));
  HADDX1 U1_1_15(.A0(A[15:15]),.B0(carry[15:15]),.C1(carry[16:16]),.SO(SUM[15:15]));
  HADDX1 U1_1_14(.A0(A[14:14]),.B0(carry[14:14]),.C1(carry[15:15]),.SO(SUM[14:14]));
  HADDX1 U1_1_13(.A0(A[13:13]),.B0(carry[13:13]),.C1(carry[14:14]),.SO(SUM[13:13]));
  HADDX1 U1_1_12(.A0(A[12:12]),.B0(carry[12:12]),.C1(carry[13:13]),.SO(SUM[12:12]));
  HADDX1 U1_1_11(.A0(A[11:11]),.B0(carry[11:11]),.C1(carry[12:12]),.SO(SUM[11:11]));
  HADDX1 U1_1_10(.A0(A[10:10]),.B0(carry[10:10]),.C1(carry[11:11]),.SO(SUM[10:10]));
  HADDX1 U1_1_9(.A0(A[9:9]),.B0(carry[9:9]),.C1(carry[10:10]),.SO(SUM[9:9]));
  HADDX1 U1_1_8(.A0(A[8:8]),.B0(carry[8:8]),.C1(carry[9:9]),.SO(SUM[8:8]));
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[24:24]),.IN2(A[24:24]),.Q(SUM[24:24]));
endmodule
module post_norm_mul_DW01_sub_1_inj (A,B,CI,DIFF,CO);
input [5:0] A ;
input [5:0] B ;
output [5:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire [6:0] carry ;
// instances
  FADDX1 U2_4(.A(A[4:4]),.B(n2),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n3),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n4),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n5),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XNOR3X1 U1(.IN1(A[5:5]),.IN2(B[5:5]),.IN3(carry[5:5]),.Q(DIFF[5:5]));
  INVX0 U2(.INP(B[4:4]),.ZN(n2));
  INVX0 U3(.INP(B[2:2]),.ZN(n4));
  INVX0 U4(.INP(B[3:3]),.ZN(n3));
  INVX0 U5(.INP(B[1:1]),.ZN(n5));
  NAND2X1 U6(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U7(.INP(A[0:0]),.ZN(n1));
  XOR2X1 U8(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module post_norm_mul_DW01_sub_2_inj (A,B,CI,DIFF,CO);
input [9:0] A ;
input [9:0] B ;
output [9:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire [10:0] carry ;
// instances
  FADDX1 U2_5(.A(A[5:5]),.B(n9),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n10),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n11),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n12),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n13),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  INVX0 U1(.INP(A[7:7]),.ZN(n5));
  INVX0 U2(.INP(A[6:6]),.ZN(n3));
  INVX0 U3(.INP(carry[9:9]),.ZN(n7));
  INVX0 U4(.INP(carry[6:6]),.ZN(n4));
  AND2X1 U5(.IN1(n5),.IN2(n2),.Q(n1));
  AND2X1 U6(.IN1(n3),.IN2(n4),.Q(n2));
  NAND2X0 U7(.IN1(n6),.IN2(n1),.QN(carry[9:9]));
  INVX0 U8(.INP(A[8:8]),.ZN(n6));
  INVX0 U9(.INP(B[5:5]),.ZN(n9));
  INVX0 U10(.INP(B[3:3]),.ZN(n11));
  INVX0 U11(.INP(B[2:2]),.ZN(n12));
  INVX0 U12(.INP(B[1:1]),.ZN(n13));
  NAND2X0 U13(.IN1(n8),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U14(.INP(A[0:0]),.ZN(n8));
  INVX0 U15(.INP(B[4:4]),.ZN(n10));
  XOR2X1 U16(.IN1(n4),.IN2(A[6:6]),.Q(DIFF[6:6]));
  XOR2X1 U17(.IN1(n2),.IN2(A[7:7]),.Q(DIFF[7:7]));
  XOR2X1 U18(.IN1(n1),.IN2(A[8:8]),.Q(DIFF[8:8]));
  XOR2X1 U19(.IN1(n7),.IN2(A[9:9]),.Q(DIFF[9:9]));
  XOR2X1 U20(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module post_norm_mul_inj (clk_i,opa_i,opb_i,exp_10_i,fract_48_i,sign_i,rmode_i,output_o,ine_o);
input [31:0] opa_i ;
input [31:0] opb_i ;
input [9:0] exp_10_i ;
input [47:0] fract_48_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input clk_i ;
input sign_i ;
output ine_o ;
wire \s_rmode_i[1]  ;
wire N332 ;
wire N333 ;
wire N334 ;
wire N341 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N346 ;
wire N347 ;
wire N348 ;
wire N349 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N365 ;
wire N366 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N377 ;
wire N378 ;
wire N379 ;
wire N380 ;
wire N381 ;
wire N382 ;
wire N383 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N394 ;
wire N395 ;
wire N396 ;
wire N397 ;
wire N398 ;
wire N399 ;
wire N400 ;
wire N401 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N411 ;
wire N412 ;
wire N413 ;
wire N414 ;
wire N415 ;
wire N416 ;
wire N417 ;
wire N418 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N433 ;
wire N434 ;
wire N435 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N450 ;
wire N451 ;
wire N452 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N462 ;
wire N463 ;
wire N464 ;
wire N465 ;
wire N466 ;
wire N467 ;
wire N468 ;
wire N469 ;
wire N475 ;
wire N476 ;
wire N477 ;
wire N478 ;
wire N479 ;
wire N480 ;
wire N481 ;
wire N482 ;
wire N483 ;
wire N484 ;
wire N485 ;
wire N486 ;
wire N492 ;
wire N493 ;
wire N494 ;
wire N495 ;
wire N496 ;
wire N497 ;
wire N498 ;
wire N499 ;
wire N500 ;
wire N501 ;
wire N502 ;
wire N503 ;
wire N509 ;
wire N510 ;
wire N511 ;
wire N512 ;
wire N513 ;
wire N514 ;
wire N515 ;
wire N516 ;
wire N517 ;
wire N518 ;
wire N519 ;
wire N520 ;
wire N526 ;
wire N527 ;
wire N528 ;
wire N529 ;
wire N530 ;
wire N531 ;
wire N532 ;
wire N533 ;
wire N534 ;
wire N535 ;
wire N536 ;
wire N537 ;
wire N543 ;
wire N544 ;
wire N545 ;
wire N546 ;
wire N547 ;
wire N548 ;
wire N549 ;
wire N550 ;
wire N551 ;
wire N552 ;
wire N553 ;
wire N554 ;
wire N560 ;
wire N561 ;
wire N562 ;
wire N563 ;
wire N564 ;
wire N565 ;
wire N566 ;
wire N567 ;
wire N568 ;
wire N569 ;
wire N570 ;
wire N571 ;
wire N577 ;
wire N578 ;
wire N579 ;
wire N580 ;
wire N581 ;
wire N582 ;
wire N583 ;
wire N584 ;
wire N585 ;
wire N586 ;
wire N587 ;
wire N588 ;
wire N594 ;
wire N595 ;
wire N596 ;
wire N597 ;
wire N598 ;
wire N599 ;
wire N600 ;
wire N601 ;
wire N602 ;
wire N603 ;
wire N604 ;
wire N605 ;
wire N611 ;
wire N612 ;
wire N613 ;
wire N614 ;
wire N615 ;
wire N616 ;
wire N617 ;
wire N618 ;
wire N619 ;
wire N620 ;
wire N621 ;
wire N622 ;
wire N629 ;
wire N630 ;
wire N631 ;
wire N632 ;
wire N633 ;
wire N634 ;
wire N635 ;
wire N636 ;
wire N637 ;
wire N638 ;
wire N645 ;
wire N646 ;
wire N647 ;
wire N648 ;
wire N649 ;
wire N650 ;
wire N651 ;
wire N652 ;
wire N653 ;
wire N654 ;
wire N655 ;
wire N662 ;
wire N663 ;
wire N664 ;
wire N665 ;
wire N666 ;
wire N667 ;
wire N668 ;
wire N669 ;
wire N670 ;
wire N671 ;
wire N672 ;
wire N673 ;
wire N679 ;
wire N680 ;
wire N681 ;
wire N682 ;
wire N683 ;
wire N684 ;
wire N685 ;
wire N686 ;
wire N687 ;
wire N688 ;
wire N689 ;
wire N690 ;
wire N696 ;
wire N697 ;
wire N698 ;
wire N699 ;
wire N700 ;
wire N701 ;
wire N702 ;
wire N703 ;
wire N704 ;
wire N705 ;
wire N706 ;
wire N707 ;
wire N713 ;
wire N714 ;
wire N715 ;
wire N716 ;
wire N717 ;
wire N718 ;
wire N719 ;
wire N720 ;
wire N721 ;
wire N722 ;
wire N723 ;
wire N724 ;
wire N730 ;
wire N731 ;
wire N732 ;
wire N733 ;
wire N734 ;
wire N735 ;
wire N736 ;
wire N737 ;
wire N738 ;
wire N739 ;
wire N740 ;
wire N747 ;
wire N748 ;
wire N749 ;
wire N750 ;
wire N751 ;
wire N752 ;
wire N753 ;
wire N754 ;
wire N755 ;
wire N756 ;
wire N757 ;
wire N758 ;
wire N764 ;
wire N765 ;
wire N766 ;
wire N767 ;
wire N768 ;
wire N769 ;
wire N770 ;
wire N771 ;
wire N772 ;
wire N773 ;
wire N774 ;
wire N775 ;
wire N781 ;
wire N782 ;
wire N783 ;
wire N784 ;
wire N785 ;
wire N786 ;
wire N787 ;
wire N788 ;
wire N789 ;
wire N790 ;
wire N791 ;
wire N792 ;
wire N798 ;
wire N799 ;
wire N800 ;
wire N801 ;
wire N802 ;
wire N803 ;
wire N804 ;
wire N805 ;
wire N806 ;
wire N807 ;
wire N808 ;
wire N815 ;
wire N816 ;
wire N817 ;
wire N818 ;
wire N819 ;
wire N820 ;
wire N821 ;
wire N822 ;
wire N823 ;
wire N824 ;
wire N825 ;
wire N826 ;
wire N832 ;
wire N833 ;
wire N834 ;
wire N835 ;
wire N836 ;
wire N837 ;
wire N838 ;
wire N839 ;
wire N840 ;
wire N841 ;
wire N842 ;
wire N849 ;
wire N850 ;
wire N851 ;
wire N852 ;
wire N853 ;
wire N854 ;
wire N855 ;
wire N856 ;
wire N857 ;
wire N858 ;
wire N859 ;
wire N860 ;
wire N866 ;
wire N867 ;
wire N868 ;
wire N869 ;
wire N870 ;
wire N871 ;
wire N872 ;
wire N873 ;
wire N874 ;
wire N875 ;
wire N876 ;
wire N883 ;
wire N884 ;
wire N885 ;
wire N886 ;
wire N887 ;
wire N888 ;
wire N889 ;
wire N890 ;
wire N891 ;
wire N892 ;
wire N893 ;
wire N894 ;
wire N900 ;
wire N901 ;
wire N902 ;
wire N903 ;
wire N904 ;
wire N905 ;
wire N906 ;
wire N907 ;
wire N908 ;
wire N909 ;
wire N910 ;
wire N918 ;
wire N919 ;
wire N920 ;
wire N921 ;
wire N922 ;
wire N923 ;
wire N924 ;
wire N925 ;
wire N926 ;
wire N927 ;
wire N934 ;
wire N935 ;
wire N936 ;
wire N937 ;
wire N938 ;
wire N939 ;
wire N940 ;
wire N941 ;
wire N942 ;
wire N943 ;
wire N944 ;
wire N951 ;
wire N952 ;
wire N953 ;
wire N954 ;
wire N955 ;
wire N956 ;
wire N957 ;
wire N958 ;
wire N959 ;
wire N960 ;
wire N961 ;
wire N968 ;
wire N969 ;
wire N970 ;
wire N971 ;
wire N972 ;
wire N973 ;
wire N974 ;
wire N975 ;
wire N976 ;
wire N977 ;
wire N978 ;
wire N979 ;
wire N985 ;
wire N986 ;
wire N987 ;
wire N988 ;
wire N989 ;
wire N990 ;
wire N991 ;
wire N992 ;
wire N993 ;
wire N994 ;
wire N995 ;
wire N996 ;
wire N1002 ;
wire N1003 ;
wire N1004 ;
wire N1005 ;
wire N1006 ;
wire N1007 ;
wire N1008 ;
wire N1009 ;
wire N1010 ;
wire N1011 ;
wire N1012 ;
wire N1013 ;
wire N1019 ;
wire N1020 ;
wire N1021 ;
wire N1022 ;
wire N1023 ;
wire N1024 ;
wire N1025 ;
wire N1026 ;
wire N1027 ;
wire N1028 ;
wire N1029 ;
wire N1036 ;
wire N1037 ;
wire N1038 ;
wire N1039 ;
wire N1040 ;
wire N1041 ;
wire N1632 ;
wire N1633 ;
wire N1634 ;
wire N1635 ;
wire N1636 ;
wire N1637 ;
wire N1664 ;
wire N1665 ;
wire N1666 ;
wire N1672 ;
wire N1673 ;
wire N1674 ;
wire N1675 ;
wire N1677 ;
wire N1678 ;
wire N1679 ;
wire N1680 ;
wire N1686 ;
wire N1687 ;
wire N1688 ;
wire N1689 ;
wire N1690 ;
wire N1692 ;
wire N1693 ;
wire N1694 ;
wire N1695 ;
wire N1696 ;
wire N1702 ;
wire N1703 ;
wire N1704 ;
wire N1705 ;
wire N1706 ;
wire N1707 ;
wire N1708 ;
wire N1709 ;
wire N1710 ;
wire N1711 ;
wire N1712 ;
wire N1718 ;
wire N1719 ;
wire N1720 ;
wire N1721 ;
wire N1722 ;
wire N1723 ;
wire N1724 ;
wire N1725 ;
wire N1726 ;
wire N1727 ;
wire N1728 ;
wire N1729 ;
wire N1734 ;
wire N1735 ;
wire N1736 ;
wire N1737 ;
wire N1738 ;
wire N1739 ;
wire N1740 ;
wire N1741 ;
wire N1742 ;
wire N1743 ;
wire N1744 ;
wire N1745 ;
wire N1750 ;
wire N1751 ;
wire N1752 ;
wire N1753 ;
wire N1754 ;
wire N1755 ;
wire N1756 ;
wire N1757 ;
wire N1758 ;
wire N1759 ;
wire N1760 ;
wire N1761 ;
wire N1766 ;
wire N1767 ;
wire N1768 ;
wire N1769 ;
wire N1770 ;
wire N1771 ;
wire N1772 ;
wire N1773 ;
wire N1774 ;
wire N1775 ;
wire N1776 ;
wire N1777 ;
wire N1782 ;
wire N1783 ;
wire N1784 ;
wire N1785 ;
wire N1786 ;
wire N1787 ;
wire N1788 ;
wire N1789 ;
wire N1790 ;
wire N1791 ;
wire N1792 ;
wire N1793 ;
wire N1798 ;
wire N1799 ;
wire N1800 ;
wire N1801 ;
wire N1802 ;
wire N1804 ;
wire N1805 ;
wire N1806 ;
wire N1807 ;
wire N1808 ;
wire N1814 ;
wire N1815 ;
wire N1816 ;
wire N1817 ;
wire N1818 ;
wire N1819 ;
wire N1820 ;
wire N1821 ;
wire N1822 ;
wire N1823 ;
wire N1824 ;
wire N1825 ;
wire N1830 ;
wire N1831 ;
wire N1832 ;
wire N1833 ;
wire N1834 ;
wire N1835 ;
wire N1836 ;
wire N1837 ;
wire N1838 ;
wire N1839 ;
wire N1840 ;
wire N1841 ;
wire N1846 ;
wire N1847 ;
wire N1848 ;
wire N1849 ;
wire N1850 ;
wire N1851 ;
wire N1852 ;
wire N1853 ;
wire N1854 ;
wire N1855 ;
wire N1856 ;
wire N1857 ;
wire N1862 ;
wire N1863 ;
wire N1864 ;
wire N1865 ;
wire N1866 ;
wire N1867 ;
wire N1868 ;
wire N1869 ;
wire N1870 ;
wire N1871 ;
wire N1872 ;
wire N1873 ;
wire N1878 ;
wire N1879 ;
wire N1880 ;
wire N1881 ;
wire N1882 ;
wire N1883 ;
wire N1884 ;
wire N1885 ;
wire N1886 ;
wire N1887 ;
wire N1888 ;
wire N1889 ;
wire N1894 ;
wire N1895 ;
wire N1896 ;
wire N1897 ;
wire N1898 ;
wire N1899 ;
wire N1900 ;
wire N1901 ;
wire N1902 ;
wire N1903 ;
wire N1904 ;
wire N1910 ;
wire N1911 ;
wire N1912 ;
wire N1913 ;
wire N1914 ;
wire N1915 ;
wire N1916 ;
wire N1917 ;
wire N1918 ;
wire N1919 ;
wire N1920 ;
wire N1926 ;
wire N1927 ;
wire N1928 ;
wire N1929 ;
wire N1930 ;
wire N1931 ;
wire N1932 ;
wire N1933 ;
wire N1934 ;
wire N1935 ;
wire N1936 ;
wire N1937 ;
wire N1942 ;
wire N1943 ;
wire N1944 ;
wire N1945 ;
wire N1946 ;
wire N1947 ;
wire N1948 ;
wire N1949 ;
wire N1950 ;
wire N1951 ;
wire N1952 ;
wire N1953 ;
wire N1958 ;
wire N1959 ;
wire N1960 ;
wire N1961 ;
wire N1962 ;
wire N1963 ;
wire N1964 ;
wire N1965 ;
wire N1966 ;
wire N1967 ;
wire N1968 ;
wire N1969 ;
wire N1975 ;
wire N1976 ;
wire N1977 ;
wire N1978 ;
wire N1979 ;
wire N1980 ;
wire N1981 ;
wire N1982 ;
wire N1983 ;
wire N1984 ;
wire N1985 ;
wire N1990 ;
wire N1991 ;
wire N1992 ;
wire N1993 ;
wire N1994 ;
wire N1995 ;
wire N1996 ;
wire N1997 ;
wire N1998 ;
wire N1999 ;
wire N2000 ;
wire N2006 ;
wire N2007 ;
wire N2008 ;
wire N2009 ;
wire N2010 ;
wire N2011 ;
wire N2012 ;
wire N2013 ;
wire N2014 ;
wire N2015 ;
wire N2016 ;
wire N2022 ;
wire N2023 ;
wire N2024 ;
wire N2025 ;
wire N2026 ;
wire N2027 ;
wire N2028 ;
wire N2029 ;
wire N2030 ;
wire N2031 ;
wire N2032 ;
wire N2033 ;
wire N2038 ;
wire N2039 ;
wire N2040 ;
wire N2041 ;
wire N2042 ;
wire N2043 ;
wire N2044 ;
wire N2045 ;
wire N2046 ;
wire N2047 ;
wire N2048 ;
wire N2054 ;
wire N2055 ;
wire N2056 ;
wire N2057 ;
wire N2058 ;
wire N2059 ;
wire N2060 ;
wire N2061 ;
wire N2062 ;
wire N2063 ;
wire N2064 ;
wire N2070 ;
wire N2071 ;
wire N2072 ;
wire N2073 ;
wire N2074 ;
wire N2075 ;
wire N2076 ;
wire N2077 ;
wire N2078 ;
wire N2079 ;
wire N2080 ;
wire N2081 ;
wire N2086 ;
wire N2087 ;
wire N2088 ;
wire N2089 ;
wire N2090 ;
wire N2091 ;
wire N2092 ;
wire N2093 ;
wire N2094 ;
wire N2095 ;
wire N2096 ;
wire N2097 ;
wire N2102 ;
wire N2103 ;
wire N2104 ;
wire N2105 ;
wire N2106 ;
wire N2107 ;
wire N2108 ;
wire N2109 ;
wire N2110 ;
wire N2111 ;
wire N2112 ;
wire N2118 ;
wire N2119 ;
wire N2120 ;
wire N2121 ;
wire N2122 ;
wire N2123 ;
wire N2124 ;
wire N2125 ;
wire N2126 ;
wire N2127 ;
wire N2128 ;
wire N2129 ;
wire N2134 ;
wire N2135 ;
wire N2136 ;
wire N2137 ;
wire N2138 ;
wire N2139 ;
wire N2140 ;
wire N2141 ;
wire N2142 ;
wire N2143 ;
wire N2144 ;
wire N2145 ;
wire N2150 ;
wire N2151 ;
wire N2152 ;
wire N2153 ;
wire N2154 ;
wire N2155 ;
wire N2156 ;
wire N2157 ;
wire N2158 ;
wire N2159 ;
wire N2160 ;
wire N2166 ;
wire N2167 ;
wire N2168 ;
wire N2169 ;
wire N2170 ;
wire N2171 ;
wire N2172 ;
wire N2173 ;
wire N2174 ;
wire N2175 ;
wire N2176 ;
wire N2182 ;
wire N2183 ;
wire N2184 ;
wire N2185 ;
wire N2186 ;
wire N2187 ;
wire N2188 ;
wire N2189 ;
wire N2190 ;
wire N2191 ;
wire N2192 ;
wire N2193 ;
wire N2198 ;
wire N2199 ;
wire N2200 ;
wire N2201 ;
wire N2202 ;
wire N2203 ;
wire N2204 ;
wire N2205 ;
wire N2206 ;
wire N2207 ;
wire N2208 ;
wire N2214 ;
wire N2215 ;
wire N2216 ;
wire N2217 ;
wire N2218 ;
wire N2219 ;
wire N2220 ;
wire N2221 ;
wire N2222 ;
wire N2223 ;
wire N2224 ;
wire N2230 ;
wire N2231 ;
wire N2232 ;
wire N2233 ;
wire N2234 ;
wire N2235 ;
wire N2236 ;
wire N2237 ;
wire N2238 ;
wire N2239 ;
wire N2240 ;
wire N2246 ;
wire N2247 ;
wire N2248 ;
wire N2249 ;
wire N2250 ;
wire N2251 ;
wire N2252 ;
wire N2253 ;
wire N2254 ;
wire N2255 ;
wire N2256 ;
wire N2262 ;
wire N2263 ;
wire N2264 ;
wire N2265 ;
wire N2266 ;
wire N2267 ;
wire N2268 ;
wire N2269 ;
wire N2270 ;
wire N2271 ;
wire N2272 ;
wire N2278 ;
wire N2279 ;
wire N2280 ;
wire N2281 ;
wire N2282 ;
wire N2284 ;
wire N2285 ;
wire N2286 ;
wire N2287 ;
wire N2288 ;
wire N2289 ;
wire N2294 ;
wire N2295 ;
wire N2296 ;
wire N2297 ;
wire N2298 ;
wire N2299 ;
wire N2300 ;
wire N2301 ;
wire N2302 ;
wire N2303 ;
wire N2304 ;
wire N2310 ;
wire N2311 ;
wire N2312 ;
wire N2313 ;
wire N2314 ;
wire N2315 ;
wire N2316 ;
wire N2317 ;
wire N2318 ;
wire N2319 ;
wire N2320 ;
wire N2326 ;
wire N2327 ;
wire N2328 ;
wire N2329 ;
wire N2330 ;
wire N2331 ;
wire N2332 ;
wire N2333 ;
wire N2334 ;
wire N2335 ;
wire N2336 ;
wire N2337 ;
wire N2343 ;
wire N2344 ;
wire N2345 ;
wire N2346 ;
wire N2347 ;
wire N2348 ;
wire N2349 ;
wire N2350 ;
wire N2351 ;
wire N2352 ;
wire N2358 ;
wire N2359 ;
wire N2360 ;
wire N2361 ;
wire N2362 ;
wire N2363 ;
wire N2974 ;
wire N2975 ;
wire N2976 ;
wire N2977 ;
wire N2978 ;
wire N2979 ;
wire N2999 ;
wire N3000 ;
wire N3001 ;
wire N3002 ;
wire N3003 ;
wire N3004 ;
wire N3005 ;
wire N3019 ;
wire N3020 ;
wire N3021 ;
wire N3022 ;
wire N3023 ;
wire N3024 ;
wire N3065 ;
wire N3066 ;
wire N3067 ;
wire N3068 ;
wire N3069 ;
wire N3070 ;
wire N3072 ;
wire N3073 ;
wire N3074 ;
wire N3075 ;
wire N3076 ;
wire N3077 ;
wire N3078 ;
wire N3081 ;
wire N3082 ;
wire N3083 ;
wire N3084 ;
wire N3085 ;
wire N3086 ;
wire N3093 ;
wire N3094 ;
wire N3095 ;
wire N3096 ;
wire N3097 ;
wire N3098 ;
wire N3099 ;
wire N3100 ;
wire N3101 ;
wire N3102 ;
wire N3103 ;
wire N3104 ;
wire N3105 ;
wire N3106 ;
wire N3107 ;
wire N3108 ;
wire N3109 ;
wire N3110 ;
wire N3111 ;
wire N3112 ;
wire N3113 ;
wire N3114 ;
wire N3115 ;
wire N3116 ;
wire N3117 ;
wire N3118 ;
wire N3119 ;
wire N3120 ;
wire N3121 ;
wire N3122 ;
wire N3123 ;
wire N3124 ;
wire N3125 ;
wire N3126 ;
wire N3127 ;
wire N3128 ;
wire N3129 ;
wire N3130 ;
wire N3131 ;
wire N3132 ;
wire N3133 ;
wire N3134 ;
wire N3135 ;
wire N3136 ;
wire N3137 ;
wire N3138 ;
wire N3139 ;
wire N3140 ;
wire N3141 ;
wire N3142 ;
wire N3143 ;
wire N3144 ;
wire N3145 ;
wire N3146 ;
wire N3147 ;
wire N3148 ;
wire N3149 ;
wire N3150 ;
wire N3151 ;
wire N3152 ;
wire N3153 ;
wire N3154 ;
wire N3155 ;
wire N3156 ;
wire N3157 ;
wire N3158 ;
wire N3159 ;
wire N3160 ;
wire N3161 ;
wire N3162 ;
wire N3163 ;
wire N3164 ;
wire N3165 ;
wire N3166 ;
wire N3167 ;
wire N3168 ;
wire N3169 ;
wire N3170 ;
wire N3171 ;
wire N3172 ;
wire N3185 ;
wire N3186 ;
wire N3187 ;
wire N3188 ;
wire N3189 ;
wire N3190 ;
wire N3191 ;
wire N3192 ;
wire N3193 ;
wire N3194 ;
wire N3195 ;
wire N3196 ;
wire N3197 ;
wire N3198 ;
wire N3199 ;
wire N3200 ;
wire N3201 ;
wire N3202 ;
wire N3203 ;
wire N3204 ;
wire N3205 ;
wire N3206 ;
wire N3207 ;
wire N3208 ;
wire N3209 ;
wire N3210 ;
wire N3211 ;
wire N3212 ;
wire N3213 ;
wire N3214 ;
wire N3215 ;
wire N3216 ;
wire N3217 ;
wire N3218 ;
wire N3219 ;
wire N3220 ;
wire N3221 ;
wire N3222 ;
wire N3223 ;
wire N3224 ;
wire N3225 ;
wire N3226 ;
wire N3227 ;
wire N3228 ;
wire N3229 ;
wire N3230 ;
wire N3231 ;
wire N3232 ;
wire N3233 ;
wire N3234 ;
wire N3235 ;
wire N3236 ;
wire N3238 ;
wire N3239 ;
wire N3240 ;
wire N3241 ;
wire N3242 ;
wire N3243 ;
wire N3244 ;
wire N3278 ;
wire N3279 ;
wire N3280 ;
wire N3281 ;
wire N3282 ;
wire N3283 ;
wire N3284 ;
wire N3285 ;
wire N3286 ;
wire N3287 ;
wire N3288 ;
wire N3289 ;
wire N3290 ;
wire N3291 ;
wire N3292 ;
wire N3293 ;
wire N3294 ;
wire N3295 ;
wire N3296 ;
wire N3297 ;
wire N3298 ;
wire N3299 ;
wire N3300 ;
wire N3301 ;
wire N3302 ;
wire N3303 ;
wire N3304 ;
wire N3305 ;
wire N3306 ;
wire N3307 ;
wire N3308 ;
wire N3309 ;
wire N3310 ;
wire N3311 ;
wire N3312 ;
wire N3313 ;
wire N3314 ;
wire N3315 ;
wire N3316 ;
wire N3317 ;
wire N3318 ;
wire N3319 ;
wire N3320 ;
wire N3321 ;
wire N3322 ;
wire N3323 ;
wire N3324 ;
wire N3325 ;
wire N3326 ;
wire N3327 ;
wire N3346 ;
wire N3347 ;
wire N3348 ;
wire N3349 ;
wire N3350 ;
wire N3351 ;
wire N3352 ;
wire N3353 ;
wire N3354 ;
wire N3532 ;
wire n68 ;
wire n69 ;
wire n118 ;
wire n119 ;
wire n122 ;
wire n123 ;
wire n130 ;
wire n137 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n152 ;
wire n154 ;
wire n156 ;
wire n158 ;
wire n160 ;
wire n162 ;
wire n164 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n177 ;
wire n182 ;
wire n189 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n204 ;
wire n206 ;
wire n208 ;
wire n210 ;
wire n212 ;
wire n214 ;
wire n215 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n229 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n235 ;
wire n236 ;
wire n238 ;
wire n244 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n351 ;
wire n352 ;
wire n354 ;
wire n355 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n406 ;
wire n407 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire n429 ;
wire n430 ;
wire n431 ;
wire n434 ;
wire n435 ;
wire n436 ;
wire n437 ;
wire n438 ;
wire n439 ;
wire n440 ;
wire n441 ;
wire n442 ;
wire n443 ;
wire n444 ;
wire n447 ;
wire n448 ;
wire n449 ;
wire n450 ;
wire n452 ;
wire n453 ;
wire n454 ;
wire n455 ;
wire n456 ;
wire n457 ;
wire n460 ;
wire n461 ;
wire n462 ;
wire n463 ;
wire n464 ;
wire n465 ;
wire n466 ;
wire n467 ;
wire n468 ;
wire n469 ;
wire n472 ;
wire n473 ;
wire n474 ;
wire n475 ;
wire n476 ;
wire n477 ;
wire n480 ;
wire n481 ;
wire n482 ;
wire n483 ;
wire n484 ;
wire n485 ;
wire n489 ;
wire n490 ;
wire n491 ;
wire n492 ;
wire n493 ;
wire n494 ;
wire n495 ;
wire n496 ;
wire n497 ;
wire n498 ;
wire n501 ;
wire n502 ;
wire n503 ;
wire n504 ;
wire n505 ;
wire n506 ;
wire n509 ;
wire n510 ;
wire n511 ;
wire n512 ;
wire n513 ;
wire n514 ;
wire n515 ;
wire n518 ;
wire n519 ;
wire n520 ;
wire n521 ;
wire n522 ;
wire n523 ;
wire n524 ;
wire n525 ;
wire n526 ;
wire n527 ;
wire n528 ;
wire n529 ;
wire n530 ;
wire n531 ;
wire n532 ;
wire n533 ;
wire n534 ;
wire n535 ;
wire n536 ;
wire n537 ;
wire n538 ;
wire n539 ;
wire n540 ;
wire n541 ;
wire n542 ;
wire n543 ;
wire n544 ;
wire n545 ;
wire n546 ;
wire n547 ;
wire n548 ;
wire n549 ;
wire n550 ;
wire n551 ;
wire n552 ;
wire n553 ;
wire n554 ;
wire n555 ;
wire n556 ;
wire n557 ;
wire n558 ;
wire n559 ;
wire n560 ;
wire n561 ;
wire n562 ;
wire n563 ;
wire n564 ;
wire n565 ;
wire n566 ;
wire n567 ;
wire n568 ;
wire n569 ;
wire n570 ;
wire n571 ;
wire n573 ;
wire n574 ;
wire n575 ;
wire n577 ;
wire n578 ;
wire n579 ;
wire n580 ;
wire n581 ;
wire n582 ;
wire n583 ;
wire n584 ;
wire n585 ;
wire n586 ;
wire n587 ;
wire n588 ;
wire n589 ;
wire n590 ;
wire n592 ;
wire n593 ;
wire n595 ;
wire n598 ;
wire n599 ;
wire n600 ;
wire n601 ;
wire n602 ;
wire n603 ;
wire n604 ;
wire n605 ;
wire n606 ;
wire n607 ;
wire n608 ;
wire n609 ;
wire n610 ;
wire n611 ;
wire n612 ;
wire n615 ;
wire n616 ;
wire n617 ;
wire n618 ;
wire n619 ;
wire n622 ;
wire n623 ;
wire n624 ;
wire n625 ;
wire n626 ;
wire n627 ;
wire n628 ;
wire n629 ;
wire n630 ;
wire n631 ;
wire n632 ;
wire n635 ;
wire n636 ;
wire n637 ;
wire n638 ;
wire n639 ;
wire n640 ;
wire n643 ;
wire n644 ;
wire n647 ;
wire n648 ;
wire n649 ;
wire n650 ;
wire n651 ;
wire n652 ;
wire n653 ;
wire n654 ;
wire n655 ;
wire n656 ;
wire n659 ;
wire n660 ;
wire n661 ;
wire n662 ;
wire n663 ;
wire n664 ;
wire n665 ;
wire n666 ;
wire n667 ;
wire n668 ;
wire n669 ;
wire n670 ;
wire n673 ;
wire n674 ;
wire n675 ;
wire n676 ;
wire n677 ;
wire n678 ;
wire n679 ;
wire n680 ;
wire n681 ;
wire n682 ;
wire n685 ;
wire n686 ;
wire n687 ;
wire n690 ;
wire n691 ;
wire n692 ;
wire n693 ;
wire n694 ;
wire n695 ;
wire n696 ;
wire n697 ;
wire n698 ;
wire n701 ;
wire n702 ;
wire n703 ;
wire n704 ;
wire n705 ;
wire n706 ;
wire n707 ;
wire n708 ;
wire n709 ;
wire n710 ;
wire n711 ;
wire n714 ;
wire n715 ;
wire n716 ;
wire n717 ;
wire n718 ;
wire n719 ;
wire n720 ;
wire n721 ;
wire n724 ;
wire n725 ;
wire n726 ;
wire n727 ;
wire n728 ;
wire n729 ;
wire n730 ;
wire n731 ;
wire n732 ;
wire n733 ;
wire n736 ;
wire n737 ;
wire n738 ;
wire n739 ;
wire n740 ;
wire n741 ;
wire n744 ;
wire n745 ;
wire n746 ;
wire n747 ;
wire n748 ;
wire n749 ;
wire n750 ;
wire n751 ;
wire n752 ;
wire n753 ;
wire n754 ;
wire n755 ;
wire n756 ;
wire n757 ;
wire n758 ;
wire n759 ;
wire n760 ;
wire n761 ;
wire n762 ;
wire n763 ;
wire n764 ;
wire n765 ;
wire n766 ;
wire n767 ;
wire n768 ;
wire n769 ;
wire n770 ;
wire n771 ;
wire n772 ;
wire n773 ;
wire n774 ;
wire n775 ;
wire n776 ;
wire n777 ;
wire n778 ;
wire n779 ;
wire n780 ;
wire n781 ;
wire n782 ;
wire n783 ;
wire n784 ;
wire n785 ;
wire n786 ;
wire n787 ;
wire n788 ;
wire n789 ;
wire n790 ;
wire n791 ;
wire n792 ;
wire n793 ;
wire n794 ;
wire n795 ;
wire n796 ;
wire n797 ;
wire n798 ;
wire n799 ;
wire n800 ;
wire n801 ;
wire n802 ;
wire n803 ;
wire N2993 ;
wire \add_197/carry[4]  ;
wire \add_197/carry[3]  ;
wire \add_197/carry[2]  ;
wire \add_197/carry[1]  ;
wire \sub_192_aco/carry[7]  ;
wire \sub_192_aco/carry[6]  ;
wire \sub_192_aco/carry[5]  ;
wire \sub_192_aco/carry[4]  ;
wire \sub_192_aco/carry[3]  ;
wire \sub_192_aco/carry[2]  ;
wire \sub_192_aco/carry[1]  ;
wire \add_140/carry[8]  ;
wire \add_140/carry[7]  ;
wire \add_140/carry[6]  ;
wire \add_140/carry[5]  ;
wire \add_140/carry[4]  ;
wire \add_140/carry[3]  ;
wire \add_140/carry[2]  ;
wire \add_140/carry[1]  ;
wire \add_105_I48_L14036_C136/carry[5]  ;
wire \add_105_I48_L14036_C136/carry[4]  ;
wire \add_105_I48_L14036_C136/carry[3]  ;
wire \add_105_I48_L14036_C136/carry[2]  ;
wire \add_105_I47_L14036_C136/carry[5]  ;
wire \add_105_I47_L14036_C136/carry[4]  ;
wire \add_105_I47_L14036_C136/carry[3]  ;
wire \add_105_I47_L14036_C136/carry[2]  ;
wire \add_105_I46_L14036_C136/carry[5]  ;
wire \add_105_I46_L14036_C136/carry[4]  ;
wire \add_105_I46_L14036_C136/carry[3]  ;
wire \add_105_I46_L14036_C136/carry[2]  ;
wire \add_105_I45_L14036_C136/carry[5]  ;
wire \add_105_I45_L14036_C136/carry[4]  ;
wire \add_105_I45_L14036_C136/carry[3]  ;
wire \add_105_I45_L14036_C136/carry[2]  ;
wire \add_105_I44_L14036_C136/carry[5]  ;
wire \add_105_I44_L14036_C136/carry[4]  ;
wire \add_105_I44_L14036_C136/carry[3]  ;
wire \add_105_I44_L14036_C136/carry[2]  ;
wire \add_105_I43_L14036_C136/carry[5]  ;
wire \add_105_I43_L14036_C136/carry[4]  ;
wire \add_105_I43_L14036_C136/carry[3]  ;
wire \add_105_I43_L14036_C136/carry[2]  ;
wire \add_105_I42_L14036_C136/carry[5]  ;
wire \add_105_I42_L14036_C136/carry[4]  ;
wire \add_105_I42_L14036_C136/carry[3]  ;
wire \add_105_I42_L14036_C136/carry[2]  ;
wire \add_105_I41_L14036_C136/carry[5]  ;
wire \add_105_I41_L14036_C136/carry[4]  ;
wire \add_105_I41_L14036_C136/carry[3]  ;
wire \add_105_I41_L14036_C136/carry[2]  ;
wire \add_105_I40_L14036_C136/carry[5]  ;
wire \add_105_I40_L14036_C136/carry[4]  ;
wire \add_105_I40_L14036_C136/carry[3]  ;
wire \add_105_I40_L14036_C136/carry[2]  ;
wire \add_105_I39_L14036_C136/carry[5]  ;
wire \add_105_I39_L14036_C136/carry[4]  ;
wire \add_105_I39_L14036_C136/carry[3]  ;
wire \add_105_I39_L14036_C136/carry[2]  ;
wire \add_105_I38_L14036_C136/carry[5]  ;
wire \add_105_I38_L14036_C136/carry[4]  ;
wire \add_105_I38_L14036_C136/carry[3]  ;
wire \add_105_I38_L14036_C136/carry[2]  ;
wire \add_105_I37_L14036_C136/carry[5]  ;
wire \add_105_I37_L14036_C136/carry[4]  ;
wire \add_105_I37_L14036_C136/carry[3]  ;
wire \add_105_I37_L14036_C136/carry[2]  ;
wire \add_105_I36_L14036_C136/carry[5]  ;
wire \add_105_I36_L14036_C136/carry[4]  ;
wire \add_105_I36_L14036_C136/carry[3]  ;
wire \add_105_I36_L14036_C136/carry[2]  ;
wire \add_105_I35_L14036_C136/carry[5]  ;
wire \add_105_I35_L14036_C136/carry[4]  ;
wire \add_105_I35_L14036_C136/carry[3]  ;
wire \add_105_I35_L14036_C136/carry[2]  ;
wire \add_105_I34_L14036_C136/carry[5]  ;
wire \add_105_I34_L14036_C136/carry[4]  ;
wire \add_105_I34_L14036_C136/carry[3]  ;
wire \add_105_I34_L14036_C136/carry[2]  ;
wire \add_105_I33_L14036_C136/carry[5]  ;
wire \add_105_I33_L14036_C136/carry[4]  ;
wire \add_105_I33_L14036_C136/carry[3]  ;
wire \add_105_I33_L14036_C136/carry[2]  ;
wire \add_105_I32_L14036_C136/carry[5]  ;
wire \add_105_I32_L14036_C136/carry[4]  ;
wire \add_105_I32_L14036_C136/carry[3]  ;
wire \add_105_I32_L14036_C136/carry[2]  ;
wire \add_105_I31_L14036_C136/carry[5]  ;
wire \add_105_I31_L14036_C136/carry[4]  ;
wire \add_105_I31_L14036_C136/carry[3]  ;
wire \add_105_I31_L14036_C136/carry[2]  ;
wire \add_105_I30_L14036_C136/carry[5]  ;
wire \add_105_I30_L14036_C136/carry[4]  ;
wire \add_105_I30_L14036_C136/carry[3]  ;
wire \add_105_I30_L14036_C136/carry[2]  ;
wire \add_105_I29_L14036_C136/carry[5]  ;
wire \add_105_I29_L14036_C136/carry[4]  ;
wire \add_105_I29_L14036_C136/carry[3]  ;
wire \add_105_I29_L14036_C136/carry[2]  ;
wire \add_105_I28_L14036_C136/carry[5]  ;
wire \add_105_I28_L14036_C136/carry[4]  ;
wire \add_105_I28_L14036_C136/carry[3]  ;
wire \add_105_I28_L14036_C136/carry[2]  ;
wire \add_105_I27_L14036_C136/carry[5]  ;
wire \add_105_I27_L14036_C136/carry[4]  ;
wire \add_105_I27_L14036_C136/carry[3]  ;
wire \add_105_I27_L14036_C136/carry[2]  ;
wire \add_105_I26_L14036_C136/carry[5]  ;
wire \add_105_I26_L14036_C136/carry[4]  ;
wire \add_105_I26_L14036_C136/carry[3]  ;
wire \add_105_I26_L14036_C136/carry[2]  ;
wire \add_105_I25_L14036_C136/carry[5]  ;
wire \add_105_I25_L14036_C136/carry[4]  ;
wire \add_105_I25_L14036_C136/carry[3]  ;
wire \add_105_I25_L14036_C136/carry[2]  ;
wire \add_105_I24_L14036_C136/carry[5]  ;
wire \add_105_I24_L14036_C136/carry[4]  ;
wire \add_105_I24_L14036_C136/carry[3]  ;
wire \add_105_I24_L14036_C136/carry[2]  ;
wire \add_105_I23_L14036_C136/carry[5]  ;
wire \add_105_I23_L14036_C136/carry[4]  ;
wire \add_105_I23_L14036_C136/carry[3]  ;
wire \add_105_I23_L14036_C136/carry[2]  ;
wire \add_105_I22_L14036_C136/carry[5]  ;
wire \add_105_I22_L14036_C136/carry[4]  ;
wire \add_105_I22_L14036_C136/carry[3]  ;
wire \add_105_I22_L14036_C136/carry[2]  ;
wire \add_105_I21_L14036_C136/carry[5]  ;
wire \add_105_I21_L14036_C136/carry[4]  ;
wire \add_105_I21_L14036_C136/carry[3]  ;
wire \add_105_I21_L14036_C136/carry[2]  ;
wire \add_105_I20_L14036_C136/carry[5]  ;
wire \add_105_I20_L14036_C136/carry[4]  ;
wire \add_105_I20_L14036_C136/carry[3]  ;
wire \add_105_I20_L14036_C136/carry[2]  ;
wire \add_105_I19_L14036_C136/carry[5]  ;
wire \add_105_I19_L14036_C136/carry[4]  ;
wire \add_105_I19_L14036_C136/carry[3]  ;
wire \add_105_I19_L14036_C136/carry[2]  ;
wire \add_105_I18_L14036_C136/carry[5]  ;
wire \add_105_I18_L14036_C136/carry[4]  ;
wire \add_105_I18_L14036_C136/carry[3]  ;
wire \add_105_I18_L14036_C136/carry[2]  ;
wire \add_105_I17_L14036_C136/carry[5]  ;
wire \add_105_I17_L14036_C136/carry[4]  ;
wire \add_105_I17_L14036_C136/carry[3]  ;
wire \add_105_I17_L14036_C136/carry[2]  ;
wire \add_105_I16_L14036_C136/carry[5]  ;
wire \add_105_I16_L14036_C136/carry[4]  ;
wire \add_105_I16_L14036_C136/carry[3]  ;
wire \add_105_I16_L14036_C136/carry[2]  ;
wire \add_105_I15_L14036_C136/carry[5]  ;
wire \add_105_I15_L14036_C136/carry[4]  ;
wire \add_105_I15_L14036_C136/carry[3]  ;
wire \add_105_I15_L14036_C136/carry[2]  ;
wire \add_105_I14_L14036_C136/carry[5]  ;
wire \add_105_I14_L14036_C136/carry[4]  ;
wire \add_105_I14_L14036_C136/carry[3]  ;
wire \add_105_I14_L14036_C136/carry[2]  ;
wire \add_105_I13_L14036_C136/carry[5]  ;
wire \add_105_I13_L14036_C136/carry[4]  ;
wire \add_105_I13_L14036_C136/carry[3]  ;
wire \add_105_I13_L14036_C136/carry[2]  ;
wire \add_105_I12_L14036_C136/carry[5]  ;
wire \add_105_I12_L14036_C136/carry[4]  ;
wire \add_105_I12_L14036_C136/carry[3]  ;
wire \add_105_I12_L14036_C136/carry[2]  ;
wire \add_105_I11_L14036_C136/carry[5]  ;
wire \add_105_I11_L14036_C136/carry[4]  ;
wire \add_105_I11_L14036_C136/carry[3]  ;
wire \add_105_I11_L14036_C136/carry[2]  ;
wire \add_105_I10_L14036_C136/carry[5]  ;
wire \add_105_I10_L14036_C136/carry[4]  ;
wire \add_105_I10_L14036_C136/carry[3]  ;
wire \add_105_I10_L14036_C136/carry[2]  ;
wire \add_105_I9_L14036_C136/carry[5]  ;
wire \add_105_I9_L14036_C136/carry[4]  ;
wire \add_105_I9_L14036_C136/carry[3]  ;
wire \add_105_I9_L14036_C136/carry[2]  ;
wire \add_105_I8_L14036_C136/carry[5]  ;
wire \add_105_I8_L14036_C136/carry[4]  ;
wire \add_105_I8_L14036_C136/carry[3]  ;
wire \add_105_I8_L14036_C136/carry[2]  ;
wire \add_105_I7_L14036_C136/carry[4]  ;
wire \add_105_I7_L14036_C136/carry[3]  ;
wire \add_105_I7_L14036_C136/carry[2]  ;
wire \add_105_I6_L14036_C136/carry[2]  ;
wire \add_105_I6_L14036_C136/carry[3]  ;
wire \add_105_I5_L14036_C136/carry[2]  ;
wire \add_90_I46_L14036_C132/carry[5]  ;
wire \add_90_I46_L14036_C132/carry[4]  ;
wire \add_90_I46_L14036_C132/carry[3]  ;
wire \add_90_I46_L14036_C132/carry[2]  ;
wire \add_90_I45_L14036_C132/carry[5]  ;
wire \add_90_I45_L14036_C132/carry[4]  ;
wire \add_90_I45_L14036_C132/carry[3]  ;
wire \add_90_I45_L14036_C132/carry[2]  ;
wire \add_90_I44_L14036_C132/carry[5]  ;
wire \add_90_I44_L14036_C132/carry[4]  ;
wire \add_90_I44_L14036_C132/carry[3]  ;
wire \add_90_I44_L14036_C132/carry[2]  ;
wire \add_90_I43_L14036_C132/carry[5]  ;
wire \add_90_I43_L14036_C132/carry[4]  ;
wire \add_90_I43_L14036_C132/carry[3]  ;
wire \add_90_I43_L14036_C132/carry[2]  ;
wire \add_90_I42_L14036_C132/carry[5]  ;
wire \add_90_I42_L14036_C132/carry[4]  ;
wire \add_90_I42_L14036_C132/carry[3]  ;
wire \add_90_I42_L14036_C132/carry[2]  ;
wire \add_90_I41_L14036_C132/carry[5]  ;
wire \add_90_I41_L14036_C132/carry[4]  ;
wire \add_90_I41_L14036_C132/carry[3]  ;
wire \add_90_I41_L14036_C132/carry[2]  ;
wire \add_90_I40_L14036_C132/carry[5]  ;
wire \add_90_I40_L14036_C132/carry[4]  ;
wire \add_90_I40_L14036_C132/carry[3]  ;
wire \add_90_I40_L14036_C132/carry[2]  ;
wire \add_90_I39_L14036_C132/carry[5]  ;
wire \add_90_I39_L14036_C132/carry[4]  ;
wire \add_90_I39_L14036_C132/carry[3]  ;
wire \add_90_I39_L14036_C132/carry[2]  ;
wire \add_90_I38_L14036_C132/carry[5]  ;
wire \add_90_I38_L14036_C132/carry[4]  ;
wire \add_90_I38_L14036_C132/carry[3]  ;
wire \add_90_I38_L14036_C132/carry[2]  ;
wire \add_90_I37_L14036_C132/carry[5]  ;
wire \add_90_I37_L14036_C132/carry[4]  ;
wire \add_90_I37_L14036_C132/carry[3]  ;
wire \add_90_I37_L14036_C132/carry[2]  ;
wire \add_90_I36_L14036_C132/carry[5]  ;
wire \add_90_I36_L14036_C132/carry[4]  ;
wire \add_90_I36_L14036_C132/carry[3]  ;
wire \add_90_I36_L14036_C132/carry[2]  ;
wire \add_90_I35_L14036_C132/carry[5]  ;
wire \add_90_I35_L14036_C132/carry[4]  ;
wire \add_90_I35_L14036_C132/carry[3]  ;
wire \add_90_I35_L14036_C132/carry[2]  ;
wire \add_90_I34_L14036_C132/carry[5]  ;
wire \add_90_I34_L14036_C132/carry[4]  ;
wire \add_90_I34_L14036_C132/carry[3]  ;
wire \add_90_I34_L14036_C132/carry[2]  ;
wire \add_90_I33_L14036_C132/carry[5]  ;
wire \add_90_I33_L14036_C132/carry[4]  ;
wire \add_90_I33_L14036_C132/carry[3]  ;
wire \add_90_I33_L14036_C132/carry[2]  ;
wire \add_90_I32_L14036_C132/carry[5]  ;
wire \add_90_I32_L14036_C132/carry[4]  ;
wire \add_90_I32_L14036_C132/carry[3]  ;
wire \add_90_I32_L14036_C132/carry[2]  ;
wire \add_90_I31_L14036_C132/carry[5]  ;
wire \add_90_I31_L14036_C132/carry[4]  ;
wire \add_90_I31_L14036_C132/carry[3]  ;
wire \add_90_I31_L14036_C132/carry[2]  ;
wire \add_90_I30_L14036_C132/carry[5]  ;
wire \add_90_I30_L14036_C132/carry[4]  ;
wire \add_90_I30_L14036_C132/carry[3]  ;
wire \add_90_I30_L14036_C132/carry[2]  ;
wire \add_90_I29_L14036_C132/carry[5]  ;
wire \add_90_I29_L14036_C132/carry[4]  ;
wire \add_90_I29_L14036_C132/carry[3]  ;
wire \add_90_I29_L14036_C132/carry[2]  ;
wire \add_90_I28_L14036_C132/carry[5]  ;
wire \add_90_I28_L14036_C132/carry[4]  ;
wire \add_90_I28_L14036_C132/carry[3]  ;
wire \add_90_I28_L14036_C132/carry[2]  ;
wire \add_90_I27_L14036_C132/carry[5]  ;
wire \add_90_I27_L14036_C132/carry[4]  ;
wire \add_90_I27_L14036_C132/carry[3]  ;
wire \add_90_I27_L14036_C132/carry[2]  ;
wire \add_90_I26_L14036_C132/carry[5]  ;
wire \add_90_I26_L14036_C132/carry[4]  ;
wire \add_90_I26_L14036_C132/carry[3]  ;
wire \add_90_I26_L14036_C132/carry[2]  ;
wire \add_90_I25_L14036_C132/carry[5]  ;
wire \add_90_I25_L14036_C132/carry[4]  ;
wire \add_90_I25_L14036_C132/carry[3]  ;
wire \add_90_I25_L14036_C132/carry[2]  ;
wire \add_90_I24_L14036_C132/carry[5]  ;
wire \add_90_I24_L14036_C132/carry[4]  ;
wire \add_90_I24_L14036_C132/carry[3]  ;
wire \add_90_I24_L14036_C132/carry[2]  ;
wire \add_90_I23_L14036_C132/carry[5]  ;
wire \add_90_I23_L14036_C132/carry[4]  ;
wire \add_90_I23_L14036_C132/carry[3]  ;
wire \add_90_I23_L14036_C132/carry[2]  ;
wire \add_90_I22_L14036_C132/carry[5]  ;
wire \add_90_I22_L14036_C132/carry[4]  ;
wire \add_90_I22_L14036_C132/carry[3]  ;
wire \add_90_I22_L14036_C132/carry[2]  ;
wire \add_90_I21_L14036_C132/carry[5]  ;
wire \add_90_I21_L14036_C132/carry[4]  ;
wire \add_90_I21_L14036_C132/carry[3]  ;
wire \add_90_I21_L14036_C132/carry[2]  ;
wire \add_90_I20_L14036_C132/carry[5]  ;
wire \add_90_I20_L14036_C132/carry[4]  ;
wire \add_90_I20_L14036_C132/carry[3]  ;
wire \add_90_I20_L14036_C132/carry[2]  ;
wire \add_90_I19_L14036_C132/carry[5]  ;
wire \add_90_I19_L14036_C132/carry[4]  ;
wire \add_90_I19_L14036_C132/carry[3]  ;
wire \add_90_I19_L14036_C132/carry[2]  ;
wire \add_90_I18_L14036_C132/carry[5]  ;
wire \add_90_I18_L14036_C132/carry[4]  ;
wire \add_90_I18_L14036_C132/carry[3]  ;
wire \add_90_I18_L14036_C132/carry[2]  ;
wire \add_90_I17_L14036_C132/carry[5]  ;
wire \add_90_I17_L14036_C132/carry[4]  ;
wire \add_90_I17_L14036_C132/carry[3]  ;
wire \add_90_I17_L14036_C132/carry[2]  ;
wire \add_90_I16_L14036_C132/carry[5]  ;
wire \add_90_I16_L14036_C132/carry[4]  ;
wire \add_90_I16_L14036_C132/carry[3]  ;
wire \add_90_I16_L14036_C132/carry[2]  ;
wire \add_90_I15_L14036_C132/carry[5]  ;
wire \add_90_I15_L14036_C132/carry[4]  ;
wire \add_90_I15_L14036_C132/carry[3]  ;
wire \add_90_I15_L14036_C132/carry[2]  ;
wire \add_90_I14_L14036_C132/carry[5]  ;
wire \add_90_I14_L14036_C132/carry[4]  ;
wire \add_90_I14_L14036_C132/carry[3]  ;
wire \add_90_I14_L14036_C132/carry[2]  ;
wire \add_90_I13_L14036_C132/carry[5]  ;
wire \add_90_I13_L14036_C132/carry[4]  ;
wire \add_90_I13_L14036_C132/carry[3]  ;
wire \add_90_I13_L14036_C132/carry[2]  ;
wire \add_90_I12_L14036_C132/carry[5]  ;
wire \add_90_I12_L14036_C132/carry[4]  ;
wire \add_90_I12_L14036_C132/carry[3]  ;
wire \add_90_I12_L14036_C132/carry[2]  ;
wire \add_90_I11_L14036_C132/carry[5]  ;
wire \add_90_I11_L14036_C132/carry[4]  ;
wire \add_90_I11_L14036_C132/carry[3]  ;
wire \add_90_I11_L14036_C132/carry[2]  ;
wire \add_90_I10_L14036_C132/carry[5]  ;
wire \add_90_I10_L14036_C132/carry[4]  ;
wire \add_90_I10_L14036_C132/carry[3]  ;
wire \add_90_I10_L14036_C132/carry[2]  ;
wire \add_90_I9_L14036_C132/carry[5]  ;
wire \add_90_I9_L14036_C132/carry[4]  ;
wire \add_90_I9_L14036_C132/carry[3]  ;
wire \add_90_I9_L14036_C132/carry[2]  ;
wire \add_90_I8_L14036_C132/carry[5]  ;
wire \add_90_I8_L14036_C132/carry[4]  ;
wire \add_90_I8_L14036_C132/carry[3]  ;
wire \add_90_I8_L14036_C132/carry[2]  ;
wire \add_90_I7_L14036_C132/carry[4]  ;
wire \add_90_I7_L14036_C132/carry[3]  ;
wire \add_90_I7_L14036_C132/carry[2]  ;
wire \add_90_I6_L14036_C132/carry[2]  ;
wire \add_90_I6_L14036_C132/carry[3]  ;
wire \add_90_I5_L14036_C132/carry[2]  ;
wire \sub_0_root_add_0_root_add_148/carry[5]  ;
wire \sub_0_root_add_0_root_add_148/carry[4]  ;
wire \sub_0_root_add_0_root_add_148/carry[3]  ;
wire \sub_0_root_add_0_root_add_148/carry[2]  ;
wire \sub_0_root_add_0_root_add_148/carry[1]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n120 ;
wire n121 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n153 ;
wire n155 ;
wire n157 ;
wire n159 ;
wire n161 ;
wire n163 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n175 ;
wire n176 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n205 ;
wire n207 ;
wire n209 ;
wire n211 ;
wire n213 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n228 ;
wire n230 ;
wire n234 ;
wire n237 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n245 ;
wire n313 ;
wire n314 ;
wire n329 ;
wire n330 ;
wire n335 ;
wire n336 ;
wire n350 ;
wire n353 ;
wire n356 ;
wire n357 ;
wire n373 ;
wire n374 ;
wire n381 ;
wire n382 ;
wire n404 ;
wire n405 ;
wire n416 ;
wire n417 ;
wire n432 ;
wire n433 ;
wire n445 ;
wire n446 ;
wire n451 ;
wire n458 ;
wire n459 ;
wire n470 ;
wire n471 ;
wire n478 ;
wire n479 ;
wire n486 ;
wire n487 ;
wire n488 ;
wire n499 ;
wire n500 ;
wire n507 ;
wire n508 ;
wire n516 ;
wire n517 ;
wire n572 ;
wire n576 ;
wire n591 ;
wire n594 ;
wire n596 ;
wire n597 ;
wire n613 ;
wire n614 ;
wire n620 ;
wire n621 ;
wire n633 ;
wire n634 ;
wire n641 ;
wire n642 ;
wire n645 ;
wire n646 ;
wire n657 ;
wire n658 ;
wire n671 ;
wire n672 ;
wire n683 ;
wire n684 ;
wire n688 ;
wire n689 ;
wire n699 ;
wire n700 ;
wire n712 ;
wire n713 ;
wire n722 ;
wire n723 ;
wire n734 ;
wire n735 ;
wire n742 ;
wire n743 ;
wire n804 ;
wire n805 ;
wire n806 ;
wire n807 ;
wire n808 ;
wire n809 ;
wire n810 ;
wire n811 ;
wire n812 ;
wire n813 ;
wire n814 ;
wire n815 ;
wire n816 ;
wire n817 ;
wire n818 ;
wire n819 ;
wire n820 ;
wire n821 ;
wire n822 ;
wire n823 ;
wire n824 ;
wire n825 ;
wire n826 ;
wire n827 ;
wire n828 ;
wire n829 ;
wire n830 ;
wire n831 ;
wire n832 ;
wire n833 ;
wire n834 ;
wire n835 ;
wire n836 ;
wire n837 ;
wire n838 ;
wire n839 ;
wire n840 ;
wire n841 ;
wire n842 ;
wire n843 ;
wire n844 ;
wire n845 ;
wire n846 ;
wire n847 ;
wire n848 ;
wire n849 ;
wire n850 ;
wire n851 ;
wire n852 ;
wire n853 ;
wire n854 ;
wire n855 ;
wire n856 ;
wire n857 ;
wire n858 ;
wire n859 ;
wire n860 ;
wire n861 ;
wire n862 ;
wire n863 ;
wire n864 ;
wire n865 ;
wire n866 ;
wire n867 ;
wire n868 ;
wire n869 ;
wire n870 ;
wire n871 ;
wire n872 ;
wire n873 ;
wire n874 ;
wire n875 ;
wire n876 ;
wire n877 ;
wire n878 ;
wire n879 ;
wire n880 ;
wire n881 ;
wire n882 ;
wire n883 ;
wire n884 ;
wire n885 ;
wire n886 ;
wire n887 ;
wire n888 ;
wire n889 ;
wire n890 ;
wire n891 ;
wire n892 ;
wire n893 ;
wire n894 ;
wire n895 ;
wire n896 ;
wire n897 ;
wire n898 ;
wire n899 ;
wire n900 ;
wire n901 ;
wire n902 ;
wire n903 ;
wire n904 ;
wire n905 ;
wire n906 ;
wire n907 ;
wire n908 ;
wire n909 ;
wire n910 ;
wire n911 ;
wire n912 ;
wire n913 ;
wire n914 ;
wire n915 ;
wire n916 ;
wire n917 ;
wire n918 ;
wire n919 ;
wire n920 ;
wire n921 ;
wire n922 ;
wire n923 ;
wire n924 ;
wire n925 ;
wire n926 ;
wire n927 ;
wire n928 ;
wire n929 ;
wire n930 ;
wire n931 ;
wire n932 ;
wire n933 ;
wire n934 ;
wire n935 ;
wire n936 ;
wire n937 ;
wire n938 ;
wire n939 ;
wire n940 ;
wire n941 ;
wire n942 ;
wire n943 ;
wire n944 ;
wire n945 ;
wire n946 ;
wire n947 ;
wire n948 ;
wire n949 ;
wire n950 ;
wire n951 ;
wire n952 ;
wire n953 ;
wire n954 ;
wire n955 ;
wire n956 ;
wire n957 ;
wire n958 ;
wire n959 ;
wire n960 ;
wire n961 ;
wire n962 ;
wire n963 ;
wire n964 ;
wire n965 ;
wire n966 ;
wire n967 ;
wire n968 ;
wire n969 ;
wire n970 ;
wire n971 ;
wire n972 ;
wire n973 ;
wire n974 ;
wire n975 ;
wire n976 ;
wire n977 ;
wire n978 ;
wire n979 ;
wire n980 ;
wire n981 ;
wire n982 ;
wire n983 ;
wire n984 ;
wire n985 ;
wire n986 ;
wire n987 ;
wire n988 ;
wire n989 ;
wire n990 ;
wire n991 ;
wire n992 ;
wire n993 ;
wire n994 ;
wire n995 ;
wire n996 ;
wire n997 ;
wire n998 ;
wire n999 ;
wire n1000 ;
wire n1001 ;
wire n1002 ;
wire n1003 ;
wire n1004 ;
wire n1005 ;
wire n1006 ;
wire n1007 ;
wire n1008 ;
wire n1009 ;
wire n1010 ;
wire n1011 ;
wire n1012 ;
wire n1013 ;
wire n1014 ;
wire n1015 ;
wire n1016 ;
wire n1017 ;
wire n1018 ;
wire n1019 ;
wire n1020 ;
wire n1021 ;
wire n1022 ;
wire n1023 ;
wire n1024 ;
wire n1025 ;
wire n1026 ;
wire n1027 ;
wire n1028 ;
wire n1029 ;
wire n1030 ;
wire n1031 ;
wire n1032 ;
wire n1033 ;
wire n1034 ;
wire n1035 ;
wire n1036 ;
wire n1037 ;
wire n1038 ;
wire n1039 ;
wire n1040 ;
wire n1041 ;
wire n1042 ;
wire n1043 ;
wire n1044 ;
wire n1045 ;
wire n1046 ;
wire n1047 ;
wire n1048 ;
wire n1049 ;
wire n1050 ;
wire n1051 ;
wire n1052 ;
wire n1053 ;
wire n1054 ;
wire n1055 ;
wire n1056 ;
wire n1057 ;
wire n1058 ;
wire n1059 ;
wire n1060 ;
wire n1061 ;
wire n1062 ;
wire n1063 ;
wire n1064 ;
wire n1065 ;
wire n1066 ;
wire n1067 ;
wire n1068 ;
wire n1069 ;
wire n1070 ;
wire n1071 ;
wire n1072 ;
wire n1073 ;
wire n1074 ;
wire n1075 ;
wire n1076 ;
wire n1077 ;
wire n1078 ;
wire n1079 ;
wire n1080 ;
wire n1081 ;
wire n1082 ;
wire n1083 ;
wire n1084 ;
wire n1085 ;
wire n1086 ;
wire n1087 ;
wire n1088 ;
wire n1089 ;
wire n1090 ;
wire n1091 ;
wire n1092 ;
wire n1093 ;
wire n1094 ;
wire n1095 ;
wire n1096 ;
wire n1097 ;
wire n1098 ;
wire n1099 ;
wire n1100 ;
wire n1101 ;
wire n1102 ;
wire n1103 ;
wire n1104 ;
wire n1105 ;
wire n1106 ;
wire n1107 ;
wire n1108 ;
wire n1109 ;
wire n1110 ;
wire n1111 ;
wire n1112 ;
wire n1113 ;
wire n1114 ;
wire n1115 ;
wire n1116 ;
wire n1117 ;
wire n1118 ;
wire n1119 ;
wire n1120 ;
wire n1121 ;
wire n1122 ;
wire n1123 ;
wire n1124 ;
wire n1125 ;
wire n1126 ;
wire n1127 ;
wire n1128 ;
wire n1129 ;
wire n1130 ;
wire n1131 ;
wire n1132 ;
wire n1133 ;
wire n1134 ;
wire n1135 ;
wire n1136 ;
wire n1137 ;
wire n1138 ;
wire n1139 ;
wire n1140 ;
wire n1141 ;
wire n1142 ;
wire n1143 ;
wire n1144 ;
wire n1145 ;
wire n1146 ;
wire n1147 ;
wire n1148 ;
wire n1149 ;
wire n1150 ;
wire n1151 ;
wire n1152 ;
wire n1153 ;
wire n1154 ;
wire n1155 ;
wire n1156 ;
wire n1157 ;
wire n1158 ;
wire n1159 ;
wire n1160 ;
wire n1161 ;
wire n1162 ;
wire n1163 ;
wire n1164 ;
wire n1165 ;
wire n1166 ;
wire n1167 ;
wire n1168 ;
wire n1169 ;
wire n1170 ;
wire n1171 ;
wire n1172 ;
wire n1173 ;
wire n1174 ;
wire n1175 ;
wire n1176 ;
wire n1177 ;
wire n1178 ;
wire n1179 ;
wire n1180 ;
wire n1181 ;
wire n1182 ;
wire n1183 ;
wire n1184 ;
wire n1185 ;
wire n1186 ;
wire n1187 ;
wire n1188 ;
wire n1189 ;
wire n1190 ;
wire n1191 ;
wire n1192 ;
wire n1193 ;
wire n1194 ;
wire n1195 ;
wire n1196 ;
wire n1197 ;
wire n1198 ;
wire n1199 ;
wire n1200 ;
wire n1201 ;
wire n1202 ;
wire n1203 ;
wire n1204 ;
wire n1205 ;
wire n1206 ;
wire n1207 ;
wire n1208 ;
wire n1209 ;
wire n1210 ;
wire n1211 ;
wire n1212 ;
wire n1213 ;
wire n1214 ;
wire n1215 ;
wire n1216 ;
wire n1217 ;
wire n1218 ;
wire n1219 ;
wire n1220 ;
wire n1221 ;
wire n1222 ;
wire n1223 ;
wire n1224 ;
wire n1225 ;
wire n1226 ;
wire n1227 ;
wire n1228 ;
wire n1229 ;
wire n1230 ;
wire n1231 ;
wire n1232 ;
wire n1233 ;
wire n1234 ;
wire n1235 ;
wire n1236 ;
wire n1237 ;
wire n1238 ;
wire n1239 ;
wire n1240 ;
wire n1241 ;
wire n1242 ;
wire n1243 ;
wire n1244 ;
wire n1245 ;
wire n1246 ;
wire n1247 ;
wire n1248 ;
wire n1249 ;
wire n1250 ;
wire n1251 ;
wire n1252 ;
wire n1253 ;
wire n1254 ;
wire n1255 ;
wire n1256 ;
wire n1257 ;
wire n1258 ;
wire n1259 ;
wire n1260 ;
wire n1261 ;
wire n1262 ;
wire n1263 ;
wire n1264 ;
wire n1265 ;
wire n1266 ;
wire n1267 ;
wire n1268 ;
wire n1269 ;
wire n1270 ;
wire n1271 ;
wire n1272 ;
wire n1273 ;
wire n1274 ;
wire n1275 ;
wire n1276 ;
wire n1277 ;
wire n1278 ;
wire n1279 ;
wire n1280 ;
wire n1281 ;
wire n1282 ;
wire n1283 ;
wire n1284 ;
wire n1285 ;
wire n1286 ;
wire n1287 ;
wire n1288 ;
wire n1289 ;
wire n1290 ;
wire n1291 ;
wire n1292 ;
wire n1293 ;
wire n1294 ;
wire n1295 ;
wire n1296 ;
wire n1297 ;
wire n1298 ;
wire n1299 ;
wire n1300 ;
wire n1301 ;
wire n1302 ;
wire n1303 ;
wire n1304 ;
wire n1305 ;
wire n1306 ;
wire n1307 ;
wire n1308 ;
wire n1309 ;
wire n1310 ;
wire n1311 ;
wire n1312 ;
wire n1313 ;
wire n1314 ;
wire n1315 ;
wire n1316 ;
wire n1317 ;
wire n1318 ;
wire n1319 ;
wire n1320 ;
wire n1321 ;
wire n1322 ;
wire n1323 ;
wire n1324 ;
wire n1325 ;
wire n1326 ;
wire n1327 ;
wire n1328 ;
wire n1329 ;
wire n1330 ;
wire n1331 ;
wire n1332 ;
wire n1333 ;
wire n1334 ;
wire n1335 ;
wire n1336 ;
wire n1337 ;
wire n1338 ;
wire n1339 ;
wire n1340 ;
wire n1341 ;
wire n1342 ;
wire n1343 ;
wire n1344 ;
wire n1345 ;
wire n1346 ;
wire n1347 ;
wire n1348 ;
wire n1349 ;
wire n1350 ;
wire n1351 ;
wire n1352 ;
wire n1353 ;
wire n1354 ;
wire n1355 ;
wire n1356 ;
wire n1357 ;
wire n1358 ;
wire n1359 ;
wire n1360 ;
wire n1361 ;
wire n1362 ;
wire n1363 ;
wire n1364 ;
wire n1365 ;
wire n1366 ;
wire n1367 ;
wire n1368 ;
wire n1369 ;
wire n1370 ;
wire n1371 ;
wire n1372 ;
wire n1373 ;
wire n1374 ;
wire n1375 ;
wire n1376 ;
wire n1377 ;
wire n1378 ;
wire n1379 ;
wire n1380 ;
wire n1381 ;
wire n1382 ;
wire n1383 ;
wire n1384 ;
wire n1385 ;
wire n1386 ;
wire n1387 ;
wire n1388 ;
wire n1389 ;
wire n1390 ;
wire n1391 ;
wire n1392 ;
wire n1393 ;
wire n1394 ;
wire n1395 ;
wire n1396 ;
wire n1397 ;
wire n1398 ;
wire n1399 ;
wire n1400 ;
wire n1401 ;
wire n1402 ;
wire n1403 ;
wire n1404 ;
wire n1405 ;
wire n1406 ;
wire n1407 ;
wire n1408 ;
wire n1409 ;
wire n1410 ;
wire n1411 ;
wire n1412 ;
wire n1413 ;
wire n1414 ;
wire n1415 ;
wire n1416 ;
wire n1417 ;
wire n1418 ;
wire n1419 ;
wire n1420 ;
wire n1421 ;
wire n1422 ;
wire n1423 ;
wire n1424 ;
wire n1425 ;
wire n1426 ;
wire n1427 ;
wire n1428 ;
wire n1429 ;
wire n1430 ;
wire n1431 ;
wire n1432 ;
wire n1433 ;
wire n1434 ;
wire n1435 ;
wire n1436 ;
wire n1437 ;
wire n1438 ;
wire n1439 ;
wire n1440 ;
wire n1441 ;
wire n1442 ;
wire n1443 ;
wire n1444 ;
wire n1445 ;
wire n1446 ;
wire n1447 ;
wire n1448 ;
wire n1449 ;
wire n1450 ;
wire n1451 ;
wire n1452 ;
wire n1453 ;
wire n1454 ;
wire n1455 ;
wire n1456 ;
wire n1457 ;
wire n1458 ;
wire n1459 ;
wire n1460 ;
wire n1461 ;
wire n1462 ;
wire n1463 ;
wire n1464 ;
wire n1465 ;
wire n1466 ;
wire n1467 ;
wire n1468 ;
wire n1469 ;
wire n1470 ;
wire n1471 ;
wire n1472 ;
wire n1473 ;
wire n1474 ;
wire n1475 ;
wire n1476 ;
wire n1477 ;
wire n1478 ;
wire n1479 ;
wire n1480 ;
wire n1481 ;
wire n1482 ;
wire n1483 ;
wire n1484 ;
wire n1485 ;
wire n1486 ;
wire n1487 ;
wire n1488 ;
wire n1489 ;
wire n1490 ;
wire n1491 ;
wire n1492 ;
wire n1493 ;
wire n1494 ;
wire n1495 ;
wire n1496 ;
wire n1497 ;
wire n1498 ;
wire n1499 ;
wire n1500 ;
wire n1501 ;
wire n1502 ;
wire n1503 ;
wire n1504 ;
wire n1505 ;
wire n1506 ;
wire n1507 ;
wire n1508 ;
wire n1509 ;
wire n1510 ;
wire n1511 ;
wire n1512 ;
wire n1513 ;
wire n1514 ;
wire n1515 ;
wire n1516 ;
wire n1517 ;
wire n1518 ;
wire n1519 ;
wire n1520 ;
wire n1521 ;
wire n1522 ;
wire n1523 ;
wire n1524 ;
wire n1525 ;
wire n1526 ;
wire n1527 ;
wire n1528 ;
wire n1529 ;
wire n1530 ;
wire n1531 ;
wire n1532 ;
wire n1533 ;
wire n1534 ;
wire n1535 ;
wire n1536 ;
wire n1537 ;
wire n1538 ;
wire n1539 ;
wire n1540 ;
wire n1541 ;
wire n1542 ;
wire n1543 ;
wire n1544 ;
wire n1545 ;
wire n1546 ;
wire n1547 ;
wire n1548 ;
wire n1549 ;
wire n1550 ;
wire n1551 ;
wire n1552 ;
wire n1553 ;
wire n1554 ;
wire n1555 ;
wire n1556 ;
wire n1557 ;
wire n1558 ;
wire n1559 ;
wire n1560 ;
wire n1561 ;
wire n1562 ;
wire n1563 ;
wire n1564 ;
wire n1565 ;
wire n1566 ;
wire n1567 ;
wire n1568 ;
wire n1569 ;
wire n1570 ;
wire n1571 ;
wire n1572 ;
wire n1573 ;
wire n1574 ;
wire n1575 ;
wire n1576 ;
wire n1577 ;
wire n1578 ;
wire n1579 ;
wire n1580 ;
wire n1581 ;
wire n1582 ;
wire n1583 ;
wire n1584 ;
wire n1585 ;
wire n1586 ;
wire n1587 ;
wire n1588 ;
wire n1589 ;
wire n1590 ;
wire n1591 ;
wire n1592 ;
wire n1593 ;
wire n1594 ;
wire n1595 ;
wire n1596 ;
wire n1597 ;
wire n1598 ;
wire n1599 ;
wire n1600 ;
wire n1601 ;
wire n1602 ;
wire n1603 ;
wire n1604 ;
wire n1605 ;
wire n1606 ;
wire n1607 ;
wire n1608 ;
wire n1609 ;
wire n1610 ;
wire n1611 ;
wire n1612 ;
wire n1613 ;
wire n1614 ;
wire n1615 ;
wire n1616 ;
wire n1617 ;
wire n1618 ;
wire n1619 ;
wire n1620 ;
wire n1621 ;
wire n1622 ;
wire n1623 ;
wire n1624 ;
wire n1625 ;
wire n1626 ;
wire n1627 ;
wire n1628 ;
wire n1629 ;
wire n1630 ;
wire n1631 ;
wire n1632 ;
wire n1633 ;
wire n1634 ;
wire n1635 ;
wire n1636 ;
wire n1637 ;
wire n1638 ;
wire n1639 ;
wire n1640 ;
wire n1641 ;
wire n1642 ;
wire n1643 ;
wire n1644 ;
wire n1645 ;
wire n1646 ;
wire n1647 ;
wire n1648 ;
wire n1649 ;
wire n1650 ;
wire n1651 ;
wire n1652 ;
wire n1653 ;
wire n1654 ;
wire n1655 ;
wire n1656 ;
wire n1657 ;
wire n1658 ;
wire n1659 ;
wire n1660 ;
wire n1661 ;
wire n1662 ;
wire n1663 ;
wire n1664 ;
wire n1665 ;
wire n1666 ;
wire n1667 ;
wire n1668 ;
wire n1669 ;
wire n1670 ;
wire n1671 ;
wire n1672 ;
wire n1673 ;
wire n1674 ;
wire n1675 ;
wire n1676 ;
wire n1677 ;
wire n1678 ;
wire n1679 ;
wire n1680 ;
wire n1681 ;
wire n1682 ;
wire n1683 ;
wire n1684 ;
wire n1685 ;
wire n1686 ;
wire n1687 ;
wire n1688 ;
wire n1689 ;
wire n1690 ;
wire n1691 ;
wire n1692 ;
wire n1693 ;
wire n1694 ;
wire n1695 ;
wire n1696 ;
wire n1697 ;
wire n1698 ;
wire n1699 ;
wire n1700 ;
wire n1701 ;
wire n1702 ;
wire n1703 ;
wire n1704 ;
wire n1705 ;
wire n1706 ;
wire n1707 ;
wire n1708 ;
wire n1709 ;
wire n1710 ;
wire n1711 ;
wire n1712 ;
wire n1713 ;
wire n1714 ;
wire n1715 ;
wire n1716 ;
wire n1717 ;
wire n1718 ;
wire n1719 ;
wire n1720 ;
wire n1721 ;
wire n1722 ;
wire n1723 ;
wire n1724 ;
wire n1725 ;
wire n1726 ;
wire n1727 ;
wire n1728 ;
wire n1729 ;
wire n1730 ;
wire n1731 ;
wire n1732 ;
wire n1733 ;
wire n1734 ;
wire n1735 ;
wire n1736 ;
wire n1737 ;
wire n1738 ;
wire n1739 ;
wire n1740 ;
wire n1741 ;
wire n1742 ;
wire n1743 ;
wire n1744 ;
wire n1745 ;
wire n1746 ;
wire n1747 ;
wire n1748 ;
wire n1749 ;
wire n1750 ;
wire n1751 ;
wire n1752 ;
wire n1753 ;
wire n1754 ;
wire n1755 ;
wire n1756 ;
wire n1757 ;
wire n1758 ;
wire n1759 ;
wire n1760 ;
wire n1761 ;
wire n1762 ;
wire n1763 ;
wire n1764 ;
wire n1765 ;
wire n1766 ;
wire n1767 ;
wire n1768 ;
wire n1769 ;
wire n1770 ;
wire n1771 ;
wire n1772 ;
wire n1773 ;
wire n1774 ;
wire n1775 ;
wire n1776 ;
wire n1777 ;
wire n1778 ;
wire n1779 ;
wire n1780 ;
wire n1781 ;
wire n1782 ;
wire n1783 ;
wire n1784 ;
wire n1785 ;
wire n1786 ;
wire n1787 ;
wire n1788 ;
wire n1789 ;
wire n1790 ;
wire n1791 ;
wire n1792 ;
wire n1793 ;
wire n1794 ;
wire n1795 ;
wire n1796 ;
wire n1797 ;
wire n1798 ;
wire n1799 ;
wire n1800 ;
wire n1801 ;
wire n1802 ;
wire n1803 ;
wire n1804 ;
wire n1805 ;
wire n1806 ;
wire n1807 ;
wire n1808 ;
wire n1809 ;
wire n1810 ;
wire n1811 ;
wire n1812 ;
wire n1813 ;
wire n1814 ;
wire n1815 ;
wire n1816 ;
wire n1817 ;
wire n1818 ;
wire n1819 ;
wire n1820 ;
wire n1821 ;
wire n1822 ;
wire n1823 ;
wire n1824 ;
wire n1825 ;
wire n1826 ;
wire n1827 ;
wire n1828 ;
wire n1829 ;
wire n1830 ;
wire n1831 ;
wire n1832 ;
wire n1833 ;
wire n1834 ;
wire n1835 ;
wire n1836 ;
wire n1837 ;
wire n1838 ;
wire n1839 ;
wire n1840 ;
wire n1841 ;
wire n1842 ;
wire n1843 ;
wire n1844 ;
wire n1845 ;
wire n1846 ;
wire n1847 ;
wire n1848 ;
wire n1849 ;
wire n1850 ;
wire n1851 ;
wire n1852 ;
wire n1853 ;
wire n1854 ;
wire n1855 ;
wire n1856 ;
wire n1857 ;
wire n1858 ;
wire n1859 ;
wire n1860 ;
wire n1861 ;
wire n1862 ;
wire n1863 ;
wire n1864 ;
wire n1865 ;
wire n1866 ;
wire n1867 ;
wire n1868 ;
wire n1869 ;
wire n1870 ;
wire n1871 ;
wire n1872 ;
wire n1873 ;
wire n1874 ;
wire n1875 ;
wire n1876 ;
wire n1877 ;
wire n1878 ;
wire n1879 ;
wire n1880 ;
wire n1881 ;
wire n1882 ;
wire n1883 ;
wire n1884 ;
wire n1885 ;
wire n1886 ;
wire n1887 ;
wire n1888 ;
wire n1889 ;
wire n1890 ;
wire n1891 ;
wire n1892 ;
wire n1893 ;
wire n1894 ;
wire n1895 ;
wire n1896 ;
wire n1897 ;
wire n1898 ;
wire n1899 ;
wire n1900 ;
wire n1901 ;
wire n1902 ;
wire n1903 ;
wire n1904 ;
wire n1905 ;
wire n1906 ;
wire n1907 ;
wire n1908 ;
wire n1909 ;
wire n1910 ;
wire n1911 ;
wire n1912 ;
wire n1913 ;
wire n1914 ;
wire n1915 ;
wire n1916 ;
wire n1917 ;
wire n1918 ;
wire n1919 ;
wire n1920 ;
wire n1921 ;
wire n1922 ;
wire n1923 ;
wire n1924 ;
wire n1925 ;
wire n1926 ;
wire n1927 ;
wire n1928 ;
wire n1929 ;
wire n1930 ;
wire n1931 ;
wire n1932 ;
wire n1933 ;
wire n1934 ;
wire n1935 ;
wire n1936 ;
wire n1937 ;
wire n1938 ;
wire n1939 ;
wire n1940 ;
wire n1941 ;
wire n1942 ;
wire n1943 ;
wire n1944 ;
wire n1945 ;
wire n1946 ;
wire n1947 ;
wire n1948 ;
wire n1949 ;
wire n1950 ;
wire n1951 ;
wire n1952 ;
wire n1953 ;
wire n1954 ;
wire n1955 ;
wire n1956 ;
wire n1957 ;
wire n1958 ;
wire n1959 ;
wire n1960 ;
wire n1961 ;
wire n1962 ;
wire n1963 ;
wire n1964 ;
wire n1965 ;
wire n1966 ;
wire n1967 ;
wire n1968 ;
wire n1969 ;
wire n1970 ;
wire n1971 ;
wire n1972 ;
wire n1973 ;
wire n1974 ;
wire n1975 ;
wire n1976 ;
wire n1977 ;
wire n1978 ;
wire n1979 ;
wire n1980 ;
wire n1981 ;
wire n1982 ;
wire n1983 ;
wire n1984 ;
wire n1985 ;
wire n1986 ;
wire n1987 ;
wire n1988 ;
wire n1989 ;
wire n1990 ;
wire n1991 ;
wire n1992 ;
wire n1993 ;
wire n1994 ;
wire n1995 ;
wire n1996 ;
wire n1997 ;
wire n1998 ;
wire n1999 ;
wire n2000 ;
wire n2001 ;
wire n2002 ;
wire n2003 ;
wire n2004 ;
wire n2005 ;
wire n2006 ;
wire n2007 ;
wire [30:0] s_opa_i ;
wire [30:0] s_opb_i ;
wire [7:0] s_expa ;
wire [7:0] s_expb ;
wire [9:0] s_exp_10_i ;
wire [47:0] s_fract_48_i ;
wire [31:0] s_output_o ;
wire [5:0] s_zeros ;
wire [5:0] s_r_zeros ;
wire [9:0] s_exp_10a ;
wire [9:0] s_exp_10b ;
wire [8:0] s_expo1 ;
wire [5:0] s_shr2 ;
wire [5:0] s_shl2 ;
wire [47:0] s_frac2a ;
wire [8:0] s_expo2b ;
wire [24:0] s_frac_rnd ;
// instances
  DFFX1 desc876(.D(opa_i[30:30]),.CLK(clk_i),.QN(n1158));
  DFFX1 desc877(.D(opa_i[29:29]),.CLK(clk_i),.QN(n1159));
  DFFX1 desc878(.D(opa_i[28:28]),.CLK(clk_i),.QN(n1160));
  DFFX1 desc879(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_opa_i[27:27]));
  DFFX1 desc880(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_opa_i[26:26]));
  DFFX1 desc881(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_opa_i[25:25]));
  DFFX1 desc882(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_opa_i[24:24]));
  DFFX1 desc883(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_opa_i[23:23]));
  DFFX1 desc884(.D(opa_i[22:22]),.CLK(clk_i),.QN(n1166));
  DFFX1 desc885(.D(opa_i[21:21]),.CLK(clk_i),.Q(s_opa_i[21:21]));
  DFFX1 desc886(.D(opa_i[20:20]),.CLK(clk_i),.Q(s_opa_i[20:20]));
  DFFX1 desc887(.D(opa_i[19:19]),.CLK(clk_i),.QN(n1152));
  DFFX1 desc888(.D(opa_i[18:18]),.CLK(clk_i),.QN(n1153));
  DFFX1 desc889(.D(opa_i[17:17]),.CLK(clk_i),.QN(n1154));
  DFFX1 desc890(.D(opa_i[16:16]),.CLK(clk_i),.Q(s_opa_i[16:16]));
  DFFX1 desc891(.D(opa_i[15:15]),.CLK(clk_i),.Q(s_opa_i[15:15]));
  DFFX1 desc892(.D(opa_i[14:14]),.CLK(clk_i),.Q(s_opa_i[14:14]));
  DFFX1 desc893(.D(opa_i[13:13]),.CLK(clk_i),.Q(s_opa_i[13:13]));
  DFFX1 desc894(.D(opa_i[12:12]),.CLK(clk_i),.Q(s_opa_i[12:12]));
  DFFX1 desc895(.D(opa_i[11:11]),.CLK(clk_i),.Q(s_opa_i[11:11]));
  DFFX1 desc896(.D(opa_i[10:10]),.CLK(clk_i),.QN(n1176));
  DFFX1 desc897(.D(opa_i[9:9]),.CLK(clk_i),.QN(n1167));
  DFFX1 desc898(.D(opa_i[8:8]),.CLK(clk_i),.QN(n1168));
  DFFX1 desc899(.D(opa_i[7:7]),.CLK(clk_i),.QN(n1169));
  DFFX1 desc900(.D(opa_i[6:6]),.CLK(clk_i),.Q(s_opa_i[6:6]));
  DFFX1 desc901(.D(opa_i[5:5]),.CLK(clk_i),.Q(s_opa_i[5:5]));
  DFFX1 desc902(.D(opa_i[4:4]),.CLK(clk_i),.Q(s_opa_i[4:4]));
  DFFX1 desc903(.D(opa_i[3:3]),.CLK(clk_i),.QN(n1164));
  DFFX1 desc904(.D(opa_i[2:2]),.CLK(clk_i),.QN(n1165));
  DFFX1 desc905(.D(opa_i[1:1]),.CLK(clk_i),.Q(s_opa_i[1:1]));
  DFFX1 desc906(.D(opa_i[0:0]),.CLK(clk_i),.QN(n1177));
  DFFX1 desc907(.D(opb_i[30:30]),.CLK(clk_i),.QN(n1161));
  DFFX1 desc908(.D(opb_i[29:29]),.CLK(clk_i),.QN(n1162));
  DFFX1 desc909(.D(opb_i[28:28]),.CLK(clk_i),.QN(n1163));
  DFFX1 desc910(.D(opb_i[27:27]),.CLK(clk_i),.Q(s_opb_i[27:27]));
  DFFX1 desc911(.D(opb_i[26:26]),.CLK(clk_i),.Q(s_opb_i[26:26]));
  DFFX1 desc912(.D(opb_i[25:25]),.CLK(clk_i),.Q(s_opb_i[25:25]));
  DFFX1 desc913(.D(opb_i[24:24]),.CLK(clk_i),.Q(s_opb_i[24:24]));
  DFFX1 desc914(.D(opb_i[23:23]),.CLK(clk_i),.Q(s_opb_i[23:23]));
  DFFX1 desc915(.D(opb_i[22:22]),.CLK(clk_i),.QN(n1172));
  DFFX1 desc916(.D(opb_i[21:21]),.CLK(clk_i),.Q(s_opb_i[21:21]));
  DFFX1 desc917(.D(opb_i[20:20]),.CLK(clk_i),.Q(s_opb_i[20:20]));
  DFFX1 desc918(.D(opb_i[19:19]),.CLK(clk_i),.QN(n1155));
  DFFX1 desc919(.D(opb_i[18:18]),.CLK(clk_i),.QN(n1156));
  DFFX1 desc920(.D(opb_i[17:17]),.CLK(clk_i),.QN(n1157));
  DFFX1 desc921(.D(opb_i[16:16]),.CLK(clk_i),.Q(s_opb_i[16:16]));
  DFFX1 desc922(.D(opb_i[15:15]),.CLK(clk_i),.Q(s_opb_i[15:15]));
  DFFX1 desc923(.D(opb_i[14:14]),.CLK(clk_i),.Q(s_opb_i[14:14]));
  DFFX1 desc924(.D(opb_i[13:13]),.CLK(clk_i),.Q(s_opb_i[13:13]));
  DFFX1 desc925(.D(opb_i[12:12]),.CLK(clk_i),.Q(s_opb_i[12:12]));
  DFFX1 desc926(.D(opb_i[11:11]),.CLK(clk_i),.Q(s_opb_i[11:11]));
  DFFX1 desc927(.D(opb_i[10:10]),.CLK(clk_i),.QN(n1178));
  DFFX1 desc928(.D(opb_i[9:9]),.CLK(clk_i),.QN(n1173));
  DFFX1 desc929(.D(opb_i[8:8]),.CLK(clk_i),.QN(n1174));
  DFFX1 desc930(.D(opb_i[7:7]),.CLK(clk_i),.QN(n1175));
  DFFX1 desc931(.D(opb_i[6:6]),.CLK(clk_i),.Q(s_opb_i[6:6]));
  DFFX1 desc932(.D(opb_i[5:5]),.CLK(clk_i),.Q(s_opb_i[5:5]));
  DFFX1 desc933(.D(opb_i[4:4]),.CLK(clk_i),.Q(s_opb_i[4:4]));
  DFFX1 desc934(.D(opb_i[3:3]),.CLK(clk_i),.QN(n1170));
  DFFX1 desc935(.D(opb_i[2:2]),.CLK(clk_i),.QN(n1171));
  DFFX1 desc936(.D(opb_i[1:1]),.CLK(clk_i),.Q(s_opb_i[1:1]));
  DFFX1 desc937(.D(opb_i[0:0]),.CLK(clk_i),.QN(n1179));
  DFFX1 desc938(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_expa[7:7]));
  DFFX1 desc939(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_expa[6:6]));
  DFFX1 desc940(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_expa[5:5]));
  DFFX1 desc941(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_expa[4:4]));
  DFFX1 desc942(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_expa[3:3]));
  DFFX1 desc943(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_expa[2:2]));
  DFFX1 desc944(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_expa[1:1]));
  DFFX1 desc945(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_expa[0:0]));
  DFFX1 desc946(.D(opb_i[30:30]),.CLK(clk_i),.Q(s_expb[7:7]));
  DFFX1 desc947(.D(opb_i[29:29]),.CLK(clk_i),.Q(s_expb[6:6]));
  DFFX1 desc948(.D(opb_i[28:28]),.CLK(clk_i),.Q(s_expb[5:5]));
  DFFX1 desc949(.D(opb_i[27:27]),.CLK(clk_i),.Q(s_expb[4:4]));
  DFFX1 desc950(.D(opb_i[26:26]),.CLK(clk_i),.Q(s_expb[3:3]));
  DFFX1 desc951(.D(opb_i[25:25]),.CLK(clk_i),.Q(s_expb[2:2]));
  DFFX1 desc952(.D(opb_i[24:24]),.CLK(clk_i),.Q(s_expb[1:1]));
  DFFX1 desc953(.D(opb_i[23:23]),.CLK(clk_i),.Q(s_expb[0:0]));
  DFFX1 desc954(.D(exp_10_i[9:9]),.CLK(clk_i),.QN(n1198));
  DFFX1 desc955(.D(exp_10_i[8:8]),.CLK(clk_i),.Q(s_exp_10_i[8:8]));
  DFFX1 desc956(.D(exp_10_i[7:7]),.CLK(clk_i),.Q(s_exp_10_i[7:7]));
  DFFX1 desc957(.D(exp_10_i[6:6]),.CLK(clk_i),.Q(s_exp_10_i[6:6]));
  DFFX1 desc958(.D(exp_10_i[5:5]),.CLK(clk_i),.Q(s_exp_10_i[5:5]));
  DFFX1 desc959(.D(exp_10_i[4:4]),.CLK(clk_i),.Q(s_exp_10_i[4:4]));
  DFFX1 desc960(.D(exp_10_i[3:3]),.CLK(clk_i),.Q(s_exp_10_i[3:3]));
  DFFX1 desc961(.D(exp_10_i[2:2]),.CLK(clk_i),.Q(s_exp_10_i[2:2]));
  DFFX1 desc962(.D(exp_10_i[1:1]),.CLK(clk_i),.Q(s_exp_10_i[1:1]));
  DFFX1 desc963(.D(exp_10_i[0:0]),.CLK(clk_i),.Q(s_exp_10_i[0:0]));
  DFFX1 desc964(.D(fract_48_i[47:47]),.CLK(clk_i),.Q(N2993),.QN(n68));
  DFFX1 desc965(.D(fract_48_i[46:46]),.CLK(clk_i),.Q(s_fract_48_i[46:46]),.QN(n69));
  DFFX1 desc966(.D(fract_48_i[45:45]),.CLK(clk_i),.Q(s_fract_48_i[45:45]),.QN(n118));
  DFFX1 desc967(.D(fract_48_i[43:43]),.CLK(clk_i),.Q(s_fract_48_i[43:43]),.QN(n122));
  DFFX1 desc968(.D(fract_48_i[41:41]),.CLK(clk_i),.Q(s_fract_48_i[41:41]),.QN(n130));
  DFFX1 desc969(.D(fract_48_i[40:40]),.CLK(clk_i),.Q(s_fract_48_i[40:40]),.QN(n137));
  DFFX1 desc970(.D(fract_48_i[39:39]),.CLK(clk_i),.Q(s_fract_48_i[39:39]),.QN(n144));
  DFFX1 desc971(.D(fract_48_i[38:38]),.CLK(clk_i),.Q(s_fract_48_i[38:38]),.QN(n145));
  DFFX1 desc972(.D(fract_48_i[37:37]),.CLK(clk_i),.Q(s_fract_48_i[37:37]),.QN(n146));
  DFFX1 desc973(.D(fract_48_i[35:35]),.CLK(clk_i),.Q(s_fract_48_i[35:35]),.QN(n154));
  DFFX1 desc974(.D(fract_48_i[34:34]),.CLK(clk_i),.Q(s_fract_48_i[34:34]),.QN(n156));
  DFFX1 desc975(.D(fract_48_i[33:33]),.CLK(clk_i),.Q(s_fract_48_i[33:33]),.QN(n158));
  DFFX1 desc976(.D(fract_48_i[32:32]),.CLK(clk_i),.Q(s_fract_48_i[32:32]),.QN(n160));
  DFFX1 desc977(.D(fract_48_i[31:31]),.CLK(clk_i),.Q(s_fract_48_i[31:31]),.QN(n162));
  DFFX1 desc978(.D(fract_48_i[29:29]),.CLK(clk_i),.Q(s_fract_48_i[29:29]),.QN(n170));
  DFFX1 desc979(.D(fract_48_i[28:28]),.CLK(clk_i),.Q(s_fract_48_i[28:28]),.QN(n171));
  DFFX1 desc980(.D(fract_48_i[27:27]),.CLK(clk_i),.Q(s_fract_48_i[27:27]),.QN(n172));
  DFFX1 desc981(.D(fract_48_i[26:26]),.CLK(clk_i),.Q(s_fract_48_i[26:26]),.QN(n173));
  DFFX1 desc982(.D(fract_48_i[25:25]),.CLK(clk_i),.Q(s_fract_48_i[25:25]),.QN(n174));
  DFFX1 desc983(.D(fract_48_i[23:23]),.CLK(clk_i),.Q(s_fract_48_i[23:23]),.QN(n182));
  DFFX1 desc984(.D(fract_48_i[22:22]),.CLK(clk_i),.Q(s_fract_48_i[22:22]),.QN(n189));
  DFFX1 desc985(.D(fract_48_i[21:21]),.CLK(clk_i),.Q(s_fract_48_i[21:21]),.QN(n196));
  DFFX1 desc986(.D(fract_48_i[20:20]),.CLK(clk_i),.Q(s_fract_48_i[20:20]),.QN(n197));
  DFFX1 desc987(.D(fract_48_i[19:19]),.CLK(clk_i),.Q(s_fract_48_i[19:19]),.QN(n198));
  DFFX1 desc988(.D(fract_48_i[17:17]),.CLK(clk_i),.Q(s_fract_48_i[17:17]),.QN(n206));
  DFFX1 desc989(.D(fract_48_i[16:16]),.CLK(clk_i),.Q(s_fract_48_i[16:16]),.QN(n208));
  DFFX1 desc990(.D(fract_48_i[15:15]),.CLK(clk_i),.Q(s_fract_48_i[15:15]),.QN(n210));
  DFFX1 desc991(.D(fract_48_i[14:14]),.CLK(clk_i),.Q(s_fract_48_i[14:14]),.QN(n212));
  DFFX1 desc992(.D(fract_48_i[13:13]),.CLK(clk_i),.Q(s_fract_48_i[13:13]),.QN(n214));
  DFFX1 desc993(.D(fract_48_i[11:11]),.CLK(clk_i),.Q(s_fract_48_i[11:11]),.QN(n221));
  DFFX1 desc994(.D(fract_48_i[10:10]),.CLK(clk_i),.Q(s_fract_48_i[10:10]),.QN(n222));
  DFFX1 desc995(.D(fract_48_i[9:9]),.CLK(clk_i),.Q(s_fract_48_i[9:9]),.QN(n223));
  DFFX1 desc996(.D(fract_48_i[8:8]),.CLK(clk_i),.Q(s_fract_48_i[8:8]),.QN(n224));
  DFFX1 desc997(.D(fract_48_i[7:7]),.CLK(clk_i),.Q(s_fract_48_i[7:7]),.QN(n225));
  DFFX1 desc998(.D(fract_48_i[4:4]),.CLK(clk_i),.Q(s_fract_48_i[4:4]),.QN(n229));
  DFFX1 desc999(.D(fract_48_i[3:3]),.CLK(clk_i),.Q(s_fract_48_i[3:3]),.QN(n231));
  DFFX1 desc1000(.D(fract_48_i[0:0]),.CLK(clk_i),.Q(s_fract_48_i[0:0]),.QN(n233));
  DFFX1 s_sign_i_reg(.D(sign_i),.CLK(clk_i),.Q(s_output_o[31:31]));
  DFFX1 desc1001(.D(rmode_i[1:1]),.CLK(clk_i),.Q(\s_rmode_i[1] ),.QN(n235));
  DFFX1 desc1002(.D(rmode_i[0:0]),.CLK(clk_i),.QN(n236));
  DFFX1 desc1003(.D(s_output_o[31:31]),.CLK(clk_i),.Q(output_o[31:31]));
  DFFX1 desc1004(.D(N1637),.CLK(clk_i),.Q(s_zeros[5:5]));
  DFFX1 desc1005(.D(N1636),.CLK(clk_i),.Q(s_zeros[4:4]));
  DFFX1 desc1006(.D(N1635),.CLK(clk_i),.Q(s_zeros[3:3]));
  DFFX1 desc1007(.D(N1634),.CLK(clk_i),.Q(s_zeros[2:2]));
  DFFX1 desc1008(.D(N1633),.CLK(clk_i),.Q(s_zeros[1:1]));
  DFFX1 desc1009(.D(N1632),.CLK(clk_i),.Q(s_zeros[0:0]));
  DFFX1 desc1010(.D(N2979),.CLK(clk_i),.Q(s_r_zeros[5:5]),.QN(n54));
  DFFX1 desc1011(.D(N2978),.CLK(clk_i),.Q(s_r_zeros[4:4]),.QN(n78));
  DFFX1 desc1012(.D(N2977),.CLK(clk_i),.Q(s_r_zeros[3:3]),.QN(n74));
  DFFX1 desc1013(.D(N2976),.CLK(clk_i),.Q(s_r_zeros[2:2]));
  DFFX1 desc1014(.D(N2975),.CLK(clk_i),.Q(s_r_zeros[1:1]),.QN(n75));
  DFFX1 desc1015(.D(N2974),.CLK(clk_i),.Q(s_r_zeros[0:0]),.QN(n238));
  DFFX1 desc1016(.D(N3078),.CLK(clk_i),.Q(s_expo1[7:7]));
  DFFX1 desc1017(.D(N3077),.CLK(clk_i),.Q(s_expo1[6:6]));
  DFFX1 desc1018(.D(N3076),.CLK(clk_i),.Q(s_expo1[5:5]));
  DFFX1 desc1019(.D(N3075),.CLK(clk_i),.Q(s_expo1[4:4]));
  DFFX1 desc1020(.D(N3074),.CLK(clk_i),.Q(s_expo1[3:3]));
  DFFX1 desc1021(.D(N3073),.CLK(clk_i),.Q(s_expo1[2:2]));
  DFFX1 desc1022(.D(N3072),.CLK(clk_i),.Q(s_expo1[1:1]));
  DFFSSRX1 desc1023(.D(s_exp_10b[0:0]),.RSTB(1'b1),.SETB(n318),.CLK(clk_i),.Q(s_expo1[0:0]));
  DFFX1 desc1024(.D(N3086),.CLK(clk_i),.Q(s_shr2[5:5]));
  DFFX1 desc1025(.D(N3085),.CLK(clk_i),.Q(s_shr2[4:4]),.QN(n79));
  DFFX1 desc1026(.D(N3084),.CLK(clk_i),.Q(s_shr2[3:3]),.QN(n77));
  DFFX1 desc1027(.D(N3082),.CLK(clk_i),.Q(s_shr2[1:1]),.QN(n73));
  DFFX1 desc1028(.D(N3081),.CLK(clk_i),.Q(s_shr2[0:0]),.QN(n72));
  DFFX1 desc1029(.D(N3070),.CLK(clk_i),.Q(s_shl2[5:5]));
  DFFX1 desc1030(.D(N3069),.CLK(clk_i),.Q(s_shl2[4:4]));
  DFFX1 desc1031(.D(N3068),.CLK(clk_i),.Q(s_shl2[3:3]));
  DFFX1 desc1032(.D(N3067),.CLK(clk_i),.Q(s_shl2[2:2]),.QN(n56));
  DFFX1 desc1033(.D(N3066),.CLK(clk_i),.Q(s_shl2[1:1]),.QN(n53));
  DFFX1 desc1034(.D(N3065),.CLK(clk_i),.Q(n55),.QN(n76));
  DFFX1 desc1035(.D(N3236),.CLK(clk_i),.Q(s_frac2a[47:47]));
  DFFX1 desc1036(.D(N3235),.CLK(clk_i),.Q(s_frac2a[46:46]));
  DFFX1 desc1037(.D(N3234),.CLK(clk_i),.Q(s_frac2a[45:45]));
  DFFX1 desc1038(.D(N3233),.CLK(clk_i),.Q(s_frac2a[44:44]));
  DFFX1 desc1039(.D(N3232),.CLK(clk_i),.Q(s_frac2a[43:43]));
  DFFX1 desc1040(.D(N3231),.CLK(clk_i),.Q(s_frac2a[42:42]));
  DFFX1 desc1041(.D(N3230),.CLK(clk_i),.Q(s_frac2a[41:41]));
  DFFX1 desc1042(.D(N3229),.CLK(clk_i),.Q(s_frac2a[40:40]));
  DFFX1 desc1043(.D(N3228),.CLK(clk_i),.Q(s_frac2a[39:39]));
  DFFX1 desc1044(.D(N3227),.CLK(clk_i),.Q(s_frac2a[38:38]));
  DFFX1 desc1045(.D(N3226),.CLK(clk_i),.Q(s_frac2a[37:37]));
  DFFX1 desc1046(.D(N3225),.CLK(clk_i),.Q(s_frac2a[36:36]));
  DFFX1 desc1047(.D(N3224),.CLK(clk_i),.Q(s_frac2a[35:35]));
  DFFX1 desc1048(.D(N3223),.CLK(clk_i),.Q(s_frac2a[34:34]));
  DFFX1 desc1049(.D(N3222),.CLK(clk_i),.Q(s_frac2a[33:33]));
  DFFX1 desc1050(.D(N3221),.CLK(clk_i),.Q(s_frac2a[32:32]));
  DFFX1 desc1051(.D(N3220),.CLK(clk_i),.Q(s_frac2a[31:31]));
  DFFX1 desc1052(.D(N3219),.CLK(clk_i),.Q(s_frac2a[30:30]));
  DFFX1 desc1053(.D(N3218),.CLK(clk_i),.Q(s_frac2a[29:29]));
  DFFX1 desc1054(.D(N3217),.CLK(clk_i),.Q(s_frac2a[28:28]));
  DFFX1 desc1055(.D(N3216),.CLK(clk_i),.Q(s_frac2a[27:27]));
  DFFX1 desc1056(.D(N3215),.CLK(clk_i),.Q(s_frac2a[26:26]));
  DFFX1 desc1057(.D(N3214),.CLK(clk_i),.Q(s_frac2a[25:25]));
  DFFX1 desc1058(.D(N3213),.CLK(clk_i),.Q(s_frac2a[24:24]));
  DFFX1 desc1059(.D(N3212),.CLK(clk_i),.Q(s_frac2a[23:23]));
  DFFX1 desc1060(.D(N3211),.CLK(clk_i),.Q(s_frac2a[22:22]));
  DFFX1 desc1061(.D(N3210),.CLK(clk_i),.Q(s_frac2a[21:21]));
  DFFX1 desc1062(.D(N3209),.CLK(clk_i),.Q(s_frac2a[20:20]));
  DFFX1 desc1063(.D(N3208),.CLK(clk_i),.QN(n1151));
  DFFX1 desc1064(.D(N3207),.CLK(clk_i),.QN(n1144));
  DFFX1 desc1065(.D(N3206),.CLK(clk_i),.QN(n1145));
  DFFX1 desc1066(.D(N3205),.CLK(clk_i),.QN(n1146));
  DFFX1 desc1067(.D(N3204),.CLK(clk_i),.Q(s_frac2a[15:15]));
  DFFX1 desc1068(.D(N3203),.CLK(clk_i),.Q(s_frac2a[14:14]));
  DFFX1 desc1069(.D(N3202),.CLK(clk_i),.Q(s_frac2a[13:13]));
  DFFX1 desc1070(.D(N3201),.CLK(clk_i),.QN(n1202));
  DFFX1 desc1071(.D(N3200),.CLK(clk_i),.QN(n1203));
  DFFX1 desc1072(.D(N3199),.CLK(clk_i),.QN(n1201));
  DFFX1 desc1073(.D(N3198),.CLK(clk_i),.QN(n1147));
  DFFX1 desc1074(.D(N3197),.CLK(clk_i),.QN(n1148));
  DFFX1 desc1075(.D(N3196),.CLK(clk_i),.QN(n1149));
  DFFX1 desc1076(.D(N3195),.CLK(clk_i),.Q(s_frac2a[6:6]));
  DFFX1 desc1077(.D(N3194),.CLK(clk_i),.Q(s_frac2a[5:5]));
  DFFX1 desc1078(.D(N3193),.CLK(clk_i),.Q(s_frac2a[4:4]));
  DFFX1 desc1079(.D(N3192),.CLK(clk_i),.Q(s_frac2a[3:3]));
  DFFX1 desc1080(.D(N3191),.CLK(clk_i),.Q(s_frac2a[2:2]));
  DFFX1 desc1081(.D(N3190),.CLK(clk_i),.QN(n1150));
  DFFX1 desc1082(.D(N3189),.CLK(clk_i),.Q(s_frac2a[0:0]));
  DFFX1 desc1083(.D(N3327),.CLK(clk_i),.Q(s_frac_rnd[24:24]),.QN(n244));
  DFFX1 ine_o_reg(.D(N3532),.CLK(clk_i),.Q(ine_o));
  DFFX1 desc1084(.D(s_output_o[30:30]),.CLK(clk_i),.Q(output_o[30:30]));
  DFFX1 desc1085(.D(s_output_o[29:29]),.CLK(clk_i),.Q(output_o[29:29]));
  DFFX1 desc1086(.D(s_output_o[28:28]),.CLK(clk_i),.Q(output_o[28:28]));
  DFFX1 desc1087(.D(s_output_o[27:27]),.CLK(clk_i),.Q(output_o[27:27]));
  DFFX1 desc1088(.D(s_output_o[26:26]),.CLK(clk_i),.Q(output_o[26:26]));
  DFFX1 desc1089(.D(s_output_o[25:25]),.CLK(clk_i),.Q(output_o[25:25]));
  DFFX1 desc1090(.D(s_output_o[24:24]),.CLK(clk_i),.Q(output_o[24:24]));
  DFFX1 desc1091(.D(s_output_o[23:23]),.CLK(clk_i),.Q(output_o[23:23]));
  DFFX1 desc1092(.D(N3326),.CLK(clk_i),.Q(s_frac_rnd[23:23]));
  DFFX1 desc1093(.D(N3325),.CLK(clk_i),.Q(s_frac_rnd[22:22]));
  DFFX1 desc1094(.D(s_output_o[22:22]),.CLK(clk_i),.Q(output_o[22:22]));
  DFFX1 desc1095(.D(N3324),.CLK(clk_i),.Q(s_frac_rnd[21:21]));
  DFFX1 desc1096(.D(s_output_o[21:21]),.CLK(clk_i),.Q(output_o[21:21]));
  DFFX1 desc1097(.D(N3323),.CLK(clk_i),.Q(s_frac_rnd[20:20]));
  DFFX1 desc1098(.D(s_output_o[20:20]),.CLK(clk_i),.Q(output_o[20:20]));
  DFFX1 desc1099(.D(N3322),.CLK(clk_i),.Q(s_frac_rnd[19:19]));
  DFFX1 desc1100(.D(s_output_o[19:19]),.CLK(clk_i),.Q(output_o[19:19]));
  DFFX1 desc1101(.D(N3321),.CLK(clk_i),.Q(s_frac_rnd[18:18]));
  DFFX1 desc1102(.D(s_output_o[18:18]),.CLK(clk_i),.Q(output_o[18:18]));
  DFFX1 desc1103(.D(N3320),.CLK(clk_i),.Q(s_frac_rnd[17:17]));
  DFFX1 desc1104(.D(s_output_o[17:17]),.CLK(clk_i),.Q(output_o[17:17]));
  DFFX1 desc1105(.D(N3319),.CLK(clk_i),.Q(s_frac_rnd[16:16]));
  DFFX1 desc1106(.D(s_output_o[16:16]),.CLK(clk_i),.Q(output_o[16:16]));
  DFFX1 desc1107(.D(N3318),.CLK(clk_i),.Q(s_frac_rnd[15:15]));
  DFFX1 desc1108(.D(s_output_o[15:15]),.CLK(clk_i),.Q(output_o[15:15]));
  DFFX1 desc1109(.D(N3317),.CLK(clk_i),.Q(s_frac_rnd[14:14]));
  DFFX1 desc1110(.D(s_output_o[14:14]),.CLK(clk_i),.Q(output_o[14:14]));
  DFFX1 desc1111(.D(N3316),.CLK(clk_i),.Q(s_frac_rnd[13:13]));
  DFFX1 desc1112(.D(s_output_o[13:13]),.CLK(clk_i),.Q(output_o[13:13]));
  DFFX1 desc1113(.D(N3315),.CLK(clk_i),.Q(s_frac_rnd[12:12]));
  DFFX1 desc1114(.D(s_output_o[12:12]),.CLK(clk_i),.Q(output_o[12:12]));
  DFFX1 desc1115(.D(N3314),.CLK(clk_i),.Q(s_frac_rnd[11:11]));
  DFFX1 desc1116(.D(s_output_o[11:11]),.CLK(clk_i),.Q(output_o[11:11]));
  DFFX1 desc1117(.D(N3313),.CLK(clk_i),.Q(s_frac_rnd[10:10]));
  DFFX1 desc1118(.D(s_output_o[10:10]),.CLK(clk_i),.Q(output_o[10:10]));
  DFFX1 desc1119(.D(N3312),.CLK(clk_i),.Q(s_frac_rnd[9:9]));
  DFFX1 desc1120(.D(s_output_o[9:9]),.CLK(clk_i),.Q(output_o[9:9]));
  DFFX1 desc1121(.D(N3311),.CLK(clk_i),.Q(s_frac_rnd[8:8]));
  DFFX1 desc1122(.D(s_output_o[8:8]),.CLK(clk_i),.Q(output_o[8:8]));
  DFFX1 desc1123(.D(N3310),.CLK(clk_i),.Q(s_frac_rnd[7:7]));
  DFFX1 desc1124(.D(s_output_o[7:7]),.CLK(clk_i),.Q(output_o[7:7]));
  DFFX1 desc1125(.D(N3309),.CLK(clk_i),.Q(s_frac_rnd[6:6]));
  DFFX1 desc1126(.D(s_output_o[6:6]),.CLK(clk_i),.Q(output_o[6:6]));
  DFFX1 desc1127(.D(N3308),.CLK(clk_i),.Q(s_frac_rnd[5:5]));
  DFFX1 desc1128(.D(s_output_o[5:5]),.CLK(clk_i),.Q(output_o[5:5]));
  DFFX1 desc1129(.D(N3307),.CLK(clk_i),.Q(s_frac_rnd[4:4]));
  DFFX1 desc1130(.D(s_output_o[4:4]),.CLK(clk_i),.Q(output_o[4:4]));
  DFFX1 desc1131(.D(N3306),.CLK(clk_i),.Q(s_frac_rnd[3:3]));
  DFFX1 desc1132(.D(s_output_o[3:3]),.CLK(clk_i),.Q(output_o[3:3]));
  DFFX1 desc1133(.D(N3305),.CLK(clk_i),.Q(s_frac_rnd[2:2]));
  DFFX1 desc1134(.D(s_output_o[2:2]),.CLK(clk_i),.Q(output_o[2:2]));
  DFFX1 desc1135(.D(N3304),.CLK(clk_i),.Q(s_frac_rnd[1:1]));
  DFFX1 desc1136(.D(s_output_o[1:1]),.CLK(clk_i),.Q(output_o[1:1]));
  DFFX1 desc1137(.D(N3303),.CLK(clk_i),.Q(s_frac_rnd[0:0]));
  DFFX1 desc1138(.D(s_output_o[0:0]),.CLK(clk_i),.Q(output_o[0:0]));
  AO22X1 U344(.IN1(s_frac_rnd[10:10]),.IN2(n246),.IN3(s_frac_rnd[9:9]),.IN4(n1218),.Q(s_output_o[9:9]));
  AO22X1 U345(.IN1(n246),.IN2(s_frac_rnd[9:9]),.IN3(s_frac_rnd[8:8]),.IN4(n247),.Q(s_output_o[8:8]));
  AO22X1 U346(.IN1(s_frac_rnd[8:8]),.IN2(n246),.IN3(s_frac_rnd[7:7]),.IN4(n1219),.Q(s_output_o[7:7]));
  AO22X1 U347(.IN1(s_frac_rnd[7:7]),.IN2(n246),.IN3(s_frac_rnd[6:6]),.IN4(n1218),.Q(s_output_o[6:6]));
  AO22X1 U348(.IN1(s_frac_rnd[6:6]),.IN2(n246),.IN3(s_frac_rnd[5:5]),.IN4(n247),.Q(s_output_o[5:5]));
  AO22X1 U349(.IN1(s_frac_rnd[5:5]),.IN2(n246),.IN3(s_frac_rnd[4:4]),.IN4(n1219),.Q(s_output_o[4:4]));
  AO22X1 U350(.IN1(s_frac_rnd[4:4]),.IN2(n246),.IN3(s_frac_rnd[3:3]),.IN4(n1218),.Q(s_output_o[3:3]));
  AO221X1 U351(.IN1(n248),.IN2(s_expo2b[7:7]),.IN3(n249),.IN4(N3353),.IN5(n250),.Q(s_output_o[30:30]));
  AO22X1 U352(.IN1(s_frac_rnd[3:3]),.IN2(n246),.IN3(s_frac_rnd[2:2]),.IN4(n247),.Q(s_output_o[2:2]));
  AO221X1 U353(.IN1(n248),.IN2(s_expo2b[6:6]),.IN3(n249),.IN4(N3352),.IN5(n250),.Q(s_output_o[29:29]));
  AO221X1 U354(.IN1(n248),.IN2(s_expo2b[5:5]),.IN3(n249),.IN4(N3351),.IN5(n250),.Q(s_output_o[28:28]));
  AO221X1 U355(.IN1(n248),.IN2(s_expo2b[4:4]),.IN3(n249),.IN4(N3350),.IN5(n250),.Q(s_output_o[27:27]));
  AO221X1 U356(.IN1(n248),.IN2(s_expo2b[3:3]),.IN3(n249),.IN4(N3349),.IN5(n250),.Q(s_output_o[26:26]));
  AO221X1 U357(.IN1(n248),.IN2(s_expo2b[2:2]),.IN3(n249),.IN4(N3348),.IN5(n250),.Q(s_output_o[25:25]));
  AO221X1 U358(.IN1(n248),.IN2(s_expo2b[1:1]),.IN3(n249),.IN4(N3347),.IN5(n250),.Q(s_output_o[24:24]));
  AO221X1 U359(.IN1(n248),.IN2(s_expo2b[0:0]),.IN3(n249),.IN4(N3346),.IN5(n250),.Q(s_output_o[23:23]));
  OAI221X1 U360(.IN1(n1335),.IN2(n251),.IN3(n1334),.IN4(n252),.IN5(n253),.QN(s_output_o[22:22]));
  NAND4X0 U361(.IN1(n1335),.IN2(n256),.IN3(n257),.IN4(n258),.QN(n255));
  AO22X1 U362(.IN1(s_frac_rnd[23:23]),.IN2(s_frac_rnd[24:24]),.IN3(s_frac_rnd[22:22]),.IN4(n244),.Q(n256));
  AO22X1 U363(.IN1(s_frac_rnd[22:22]),.IN2(n246),.IN3(s_frac_rnd[21:21]),.IN4(n1219),.Q(s_output_o[21:21]));
  AO22X1 U364(.IN1(s_frac_rnd[21:21]),.IN2(n246),.IN3(s_frac_rnd[20:20]),.IN4(n1218),.Q(s_output_o[20:20]));
  AO22X1 U365(.IN1(s_frac_rnd[2:2]),.IN2(n246),.IN3(s_frac_rnd[1:1]),.IN4(n247),.Q(s_output_o[1:1]));
  AO22X1 U366(.IN1(s_frac_rnd[20:20]),.IN2(n246),.IN3(s_frac_rnd[19:19]),.IN4(n1219),.Q(s_output_o[19:19]));
  AO22X1 U367(.IN1(s_frac_rnd[19:19]),.IN2(n246),.IN3(s_frac_rnd[18:18]),.IN4(n1218),.Q(s_output_o[18:18]));
  AO22X1 U368(.IN1(s_frac_rnd[18:18]),.IN2(n246),.IN3(s_frac_rnd[17:17]),.IN4(n247),.Q(s_output_o[17:17]));
  AO22X1 U369(.IN1(s_frac_rnd[17:17]),.IN2(n246),.IN3(s_frac_rnd[16:16]),.IN4(n1219),.Q(s_output_o[16:16]));
  AO22X1 U370(.IN1(s_frac_rnd[16:16]),.IN2(n246),.IN3(s_frac_rnd[15:15]),.IN4(n1218),.Q(s_output_o[15:15]));
  AO22X1 U371(.IN1(s_frac_rnd[15:15]),.IN2(n246),.IN3(s_frac_rnd[14:14]),.IN4(n247),.Q(s_output_o[14:14]));
  AO22X1 U372(.IN1(s_frac_rnd[14:14]),.IN2(n246),.IN3(s_frac_rnd[13:13]),.IN4(n1219),.Q(s_output_o[13:13]));
  AO22X1 U373(.IN1(s_frac_rnd[13:13]),.IN2(n246),.IN3(s_frac_rnd[12:12]),.IN4(n1218),.Q(s_output_o[12:12]));
  AO22X1 U374(.IN1(s_frac_rnd[12:12]),.IN2(n246),.IN3(s_frac_rnd[11:11]),.IN4(n247),.Q(s_output_o[11:11]));
  AO22X1 U375(.IN1(s_frac_rnd[11:11]),.IN2(n246),.IN3(s_frac_rnd[10:10]),.IN4(n1219),.Q(s_output_o[10:10]));
  AO22X1 U376(.IN1(s_frac_rnd[1:1]),.IN2(n246),.IN3(s_frac_rnd[0:0]),.IN4(n1218),.Q(s_output_o[0:0]));
  NAND4X0 U379(.IN1(s_r_zeros[4:4]),.IN2(n238),.IN3(s_r_zeros[5:5]),.IN4(n264),.QN(n257));
  NOR3X0 U380(.IN1(s_r_zeros[1:1]),.IN2(s_r_zeros[3:3]),.IN3(s_r_zeros[2:2]),.QN(n264));
  NOR3X0 U381(.IN1(n266),.IN2(n262),.IN3(n261),.QN(N3532));
  NOR4X0 U382(.IN1(s_opb_i[27:27]),.IN2(s_opb_i[26:26]),.IN3(n267),.IN4(n268),.QN(n261));
  OR4X1 U383(.IN1(s_opb_i[23:23]),.IN2(n260),.IN3(s_opb_i[25:25]),.IN4(s_opb_i[24:24]),.Q(n268));
  NAND4X0 U384(.IN1(n269),.IN2(n270),.IN3(n271),.IN4(n272),.QN(n260));
  NOR4X0 U385(.IN1(n273),.IN2(s_opb_i[4:4]),.IN3(s_opb_i[6:6]),.IN4(s_opb_i[5:5]),.QN(n272));
  NOR4X0 U387(.IN1(n274),.IN2(s_opb_i[1:1]),.IN3(s_opb_i[21:21]),.IN4(s_opb_i[20:20]),.QN(n271));
  NOR4X0 U389(.IN1(n275),.IN2(s_opb_i[14:14]),.IN3(s_opb_i[16:16]),.IN4(s_opb_i[15:15]),.QN(n270));
  NOR4X0 U391(.IN1(n276),.IN2(s_opb_i[11:11]),.IN3(s_opb_i[13:13]),.IN4(s_opb_i[12:12]),.QN(n269));
  NOR4X0 U394(.IN1(s_opa_i[27:27]),.IN2(s_opa_i[26:26]),.IN3(n277),.IN4(n278),.QN(n262));
  OR4X1 U395(.IN1(s_opa_i[23:23]),.IN2(n259),.IN3(s_opa_i[25:25]),.IN4(s_opa_i[24:24]),.Q(n278));
  NAND4X0 U396(.IN1(n279),.IN2(n280),.IN3(n281),.IN4(n282),.QN(n259));
  NOR4X0 U397(.IN1(n283),.IN2(s_opa_i[4:4]),.IN3(s_opa_i[6:6]),.IN4(s_opa_i[5:5]),.QN(n282));
  NOR4X0 U399(.IN1(n284),.IN2(s_opa_i[1:1]),.IN3(s_opa_i[21:21]),.IN4(s_opa_i[20:20]),.QN(n281));
  NOR4X0 U401(.IN1(n285),.IN2(s_opa_i[14:14]),.IN3(s_opa_i[16:16]),.IN4(s_opa_i[15:15]),.QN(n280));
  NOR4X0 U403(.IN1(n286),.IN2(s_opa_i[11:11]),.IN3(s_opa_i[13:13]),.IN4(s_opa_i[12:12]),.QN(n279));
  AND2X1 U406(.IN1(n258),.IN2(n287),.Q(n266));
  AO21X1 U407(.IN1(n288),.IN2(n289),.IN3(n265),.Q(n258));
  OR2X1 U408(.IN1(n290),.IN2(n291),.Q(n252));
  NAND4X0 U409(.IN1(s_expb[7:7]),.IN2(s_expb[6:6]),.IN3(s_expb[5:5]),.IN4(s_expb[4:4]),.QN(n291));
  NAND4X0 U410(.IN1(s_expb[3:3]),.IN2(s_expb[2:2]),.IN3(s_expb[1:1]),.IN4(s_expb[0:0]),.QN(n290));
  OR2X1 U411(.IN1(n292),.IN2(n293),.Q(n254));
  NAND4X0 U412(.IN1(s_expa[7:7]),.IN2(s_expa[6:6]),.IN3(s_expa[5:5]),.IN4(s_expa[4:4]),.QN(n293));
  NAND4X0 U413(.IN1(s_expa[3:3]),.IN2(s_expa[2:2]),.IN3(s_expa[1:1]),.IN4(s_expa[0:0]),.QN(n292));
  NAND4X0 U414(.IN1(s_expo2b[3:3]),.IN2(s_expo2b[2:2]),.IN3(n294),.IN4(n295),.QN(n289));
  AND4X1 U415(.IN1(s_expo2b[4:4]),.IN2(s_expo2b[5:5]),.IN3(s_expo2b[6:6]),.IN4(s_expo2b[7:7]),.Q(n295));
  AND3X1 U416(.IN1(s_expo2b[1:1]),.IN2(n1331),.IN3(s_expo2b[0:0]),.Q(n294));
  NAND4X0 U417(.IN1(s_frac_rnd[24:24]),.IN2(N3353),.IN3(n296),.IN4(n297),.QN(n288));
  NOR4X0 U418(.IN1(n298),.IN2(n1332),.IN3(N3354),.IN4(s_expo2b[0:0]),.QN(n297));
  AND3X1 U419(.IN1(N3351),.IN2(N3350),.IN3(N3352),.Q(n296));
  AO22X1 U420(.IN1(N3302),.IN2(n1257),.IN3(s_frac2a[47:47]),.IN4(n1256),.Q(N3327));
  AO22X1 U421(.IN1(N3301),.IN2(n1257),.IN3(n299),.IN4(s_frac2a[46:46]),.Q(N3326));
  AO22X1 U422(.IN1(N3300),.IN2(n1257),.IN3(s_frac2a[45:45]),.IN4(n1255),.Q(N3325));
  AO22X1 U423(.IN1(N3299),.IN2(n1257),.IN3(s_frac2a[44:44]),.IN4(n1255),.Q(N3324));
  AO22X1 U424(.IN1(N3298),.IN2(n1259),.IN3(s_frac2a[43:43]),.IN4(n1255),.Q(N3323));
  AO22X1 U425(.IN1(N3297),.IN2(n1258),.IN3(s_frac2a[42:42]),.IN4(n1255),.Q(N3322));
  AO22X1 U426(.IN1(N3296),.IN2(n1259),.IN3(s_frac2a[41:41]),.IN4(n1255),.Q(N3321));
  AO22X1 U427(.IN1(N3295),.IN2(n1258),.IN3(s_frac2a[40:40]),.IN4(n1255),.Q(N3320));
  AO22X1 U428(.IN1(N3294),.IN2(n1259),.IN3(s_frac2a[39:39]),.IN4(n1255),.Q(N3319));
  AO22X1 U429(.IN1(N3293),.IN2(n1258),.IN3(s_frac2a[38:38]),.IN4(n1255),.Q(N3318));
  AO22X1 U430(.IN1(N3292),.IN2(n1259),.IN3(s_frac2a[37:37]),.IN4(n1255),.Q(N3317));
  AO22X1 U431(.IN1(N3291),.IN2(n1258),.IN3(s_frac2a[36:36]),.IN4(n1255),.Q(N3316));
  AO22X1 U432(.IN1(N3290),.IN2(n1258),.IN3(s_frac2a[35:35]),.IN4(n1255),.Q(N3315));
  AO22X1 U433(.IN1(N3289),.IN2(n1258),.IN3(s_frac2a[34:34]),.IN4(n1256),.Q(N3314));
  AO22X1 U434(.IN1(N3288),.IN2(n1258),.IN3(s_frac2a[33:33]),.IN4(n1256),.Q(N3313));
  AO22X1 U435(.IN1(N3287),.IN2(n1258),.IN3(s_frac2a[32:32]),.IN4(n1256),.Q(N3312));
  AO22X1 U436(.IN1(N3286),.IN2(n1258),.IN3(s_frac2a[31:31]),.IN4(n1256),.Q(N3311));
  AO22X1 U437(.IN1(N3285),.IN2(n1258),.IN3(s_frac2a[30:30]),.IN4(n1256),.Q(N3310));
  AO22X1 U438(.IN1(N3284),.IN2(n1259),.IN3(s_frac2a[29:29]),.IN4(n1256),.Q(N3309));
  AO22X1 U439(.IN1(N3283),.IN2(n1259),.IN3(s_frac2a[28:28]),.IN4(n1256),.Q(N3308));
  AO22X1 U440(.IN1(N3282),.IN2(n1259),.IN3(s_frac2a[27:27]),.IN4(n1256),.Q(N3307));
  AO22X1 U441(.IN1(N3281),.IN2(n1259),.IN3(s_frac2a[26:26]),.IN4(n1256),.Q(N3306));
  AO22X1 U442(.IN1(N3280),.IN2(n1259),.IN3(s_frac2a[25:25]),.IN4(n1256),.Q(N3305));
  AO22X1 U443(.IN1(N3279),.IN2(n1259),.IN3(s_frac2a[24:24]),.IN4(n1256),.Q(N3304));
  AO22X1 U444(.IN1(N3278),.IN2(n1259),.IN3(s_frac2a[23:23]),.IN4(n1255),.Q(N3303));
  NAND4X0 U445(.IN1(s_frac2a[22:22]),.IN2(n302),.IN3(n236),.IN4(n235),.QN(n301));
  OR3X1 U446(.IN1(s_frac2a[21:21]),.IN2(s_frac2a[23:23]),.IN3(n303),.Q(n302));
  NAND3X0 U447(.IN1(\s_rmode_i[1] ),.IN2(n304),.IN3(s_output_o[31:31]),.QN(n305));
  NOR3X0 U448(.IN1(s_frac2a[21:21]),.IN2(s_frac2a[22:22]),.IN3(n303),.QN(n287));
  NAND4X0 U449(.IN1(n306),.IN2(n307),.IN3(n308),.IN4(n309),.QN(n303));
  NOR4X0 U450(.IN1(n310),.IN2(s_frac2a[4:4]),.IN3(s_frac2a[6:6]),.IN4(s_frac2a[5:5]),.QN(n309));
  NOR4X0 U452(.IN1(n311),.IN2(s_frac2a[20:20]),.IN3(s_frac2a[3:3]),.IN4(s_frac2a[2:2]),.QN(n308));
  NOR4X0 U454(.IN1(n312),.IN2(s_frac2a[13:13]),.IN3(s_frac2a[15:15]),.IN4(s_frac2a[14:14]),.QN(n307));
  AO22X1 U458(.IN1(N3140),.IN2(n1247),.IN3(N3188),.IN4(n1246),.Q(N3236));
  AO22X1 U459(.IN1(N3139),.IN2(n1247),.IN3(N3187),.IN4(n1246),.Q(N3235));
  AO22X1 U460(.IN1(N3138),.IN2(n1247),.IN3(N3186),.IN4(n1246),.Q(N3234));
  AO22X1 U461(.IN1(N3137),.IN2(n1248),.IN3(N3185),.IN4(n1246),.Q(N3233));
  AO22X1 U462(.IN1(N3136),.IN2(n1248),.IN3(n1391),.IN4(n1246),.Q(N3232));
  AO22X1 U463(.IN1(N3135),.IN2(n1248),.IN3(n1395),.IN4(n1246),.Q(N3231));
  AO22X1 U464(.IN1(N3134),.IN2(n1248),.IN3(n1400),.IN4(n1246),.Q(N3230));
  AO22X1 U465(.IN1(N3133),.IN2(n1248),.IN3(n1407),.IN4(n1246),.Q(N3229));
  AO22X1 U466(.IN1(N3132),.IN2(n1248),.IN3(n1412),.IN4(n1246),.Q(N3228));
  AO22X1 U467(.IN1(N3131),.IN2(n1248),.IN3(n1416),.IN4(n1246),.Q(N3227));
  AO22X1 U468(.IN1(N3130),.IN2(n1249),.IN3(n1420),.IN4(n1246),.Q(N3226));
  AO22X1 U469(.IN1(N3129),.IN2(n1249),.IN3(n1424),.IN4(n1246),.Q(N3225));
  AO22X1 U470(.IN1(N3128),.IN2(n1249),.IN3(n1433),.IN4(n1245),.Q(N3224));
  AO22X1 U471(.IN1(N3127),.IN2(n1249),.IN3(n1437),.IN4(n1245),.Q(N3223));
  AO22X1 U472(.IN1(N3126),.IN2(n1249),.IN3(n1441),.IN4(n1245),.Q(N3222));
  AO22X1 U473(.IN1(N3125),.IN2(n1249),.IN3(n1445),.IN4(n1245),.Q(N3221));
  AO22X1 U474(.IN1(N3124),.IN2(n1249),.IN3(N3172),.IN4(n1245),.Q(N3220));
  AO22X1 U475(.IN1(N3123),.IN2(n1250),.IN3(N3171),.IN4(n1245),.Q(N3219));
  AO22X1 U476(.IN1(N3122),.IN2(n1250),.IN3(N3170),.IN4(n1245),.Q(N3218));
  AO22X1 U477(.IN1(N3121),.IN2(n1250),.IN3(N3169),.IN4(n1245),.Q(N3217));
  AO22X1 U478(.IN1(N3120),.IN2(n1250),.IN3(N3168),.IN4(n1245),.Q(N3216));
  AO22X1 U479(.IN1(N3119),.IN2(n1250),.IN3(N3167),.IN4(n1245),.Q(N3215));
  AO22X1 U480(.IN1(N3118),.IN2(n1250),.IN3(N3166),.IN4(n1245),.Q(N3214));
  AO22X1 U481(.IN1(N3117),.IN2(n1250),.IN3(N3165),.IN4(n1245),.Q(N3213));
  AO22X1 U482(.IN1(N3116),.IN2(n1251),.IN3(N3164),.IN4(n1244),.Q(N3212));
  AO22X1 U483(.IN1(N3115),.IN2(n1251),.IN3(N3163),.IN4(n1244),.Q(N3211));
  AO22X1 U484(.IN1(N3114),.IN2(n1251),.IN3(N3162),.IN4(n1244),.Q(N3210));
  AO22X1 U485(.IN1(N3113),.IN2(n1251),.IN3(N3161),.IN4(n1244),.Q(N3209));
  AO22X1 U486(.IN1(N3112),.IN2(n1251),.IN3(N3160),.IN4(n1244),.Q(N3208));
  AO22X1 U487(.IN1(N3111),.IN2(n1251),.IN3(N3159),.IN4(n1244),.Q(N3207));
  AO22X1 U488(.IN1(N3110),.IN2(n1251),.IN3(N3158),.IN4(n1244),.Q(N3206));
  AO22X1 U489(.IN1(N3109),.IN2(n1252),.IN3(N3157),.IN4(n1244),.Q(N3205));
  AO22X1 U490(.IN1(N3108),.IN2(n1252),.IN3(N3156),.IN4(n1244),.Q(N3204));
  AO22X1 U491(.IN1(N3107),.IN2(n1252),.IN3(N3155),.IN4(n1244),.Q(N3203));
  AO22X1 U492(.IN1(N3106),.IN2(n1252),.IN3(N3154),.IN4(n1244),.Q(N3202));
  AO22X1 U493(.IN1(N3105),.IN2(n1252),.IN3(N3153),.IN4(n1244),.Q(N3201));
  AO22X1 U494(.IN1(N3104),.IN2(n1252),.IN3(N3152),.IN4(n1243),.Q(N3200));
  AO22X1 U495(.IN1(N3103),.IN2(n1252),.IN3(N3151),.IN4(n1243),.Q(N3199));
  AO22X1 U496(.IN1(N3102),.IN2(n1253),.IN3(N3150),.IN4(n1243),.Q(N3198));
  AO22X1 U497(.IN1(N3101),.IN2(n1253),.IN3(N3149),.IN4(n1243),.Q(N3197));
  AO22X1 U498(.IN1(N3100),.IN2(n1253),.IN3(N3148),.IN4(n1243),.Q(N3196));
  AO22X1 U499(.IN1(N3099),.IN2(n1253),.IN3(N3147),.IN4(n1243),.Q(N3195));
  AO22X1 U500(.IN1(N3098),.IN2(n1253),.IN3(N3146),.IN4(n1243),.Q(N3194));
  AO22X1 U501(.IN1(N3097),.IN2(n1253),.IN3(N3145),.IN4(n1243),.Q(N3193));
  AO22X1 U502(.IN1(N3096),.IN2(n1253),.IN3(N3144),.IN4(n1243),.Q(N3192));
  AO22X1 U503(.IN1(N3095),.IN2(n1254),.IN3(N3143),.IN4(n1243),.Q(N3191));
  AO22X1 U504(.IN1(N3094),.IN2(n1254),.IN3(N3142),.IN4(n1243),.Q(N3190));
  AO22X1 U505(.IN1(N3093),.IN2(n1254),.IN3(N3141),.IN4(n1243),.Q(N3189));
  OR3X1 U507(.IN1(n1286),.IN2(n1280),.IN3(s_shr2[3:3]),.Q(n315));
  AO21X1 U508(.IN1(N3004),.IN2(n316),.IN3(n317),.Q(N3086));
  AO21X1 U509(.IN1(N3003),.IN2(n316),.IN3(n317),.Q(N3085));
  AO21X1 U510(.IN1(N3002),.IN2(n316),.IN3(n317),.Q(N3084));
  AO21X1 U511(.IN1(N3001),.IN2(n316),.IN3(n317),.Q(N3083));
  AO21X1 U512(.IN1(N3000),.IN2(n316),.IN3(n317),.Q(N3082));
  AO221X1 U513(.IN1(N2993),.IN2(n318),.IN3(N2999),.IN4(n316),.IN5(n317),.Q(N3081));
  AND2X1 U514(.IN1(N3005),.IN2(n316),.Q(n317));
  AO21X1 U515(.IN1(s_exp_10b[7:7]),.IN2(n319),.IN3(n320),.Q(N3078));
  AO21X1 U516(.IN1(s_exp_10b[6:6]),.IN2(n319),.IN3(n320),.Q(N3077));
  AO21X1 U517(.IN1(s_exp_10b[5:5]),.IN2(n319),.IN3(n320),.Q(N3076));
  AO21X1 U518(.IN1(s_exp_10b[4:4]),.IN2(n319),.IN3(n320),.Q(N3075));
  AO21X1 U519(.IN1(s_exp_10b[3:3]),.IN2(n319),.IN3(n320),.Q(N3074));
  AO21X1 U520(.IN1(s_exp_10b[2:2]),.IN2(n319),.IN3(n320),.Q(N3073));
  AO21X1 U521(.IN1(s_exp_10b[1:1]),.IN2(n319),.IN3(n320),.Q(N3072));
  AND2X1 U522(.IN1(s_exp_10b[8:8]),.IN2(n319),.Q(n320));
  AO22X1 U523(.IN1(s_zeros[5:5]),.IN2(n318),.IN3(N3024),.IN4(n321),.Q(N3070));
  AO22X1 U524(.IN1(s_zeros[4:4]),.IN2(n318),.IN3(N3023),.IN4(n321),.Q(N3069));
  AO22X1 U525(.IN1(s_zeros[3:3]),.IN2(n318),.IN3(N3022),.IN4(n321),.Q(N3068));
  AO22X1 U526(.IN1(s_zeros[2:2]),.IN2(n318),.IN3(N3021),.IN4(n321),.Q(N3067));
  AO22X1 U527(.IN1(s_zeros[1:1]),.IN2(n318),.IN3(N3020),.IN4(n321),.Q(N3066));
  AO22X1 U528(.IN1(s_zeros[0:0]),.IN2(n318),.IN3(N3019),.IN4(n321),.Q(N3065));
  NOR4X0 U529(.IN1(n324),.IN2(n325),.IN3(s_exp_10b[5:5]),.IN4(s_exp_10b[4:4]),.QN(n323));
  OR3X1 U530(.IN1(s_exp_10b[7:7]),.IN2(s_exp_10b[8:8]),.IN3(s_exp_10b[6:6]),.Q(n325));
  OR4X1 U531(.IN1(s_exp_10b[0:0]),.IN2(s_exp_10b[1:1]),.IN3(s_exp_10b[2:2]),.IN4(s_exp_10b[3:3]),.Q(n324));
  NOR4X0 U533(.IN1(n328),.IN2(s_exp_10a[6:6]),.IN3(s_exp_10a[8:8]),.IN4(s_exp_10a[7:7]),.QN(n327));
  OR2X1 U534(.IN1(s_exp_10a[5:5]),.IN2(s_exp_10a[4:4]),.Q(n328));
  NOR4X0 U535(.IN1(s_exp_10a[3:3]),.IN2(s_exp_10a[2:2]),.IN3(s_exp_10a[1:1]),.IN4(s_exp_10a[0:0]),.QN(n326));
  AOI222X1 U540(.IN1(n1010),.IN2(n343),.IN3(n594),.IN4(n1210),.IN5(n913),.IN6(n344),.QN(n342));
  AOI22X1 U541(.IN1(n919),.IN2(n345),.IN3(N1873),.IN4(n346),.QN(n341));
  AO21X1 U542(.IN1(n348),.IN2(n349),.IN3(n1486),.Q(n339));
  AO22X1 U547(.IN1(n362),.IN2(n1052),.IN3(n363),.IN4(n995),.Q(n361));
  NAND4X0 U548(.IN1(n364),.IN2(n365),.IN3(n366),.IN4(n367),.QN(n360));
  AOI222X1 U549(.IN1(N2129),.IN2(n368),.IN3(n1080),.IN4(n1216),.IN5(n1065),.IN6(n369),.QN(n367));
  AOI22X1 U550(.IN1(n1016),.IN2(n370),.IN3(n1061),.IN4(n371),.QN(n366));
  OA22X1 U553(.IN1(n1321),.IN2(n379),.IN3(n1320),.IN4(n380),.Q(n378));
  AOI222X1 U557(.IN1(N1937),.IN2(n389),.IN3(n999),.IN4(n1213),.IN5(n1029),.IN6(n390),.QN(n348));
  AO221X1 U558(.IN1(n334),.IN2(n176),.IN3(n1222),.IN4(N1696),.IN5(n393),.Q(n392));
  AO22X1 U559(.IN1(n332),.IN2(n945),.IN3(n333),.IN4(n898),.Q(n393));
  AO221X1 U560(.IN1(n1501),.IN2(n1040),.IN3(n394),.IN4(n1500),.IN5(n395),.Q(n391));
  AO22X1 U561(.IN1(n337),.IN2(n951),.IN3(n338),.IN4(n912),.Q(n395));
  NAND4X0 U562(.IN1(n396),.IN2(n397),.IN3(n398),.IN4(n399),.QN(n394));
  AOI222X1 U563(.IN1(n207),.IN2(n343),.IN3(n1092),.IN4(n1211),.IN5(n891),.IN6(n344),.QN(n399));
  AO21X1 U565(.IN1(n400),.IN2(n401),.IN3(n1486),.Q(n396));
  OA221X1 U566(.IN1(n351),.IN2(n402),.IN3(n1326),.IN4(n352),.IN5(n403),.Q(n401));
  OA22X1 U567(.IN1(n1328),.IN2(n354),.IN3(n1327),.IN4(n355),.Q(n403));
  AO22X1 U570(.IN1(n362),.IN2(n807),.IN3(n363),.IN4(n645),.Q(n407));
  NAND4X0 U571(.IN1(n408),.IN2(n409),.IN3(n410),.IN4(n411),.QN(n406));
  AO21X1 U574(.IN1(n412),.IN2(n413),.IN3(n1435),.Q(n408));
  OA221X1 U575(.IN1(n414),.IN2(n376),.IN3(n1034),.IN4(n377),.IN5(n415),.Q(n413));
  OA22X1 U576(.IN1(n1325),.IN2(n379),.IN3(n1324),.IN4(n380),.Q(n415));
  AOI222X1 U580(.IN1(n175),.IN2(n389),.IN3(n996),.IN4(n1214),.IN5(n26),.IN6(n390),.QN(n400));
  AO221X1 U581(.IN1(n334),.IN2(n927),.IN3(n1222),.IN4(n1013),.IN5(n420),.Q(n419));
  AO22X1 U582(.IN1(n332),.IN2(n939),.IN3(n333),.IN4(n61),.Q(n420));
  AO221X1 U583(.IN1(n1501),.IN2(n1014),.IN3(n421),.IN4(n1500),.IN5(n422),.Q(n418));
  AO22X1 U584(.IN1(n337),.IN2(n203),.IN3(n338),.IN4(n1102),.Q(n422));
  NAND4X0 U585(.IN1(n423),.IN2(n424),.IN3(n425),.IN4(n426),.QN(n421));
  AOI222X1 U586(.IN1(n924),.IN2(n343),.IN3(n1142),.IN4(n1210),.IN5(n810),.IN6(n344),.QN(n426));
  AOI22X1 U587(.IN1(n28),.IN2(n345),.IN3(n1140),.IN4(n346),.QN(n425));
  AO21X1 U588(.IN1(n427),.IN2(n428),.IN3(n1486),.Q(n423));
  OA221X1 U589(.IN1(n430),.IN2(n351),.IN3(n1467),.IN4(n352),.IN5(n431),.Q(n428));
  OA22X1 U590(.IN1(n1474),.IN2(n354),.IN3(n1469),.IN4(n355),.Q(n431));
  AO22X1 U593(.IN1(n362),.IN2(n1086),.IN3(n363),.IN4(n185),.Q(n435));
  NAND4X0 U594(.IN1(n436),.IN2(n437),.IN3(n438),.IN4(n439),.QN(n434));
  AO21X1 U597(.IN1(n440),.IN2(n441),.IN3(n1435),.Q(n436));
  OA221X1 U598(.IN1(n376),.IN2(n443),.IN3(n959),.IN4(n377),.IN5(n444),.Q(n441));
  OA22X1 U599(.IN1(n1409),.IN2(n379),.IN3(n1402),.IN4(n380),.Q(n444));
  OA22X1 U606(.IN1(n1502),.IN2(n450),.IN3(n457),.IN4(n449),.Q(n456));
  AO22X1 U609(.IN1(n346),.IN2(n1049),.IN3(n345),.IN4(n149),.Q(n461));
  NAND4X0 U610(.IN1(n462),.IN2(n463),.IN3(n464),.IN4(n465),.QN(n460));
  AOI222X1 U611(.IN1(n809),.IN2(n389),.IN3(n1050),.IN4(n1214),.IN5(n27),.IN6(n390),.QN(n465));
  OA22X1 U612(.IN1(n1475),.IN2(n354),.IN3(n1470),.IN4(n355),.Q(n464));
  AO21X1 U613(.IN1(n466),.IN2(n467),.IN3(n351),.Q(n462));
  OA221X1 U614(.IN1(n447),.IN2(n468),.IN3(n1455),.IN4(n448),.IN5(n469),.Q(n467));
  AOI22X1 U615(.IN1(n205),.IN2(n363),.IN3(N2062),.IN4(n362),.QN(n469));
  AO22X1 U618(.IN1(n371),.IN2(n960),.IN3(n370),.IN4(n877),.Q(n473));
  OA22X1 U621(.IN1(n1397),.IN2(n377),.IN3(n477),.IN4(n376),.Q(n475));
  OA22X1 U624(.IN1(n870),.IN2(n379),.IN3(n1403),.IN4(n380),.Q(n474));
  AOI22X1 U626(.IN1(n916),.IN2(n338),.IN3(n843),.IN4(n337),.QN(n455));
  AOI22X1 U627(.IN1(n1001),.IN2(n333),.IN3(n955),.IN4(n332),.QN(n454));
  AOI22X1 U628(.IN1(n230),.IN2(n334),.IN3(n163),.IN4(n1222),.QN(n453));
  AO22X1 U629(.IN1(n331),.IN2(n480),.IN3(n481),.IN4(n1134),.Q(N2975));
  NAND4X0 U630(.IN1(n482),.IN2(n483),.IN3(n484),.IN4(n485),.QN(n480));
  NAND4X0 U635(.IN1(n491),.IN2(n492),.IN3(n493),.IN4(n494),.QN(n489));
  OA22X1 U637(.IN1(n1476),.IN2(n354),.IN3(n1471),.IN4(n355),.Q(n493));
  AO21X1 U638(.IN1(n495),.IN2(n496),.IN3(n351),.Q(n491));
  OA221X1 U639(.IN1(n447),.IN2(n497),.IN3(n1456),.IN4(n448),.IN5(n498),.Q(n496));
  AOI22X1 U640(.IN1(n932),.IN2(n363),.IN3(N2061),.IN4(n362),.QN(n498));
  AO22X1 U643(.IN1(n371),.IN2(n829),.IN3(n370),.IN4(n973),.Q(n502));
  AOI222X1 U645(.IN1(n479),.IN2(n387),.IN3(n199),.IN4(s_fract_48_i[36:36]),.IN5(n846),.IN6(n388),.QN(n505));
  OA22X1 U646(.IN1(n181),.IN2(n377),.IN3(n506),.IN4(n376),.Q(n504));
  OA22X1 U649(.IN1(n1410),.IN2(n379),.IN3(n1404),.IN4(n380),.Q(n503));
  AOI222X1 U650(.IN1(n963),.IN2(n359),.IN3(n417),.IN4(n1289),.IN5(n985),.IN6(n358),.QN(n495));
  AOI22X1 U651(.IN1(n153),.IN2(n338),.IN3(n1091),.IN4(n337),.QN(n484));
  AOI22X1 U652(.IN1(n998),.IN2(n333),.IN3(n953),.IN4(n332),.QN(n483));
  AO22X1 U654(.IN1(n509),.IN2(n233),.IN3(n331),.IN4(n510),.Q(N2974));
  NAND4X0 U655(.IN1(n511),.IN2(n512),.IN3(n513),.IN4(n514),.QN(n510));
  OA22X1 U656(.IN1(N1798),.IN2(n450),.IN3(n515),.IN4(n449),.Q(n514));
  AO22X1 U659(.IN1(n346),.IN2(N1868),.IN3(n345),.IN4(N1852),.Q(n521));
  NAND4X0 U660(.IN1(n524),.IN2(n525),.IN3(n526),.IN4(n527),.QN(n520));
  AOI222X1 U661(.IN1(N1932),.IN2(n389),.IN3(N1900),.IN4(n1214),.IN5(N1916),.IN6(n390),.QN(n527));
  AND2X1 U662(.IN1(n528),.IN2(n204),.Q(n390));
  OA22X1 U663(.IN1(N1958),.IN2(n354),.IN3(n1472),.IN4(n355),.Q(n526));
  OR2X1 U664(.IN1(n530),.IN2(n531),.Q(n355));
  AO21X1 U665(.IN1(n532),.IN2(n533),.IN3(n351),.Q(n524));
  OA221X1 U666(.IN1(n534),.IN2(n447),.IN3(N2086),.IN4(n448),.IN5(n535),.Q(n533));
  AOI22X1 U667(.IN1(N2044),.IN2(n363),.IN3(N2060),.IN4(n362),.QN(n535));
  AND2X1 U668(.IN1(n538),.IN2(n536),.Q(n363));
  AO222X1 U669(.IN1(n369),.IN2(N2108),.IN3(n1216),.IN4(N2092),.IN5(n368),.IN6(N2124),.Q(n540));
  AO221X1 U670(.IN1(n372),.IN2(N2172),.IN3(n442),.IN4(n543),.IN5(n544),.Q(n539));
  AO22X1 U671(.IN1(n371),.IN2(N2156),.IN3(n370),.IN4(N2140),.Q(n544));
  NAND3X0 U672(.IN1(n547),.IN2(n548),.IN3(n549),.QN(n543));
  AOI222X1 U673(.IN1(N2220),.IN2(n387),.IN3(N2188),.IN4(s_fract_48_i[36:36]),.IN5(N2204),.IN6(n388),.QN(n549));
  AND2X1 U674(.IN1(n550),.IN2(n152),.Q(n388));
  OA22X1 U675(.IN1(N2278),.IN2(n377),.IN3(n552),.IN4(n376),.Q(n548));
  AO222X1 U676(.IN1(n383),.IN2(N2300),.IN3(n1231),.IN4(N2284),.IN5(n384),.IN6(N2316),.Q(n554));
  AND2X1 U677(.IN1(n555),.IN2(n556),.Q(n384));
  AO222X1 U678(.IN1(N2358),.IN2(n1336),.IN3(n385),.IN4(N2332),.IN5(n386),.IN6(N2348),.Q(n553));
  AND2X1 U679(.IN1(n557),.IN2(n558),.Q(n386));
  OA22X1 U681(.IN1(N2246),.IN2(n379),.IN3(N2262),.IN4(n380),.Q(n547));
  OR2X1 U682(.IN1(n560),.IN2(n559),.Q(n380));
  AOI222X1 U683(.IN1(N2028),.IN2(n359),.IN3(N1996),.IN4(n1289),.IN5(N2012),.IN6(n358),.QN(n532));
  AND2X1 U684(.IN1(n561),.IN2(n177),.Q(n358));
  AOI22X1 U685(.IN1(N1756),.IN2(n338),.IN3(N1772),.IN4(n337),.QN(n513));
  AND2X1 U686(.IN1(n564),.IN2(n563),.Q(n338));
  AOI22X1 U687(.IN1(N1708),.IN2(n333),.IN3(N1724),.IN4(n332),.QN(n512));
  AND2X1 U688(.IN1(n565),.IN2(n566),.Q(n332));
  AOI22X1 U689(.IN1(N1740),.IN2(n334),.IN3(N1692),.IN4(n1220),.QN(n511));
  AO21X1 U690(.IN1(n567),.IN2(n452),.IN3(n1137),.Q(n509));
  AND2X1 U691(.IN1(n481),.IN2(n1136),.Q(n567));
  AO22X1 U693(.IN1(N2346),.IN2(n69),.IN3(n1205),.IN4(n991),.Q(N2352));
  AO22X1 U694(.IN1(N2345),.IN2(n69),.IN3(n1205),.IN4(n11),.Q(N2351));
  AO22X1 U695(.IN1(N2344),.IN2(n69),.IN3(n1205),.IN4(n892),.Q(N2350));
  AO22X1 U696(.IN1(N2343),.IN2(n69),.IN3(n1205),.IN4(n42),.Q(N2349));
  AO22X1 U697(.IN1(n35),.IN2(n69),.IN3(n1205),.IN4(N2332),.Q(N2348));
  AO22X1 U703(.IN1(N2326),.IN2(n118),.IN3(s_fract_48_i[45:45]),.IN4(N2316),.Q(N2332));
  AO22X1 U708(.IN1(N2311),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n896),.Q(N2317));
  AO22X1 U715(.IN1(N2294),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(N2284),.Q(N2300));
  AO22X1 U717(.IN1(N2282),.IN2(n123),.IN3(n1229),.IN4(n1042),.Q(N2288));
  AO22X1 U719(.IN1(N2280),.IN2(n123),.IN3(n1231),.IN4(N2270),.Q(N2286));
  AO22X1 U721(.IN1(N2278),.IN2(n123),.IN3(n1231),.IN4(N2268),.Q(N2284));
  AO22X1 U727(.IN1(N2262),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(N2252),.Q(N2268));
  AO22X1 U733(.IN1(N2246),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N2236),.Q(N2252));
  AO22X1 U739(.IN1(N2230),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(N2220),.Q(N2236));
  AO22X1 U744(.IN1(N2215),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n846),.Q(N2221));
  AO22X1 U745(.IN1(N2214),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(N2204),.Q(N2220));
  AO22X1 U751(.IN1(N2198),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N2188),.Q(N2204));
  AO22X1 U756(.IN1(N2183),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n699),.Q(N2189));
  AO22X1 U757(.IN1(N2182),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(N2172),.Q(N2188));
  AO22X1 U762(.IN1(N2167),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n829),.Q(N2173));
  AO22X1 U763(.IN1(N2166),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(N2156),.Q(N2172));
  AO22X1 U765(.IN1(N2154),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n1125),.Q(N2160));
  AO22X1 U767(.IN1(N2152),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n877),.Q(N2158));
  AO22X1 U768(.IN1(N2151),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n973),.Q(N2157));
  AO22X1 U769(.IN1(N2150),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(N2140),.Q(N2156));
  AO22X1 U775(.IN1(N2134),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N2124),.Q(N2140));
  AO22X1 U781(.IN1(N2118),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(N2108),.Q(N2124));
  AO22X1 U786(.IN1(N2103),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n965),.Q(N2109));
  AO22X1 U787(.IN1(N2102),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(N2092),.Q(N2108));
  AO22X1 U789(.IN1(N2090),.IN2(n164),.IN3(n1217),.IN4(n33),.Q(N2096));
  AO22X1 U791(.IN1(N2088),.IN2(n164),.IN3(n1217),.IN4(n132),.Q(N2094));
  AO22X1 U792(.IN1(N2087),.IN2(n164),.IN3(n1216),.IN4(n915),.Q(N2093));
  AO22X1 U793(.IN1(N2086),.IN2(n164),.IN3(n1216),.IN4(N2076),.Q(N2092));
  AO22X1 U799(.IN1(N2070),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N2060),.Q(N2076));
  AO22X1 U805(.IN1(N2054),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(N2044),.Q(N2060));
  AO22X1 U810(.IN1(N2039),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n963),.Q(N2045));
  AO22X1 U811(.IN1(N2038),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(N2028),.Q(N2044));
  AO22X1 U816(.IN1(N2023),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n985),.Q(N2029));
  AO22X1 U817(.IN1(N2022),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(N2012),.Q(N2028));
  AO22X1 U823(.IN1(N2006),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(N1996),.Q(N2012));
  AO22X1 U827(.IN1(N1992),.IN2(n177),.IN3(n1290),.IN4(n683),.Q(N1998));
  AO22X1 U828(.IN1(N1991),.IN2(n177),.IN3(n1290),.IN4(n947),.Q(N1997));
  AO22X1 U829(.IN1(N1990),.IN2(n177),.IN3(n1290),.IN4(N1980),.Q(N1996));
  AO22X1 U834(.IN1(N1975),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1041),.Q(N1981));
  AO22X1 U835(.IN1(n1472),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(N1964),.Q(N1980));
  AO22X1 U836(.IN1(N1963),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N1953),.Q(N1969));
  AO22X1 U839(.IN1(N1960),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n188),.Q(N1966));
  AO22X1 U840(.IN1(N1959),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N1949),.Q(N1965));
  AO22X1 U841(.IN1(N1958),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N1948),.Q(N1964));
  AO22X1 U843(.IN1(N1946),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n175),.Q(N1952));
  AO22X1 U847(.IN1(N1942),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(N1932),.Q(N1948));
  AO22X1 U852(.IN1(N1927),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n885),.Q(N1933));
  AO22X1 U853(.IN1(N1926),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(N1916),.Q(N1932));
  AO22X1 U859(.IN1(N1910),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(N1900),.Q(N1916));
  AO22X1 U861(.IN1(n204),.IN2(N1898),.IN3(n1213),.IN4(n187),.Q(N1904));
  AO22X1 U863(.IN1(N1896),.IN2(n204),.IN3(n1213),.IN4(n887),.Q(N1902));
  AO22X1 U864(.IN1(N1895),.IN2(n204),.IN3(n1214),.IN4(n925),.Q(N1901));
  AO22X1 U865(.IN1(N1894),.IN2(n204),.IN3(n1214),.IN4(N1884),.Q(N1900));
  AO22X1 U871(.IN1(N1878),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(N1868),.Q(N1884));
  AO22X1 U876(.IN1(N1863),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n954),.Q(N1869));
  AO22X1 U877(.IN1(N1862),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(N1852),.Q(N1868));
  AO22X1 U882(.IN1(N1847),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n157),.Q(N1853));
  AO22X1 U883(.IN1(N1846),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(N1836),.Q(N1852));
  AO22X1 U889(.IN1(N1830),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(N1820),.Q(N1836));
  AO22X1 U894(.IN1(N1815),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n890),.Q(N1821));
  AO22X1 U895(.IN1(N1814),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(N1804),.Q(N1820));
  AO22X1 U897(.IN1(N1802),.IN2(n215),.IN3(n1211),.IN4(n1040),.Q(N1808));
  AO22X1 U901(.IN1(N1798),.IN2(n215),.IN3(n1210),.IN4(N1788),.Q(N1804));
  AO22X1 U905(.IN1(n221),.IN2(N1784),.IN3(s_fract_48_i[11:11]),.IN4(n843),.Q(N1790));
  AO22X1 U907(.IN1(N1782),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(N1772),.Q(N1788));
  AO22X1 U913(.IN1(N1766),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(N1756),.Q(N1772));
  AO22X1 U919(.IN1(N1750),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(N1740),.Q(N1756));
  AO22X1 U922(.IN1(N1737),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n939),.Q(N1743));
  AO22X1 U925(.IN1(N1734),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(N1724),.Q(N1740));
  AO22X1 U931(.IN1(N1718),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(N1708),.Q(N1724));
  AO22X1 U933(.IN1(N1706),.IN2(n226),.IN3(n1226),.IN4(N1696),.Q(N1712));
  AO22X1 U935(.IN1(N1704),.IN2(n226),.IN3(n1227),.IN4(n163),.Q(N1710));
  AO22X1 U936(.IN1(N1703),.IN2(n226),.IN3(n1225),.IN4(n993),.Q(N1709));
  AO22X1 U937(.IN1(N1702),.IN2(n226),.IN3(n1227),.IN4(N1692),.Q(N1708));
  AO22X1 U940(.IN1(N1689),.IN2(n227),.IN3(N1680),.IN4(n1221),.Q(N1695));
  AO22X1 U941(.IN1(n227),.IN2(N1688),.IN3(n1223),.IN4(n1132),.Q(N1694));
  AO22X1 U942(.IN1(N1687),.IN2(n227),.IN3(n1223),.IN4(n1024),.Q(N1693));
  AO22X1 U943(.IN1(N1686),.IN2(n227),.IN3(n1222),.IN4(N1677),.Q(N1692));
  AND2X1 U945(.IN1(N1675),.IN2(n229),.Q(N1680));
  AO22X1 U946(.IN1(N1674),.IN2(n229),.IN3(N1666),.IN4(s_fract_48_i[4:4]),.Q(N1679));
  AO22X1 U947(.IN1(N1673),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1134),.Q(N1678));
  AO22X1 U948(.IN1(N1672),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(N1664),.Q(N1677));
  AND2X1 U950(.IN1(n1208),.IN2(n570),.Q(N1666));
  XOR2X1 U951(.IN1(n570),.IN2(n569),.Q(N1665));
  AO21X1 U952(.IN1(n1137),.IN2(n232),.IN3(n481),.Q(n570));
  XNOR2X1 U955(.IN1(n233),.IN2(s_fract_48_i[1:1]),.Q(n568));
  NAND4X0 U958(.IN1(n580),.IN2(n581),.IN3(n582),.IN4(n583),.QN(n579));
  AOI222X1 U959(.IN1(n861),.IN2(n584),.IN3(n889),.IN4(n585),.IN5(n844),.IN6(n586),.QN(n583));
  AOI22X1 U960(.IN1(n831),.IN2(s_fract_48_i[36:36]),.IN3(n841),.IN4(n587),.QN(n582));
  AO21X1 U961(.IN1(n589),.IN2(n590),.IN3(n1427),.Q(n580));
  AO22X1 U966(.IN1(n603),.IN2(n1057),.IN3(n1290),.IN4(n1036),.Q(n602));
  NAND4X0 U967(.IN1(n604),.IN2(n605),.IN3(n606),.IN4(n607),.QN(n601));
  AOI222X1 U968(.IN1(n1051),.IN2(n608),.IN3(n1005),.IN4(n609),.IN5(n1012),.IN6(n610),.QN(n607));
  AOI22X1 U969(.IN1(n1076),.IN2(n1213),.IN3(n1022),.IN4(n611),.QN(n606));
  AOI22X1 U972(.IN1(n1044),.IN2(n1211),.IN3(n936),.IN4(n619),.QN(n618));
  OA222X1 U976(.IN1(n1317),.IN2(n630),.IN3(n1316),.IN4(n631),.IN5(n1315),.IN6(n632),.Q(n589));
  NAND4X0 U979(.IN1(n637),.IN2(n638),.IN3(n639),.IN4(n640),.QN(n636));
  AOI222X1 U980(.IN1(n944),.IN2(n584),.IN3(n1119),.IN4(n585),.IN5(n1107),.IN6(n586),.QN(n640));
  AOI22X1 U984(.IN1(n572),.IN2(n1216),.IN3(n209),.IN4(n595),.QN(n644));
  NAND4X0 U988(.IN1(n649),.IN2(n650),.IN3(n651),.IN4(n652),.QN(n647));
  AOI222X1 U989(.IN1(n66),.IN2(n608),.IN3(n381),.IN4(n609),.IN5(n478),.IN6(n610),.QN(n652));
  AOI22X1 U990(.IN1(n1063),.IN2(n1214),.IN3(n633),.IN4(n611),.QN(n651));
  AO21X1 U991(.IN1(n653),.IN2(n654),.IN3(n1480),.Q(n649));
  OA221X1 U992(.IN1(n655),.IN2(n616),.IN3(n1099),.IN4(n617),.IN5(n656),.Q(n654));
  AOI22X1 U993(.IN1(n1035),.IN2(n1210),.IN3(n929),.IN4(n619),.QN(n656));
  OA222X1 U996(.IN1(n1318),.IN2(n627),.IN3(n1058),.IN4(n628),.IN5(n1053),.IN6(n629),.Q(n653));
  AO222X1 U998(.IN1(n575),.IN2(n1066),.IN3(n577),.IN4(n904),.IN5(n574),.IN6(n58),.Q(n660));
  AO222X1 U999(.IN1(n578),.IN2(n830),.IN3(n635),.IN4(n876),.IN5(n1387),.IN6(n662),.Q(n659));
  NAND4X0 U1000(.IN1(n663),.IN2(n664),.IN3(n665),.IN4(n666),.QN(n662));
  AOI222X1 U1001(.IN1(n1069),.IN2(n584),.IN3(n597),.IN4(n585),.IN5(n1106),.IN6(n586),.QN(n666));
  AO21X1 U1003(.IN1(n667),.IN2(n668),.IN3(n1427),.Q(n663));
  OA221X1 U1004(.IN1(n592),.IN2(n669),.IN3(n1045),.IN4(n593),.IN5(n670),.Q(n668));
  AOI22X1 U1005(.IN1(n350),.IN2(n1216),.IN3(n806),.IN4(n595),.QN(n670));
  AO22X1 U1008(.IN1(n603),.IN2(n1064),.IN3(n1290),.IN4(n1075),.Q(n674));
  NAND4X0 U1009(.IN1(n675),.IN2(n676),.IN3(n677),.IN4(n678),.QN(n673));
  AOI222X1 U1010(.IN1(n1083),.IN2(n608),.IN3(n432),.IN4(n609),.IN5(n382),.IN6(n610),.QN(n678));
  AOI22X1 U1011(.IN1(n989),.IN2(n1213),.IN3(n634),.IN4(n611),.QN(n677));
  AO21X1 U1012(.IN1(n679),.IN2(n680),.IN3(n1480),.Q(n675));
  OA221X1 U1013(.IN1(n616),.IN2(n681),.IN3(n1358),.IN4(n617),.IN5(n682),.Q(n680));
  AOI22X1 U1014(.IN1(n840),.IN2(n1210),.IN3(n169),.IN4(n619),.QN(n682));
  OA222X1 U1017(.IN1(n1361),.IN2(n627),.IN3(n1360),.IN4(n628),.IN5(n1359),.IN6(n629),.Q(n679));
  OA222X1 U1018(.IN1(n1363),.IN2(n630),.IN3(n871),.IN4(n631),.IN5(n1362),.IN6(n632),.Q(n667));
  AOI222X1 U1023(.IN1(n894),.IN2(n584),.IN3(n202),.IN4(n585),.IN5(n931),.IN6(n586),.QN(n693));
  AOI22X1 U1024(.IN1(n811),.IN2(s_fract_48_i[36:36]),.IN3(n186),.IN4(n587),.QN(n692));
  AO21X1 U1025(.IN1(n694),.IN2(n695),.IN3(n1427),.Q(n690));
  OA221X1 U1026(.IN1(n592),.IN2(n697),.IN3(n1367),.IN4(n593),.IN5(n698),.Q(n695));
  AOI22X1 U1027(.IN1(n908),.IN2(n1217),.IN3(n451),.IN4(n595),.QN(n698));
  AO22X1 U1030(.IN1(n603),.IN2(n976),.IN3(n1289),.IN4(n576),.Q(n702));
  NAND4X0 U1031(.IN1(n703),.IN2(n704),.IN3(n705),.IN4(n706),.QN(n701));
  AOI222X1 U1032(.IN1(n835),.IN2(n608),.IN3(n357),.IN4(n609),.IN5(n900),.IN6(n610),.QN(n706));
  AOI22X1 U1033(.IN1(n657),.IN2(n1214),.IN3(n980),.IN4(n611),.QN(n705));
  AO21X1 U1034(.IN1(n707),.IN2(n708),.IN3(n1480),.Q(n703));
  OA221X1 U1035(.IN1(n616),.IN2(n710),.IN3(n1364),.IN4(n617),.IN5(n711),.Q(n708));
  OA222X1 U1039(.IN1(n1366),.IN2(n627),.IN3(n1365),.IN4(n628),.IN5(n159),.IN6(n629),.Q(n707));
  OA222X1 U1040(.IN1(n1370),.IN2(n630),.IN3(n1369),.IN4(n631),.IN5(n1368),.IN6(n632),.Q(n694));
  AO221X1 U1041(.IN1(n716),.IN2(s_fract_48_i[44:44]),.IN3(n717),.IN4(n661),.IN5(n718),.Q(N1633));
  AOI222X1 U1042(.IN1(n1387),.IN2(n721),.IN3(n1104),.IN4(n635),.IN5(n821),.IN6(n578),.QN(n720));
  AO22X1 U1046(.IN1(n587),.IN2(n713),.IN3(s_fract_48_i[36:36]),.IN4(n863),.Q(n725));
  NAND4X0 U1047(.IN1(n726),.IN2(n727),.IN3(n728),.IN4(n729),.QN(n724));
  OA222X1 U1048(.IN1(n1378),.IN2(n630),.IN3(n1377),.IN4(n631),.IN5(n1376),.IN6(n632),.Q(n729));
  AOI22X1 U1049(.IN1(n921),.IN2(n1217),.IN3(n834),.IN4(n595),.QN(n728));
  AO21X1 U1050(.IN1(n730),.IN2(n731),.IN3(n592),.Q(n726));
  OA221X1 U1051(.IN1(n714),.IN2(n732),.IN3(n1375),.IN4(n715),.IN5(n733),.Q(n731));
  AOI22X1 U1052(.IN1(n1020),.IN2(n1290),.IN3(n507),.IN4(n603),.QN(n733));
  OA222X1 U1057(.IN1(n1374),.IN2(n627),.IN3(n1373),.IN4(n628),.IN5(n1372),.IN6(n629),.Q(n740));
  AOI22X1 U1058(.IN1(n45),.IN2(n1211),.IN3(n854),.IN4(n619),.QN(n739));
  OA22X1 U1059(.IN1(n1371),.IN2(n617),.IN3(n741),.IN4(n616),.Q(n738));
  AOI222X1 U1062(.IN1(n875),.IN2(n600),.IN3(n1003),.IN4(n599),.IN5(n105),.IN6(n598),.QN(n730));
  AO221X1 U1064(.IN1(n744),.IN2(n949),.IN3(n661),.IN4(n746),.IN5(n718),.Q(N1632));
  AOI222X1 U1065(.IN1(n749),.IN2(n1387),.IN3(N362),.IN4(n635),.IN5(N430),.IN6(n578),.QN(n748));
  AND2X1 U1066(.IN1(n750),.IN2(n751),.Q(n578));
  OR2X1 U1067(.IN1(n753),.IN2(n754),.Q(n749));
  AO222X1 U1068(.IN1(n586),.IN2(N515),.IN3(n585),.IN4(N498),.IN5(n584),.IN6(N481),.Q(n754));
  AO221X1 U1069(.IN1(n588),.IN2(N532),.IN3(n696),.IN4(n758),.IN5(n759),.Q(n753));
  AO22X1 U1070(.IN1(n587),.IN2(N464),.IN3(s_fract_48_i[36:36]),.IN4(N447),.Q(n759));
  NAND4X0 U1071(.IN1(n761),.IN2(n762),.IN3(n763),.IN4(n764),.QN(n758));
  OA222X1 U1072(.IN1(N594),.IN2(n630),.IN3(N611),.IN4(n631),.IN5(n1380),.IN6(n632),.Q(n764));
  OR2X1 U1073(.IN1(n765),.IN2(n766),.Q(n632));
  OR2X1 U1074(.IN1(n768),.IN2(n767),.Q(n630));
  AOI22X1 U1075(.IN1(N549),.IN2(n1216),.IN3(N566),.IN4(n595),.QN(n763));
  AND2X1 U1076(.IN1(n768),.IN2(n164),.Q(n595));
  AO21X1 U1077(.IN1(n769),.IN2(n770),.IN3(n592),.Q(n761));
  OA221X1 U1078(.IN1(n771),.IN2(n714),.IN3(N747),.IN4(n715),.IN5(n772),.Q(n770));
  AOI22X1 U1079(.IN1(N651),.IN2(n1290),.IN3(N668),.IN4(n603),.QN(n772));
  AND2X1 U1080(.IN1(n773),.IN2(n177),.Q(n603));
  AO222X1 U1081(.IN1(n610),.IN2(N821),.IN3(n609),.IN4(N804),.IN5(n608),.IN6(N787),.Q(n776));
  AO221X1 U1082(.IN1(n612),.IN2(N838),.IN3(n709),.IN4(n780),.IN5(n781),.Q(n775));
  AO22X1 U1083(.IN1(n611),.IN2(N770),.IN3(n1213),.IN4(N753),.Q(n781));
  NAND3X0 U1084(.IN1(n783),.IN2(n784),.IN3(n785),.QN(n780));
  OA222X1 U1085(.IN1(N900),.IN2(n627),.IN3(n1379),.IN4(n628),.IN5(N934),.IN6(n629),.Q(n785));
  OR2X1 U1086(.IN1(n786),.IN2(n787),.Q(n629));
  OR2X1 U1087(.IN1(n789),.IN2(n788),.Q(n627));
  AOI22X1 U1088(.IN1(N855),.IN2(n1210),.IN3(N872),.IN4(n619),.QN(n784));
  AND2X1 U1089(.IN1(n789),.IN2(n215),.Q(n619));
  OA22X1 U1090(.IN1(N951),.IN2(n617),.IN3(n790),.IN4(n616),.Q(n783));
  AO222X1 U1091(.IN1(n622),.IN2(N974),.IN3(n1226),.IN4(N957),.IN5(n623),.IN6(N991),.Q(n792));
  AND2X1 U1092(.IN1(n793),.IN2(n226),.Q(n622));
  AO222X1 U1093(.IN1(N1036),.IN2(n624),.IN3(n625),.IN4(N1008),.IN5(n626),.IN6(N1025),.Q(n791));
  AND2X1 U1094(.IN1(n794),.IN2(n795),.Q(n625));
  NOR3X0 U1095(.IN1(n1207),.IN2(s_fract_48_i[2:2]),.IN3(n795),.QN(n624));
  AOI222X1 U1096(.IN1(N685),.IN2(n600),.IN3(N702),.IN4(n599),.IN5(N719),.IN6(n598),.QN(n769));
  AND2X1 U1097(.IN1(n797),.IN2(n796),.Q(n599));
  AND2X1 U1099(.IN1(n799),.IN2(n798),.Q(n577));
  AND2X1 U1100(.IN1(n800),.IN2(n68),.Q(n716));
  AO22X1 U1102(.IN1(N1023),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(n1126),.Q(N1029));
  AO22X1 U1103(.IN1(N1022),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(n70),.Q(N1028));
  AO22X1 U1106(.IN1(N1019),.IN2(n232),.IN3(s_fract_48_i[2:2]),.IN4(N1008),.Q(N1025));
  AO22X1 U1109(.IN1(N973),.IN2(n227),.IN3(n1223),.IN4(n974),.Q(N979));
  AO22X1 U1116(.IN1(N854),.IN2(n215),.IN3(n1211),.IN4(n1002),.Q(N860));
  AO22X1 U1127(.IN1(N667),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1036),.Q(N673));
  AO22X1 U1130(.IN1(N616),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1084),.Q(N622));
  AO22X1 U1134(.IN1(N548),.IN2(n164),.IN3(n1217),.IN4(n865),.Q(N554));
  AO22X1 U1142(.IN1(N412),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(N401),.Q(N418));
  AO22X1 U1148(.IN1(N972),.IN2(n227),.IN3(n1220),.IN4(n1115),.Q(N978));
  AO22X1 U1149(.IN1(N955),.IN2(n226),.IN3(n1224),.IN4(n1105),.Q(N961));
  AO22X1 U1154(.IN1(N870),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1035),.Q(N876));
  AO22X1 U1156(.IN1(N836),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n478),.Q(N842));
  AO22X1 U1161(.IN1(N751),.IN2(n204),.IN3(n1213),.IN4(n1121),.Q(N757));
  AO22X1 U1163(.IN1(N717),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n992),.Q(N723));
  AO22X1 U1169(.IN1(N615),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n983),.Q(N621));
  AO22X1 U1173(.IN1(N547),.IN2(n164),.IN3(n1216),.IN4(n922),.Q(N553));
  AO22X1 U1174(.IN1(N530),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1107),.Q(N536));
  AO22X1 U1188(.IN1(N971),.IN2(n227),.IN3(n1220),.IN4(n860),.Q(N977));
  AO22X1 U1190(.IN1(N937),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1103),.Q(N943));
  AO22X1 U1195(.IN1(N852),.IN2(n215),.IN3(n1210),.IN4(n613),.Q(N858));
  AO22X1 U1201(.IN1(N750),.IN2(n204),.IN3(n1214),.IN4(n1070),.Q(N756));
  AO22X1 U1202(.IN1(N733),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1067),.Q(N739));
  AO22X1 U1203(.IN1(N716),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n956),.Q(N722));
  AO22X1 U1206(.IN1(N665),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1075),.Q(N671));
  AO22X1 U1210(.IN1(N597),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n486),.Q(N603));
  AO22X1 U1213(.IN1(N546),.IN2(n164),.IN3(n1216),.IN4(n1087),.Q(N552));
  AO22X1 U1214(.IN1(N529),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1106),.Q(N535));
  AND2X1 U1225(.IN1(N344),.IN2(n123),.Q(N349));
  AO22X1 U1228(.IN1(N970),.IN2(n227),.IN3(n1220),.IN4(n1090),.Q(N976));
  AO22X1 U1229(.IN1(N953),.IN2(n226),.IN3(n1224),.IN4(n1093),.Q(N959));
  AO22X1 U1235(.IN1(N851),.IN2(n215),.IN3(n1210),.IN4(n220),.Q(N857));
  AO22X1 U1236(.IN1(N834),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n900),.Q(N840));
  AO22X1 U1241(.IN1(N749),.IN2(n204),.IN3(n1213),.IN4(n958),.Q(N755));
  AO22X1 U1243(.IN1(N715),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n500),.Q(N721));
  AO22X1 U1246(.IN1(N664),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n576),.Q(N670));
  AO22X1 U1250(.IN1(N596),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1031),.Q(N602));
  AO22X1 U1253(.IN1(N545),.IN2(n164),.IN3(n1216),.IN4(n820),.Q(N551));
  AO22X1 U1265(.IN1(N343),.IN2(n123),.IN3(n1228),.IN4(N334),.Q(N348));
  AND2X1 U1266(.IN1(n1133),.IN2(n802),.Q(N334));
  AO22X1 U1268(.IN1(N986),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n40),.Q(N992));
  AO22X1 U1270(.IN1(N952),.IN2(n226),.IN3(n1225),.IN4(N941),.Q(N958));
  AO22X1 U1271(.IN1(N935),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(N924),.Q(N941));
  AO22X1 U1272(.IN1(N918),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n166),.Q(N924));
  AO22X1 U1274(.IN1(N884),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n854),.Q(N890));
  AO22X1 U1276(.IN1(N850),.IN2(n215),.IN3(n1211),.IN4(n878),.Q(N856));
  AO22X1 U1278(.IN1(N816),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n804),.Q(N822));
  AO22X1 U1283(.IN1(N731),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n105),.Q(N737));
  AO22X1 U1287(.IN1(N663),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1020),.Q(N669));
  AO22X1 U1289(.IN1(N629),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n994),.Q(N635));
  AO22X1 U1292(.IN1(N578),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n834),.Q(N584));
  AO22X1 U1294(.IN1(N544),.IN2(n164),.IN3(n1217),.IN4(n1081),.Q(N550));
  AO22X1 U1295(.IN1(N527),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1074),.Q(N533));
  AO22X1 U1297(.IN1(N493),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n839),.Q(N499));
  AO22X1 U1302(.IN1(N408),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n815),.Q(N414));
  AO22X1 U1306(.IN1(N342),.IN2(n123),.IN3(n1228),.IN4(N333),.Q(N347));
  AO21X1 U1308(.IN1(n949),.IN2(n119),.IN3(n800),.Q(n802));
  AO22X1 U1309(.IN1(N1002),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(N991),.Q(N1008));
  AO22X1 U1310(.IN1(N985),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(N974),.Q(N991));
  AO22X1 U1311(.IN1(N968),.IN2(n227),.IN3(n1221),.IN4(N957),.Q(N974));
  AO22X1 U1312(.IN1(N951),.IN2(n226),.IN3(n1225),.IN4(N940),.Q(N957));
  AO22X1 U1313(.IN1(N934),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(N923),.Q(N940));
  AO22X1 U1314(.IN1(n1379),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(N906),.Q(N923));
  AO22X1 U1315(.IN1(N900),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(N889),.Q(N906));
  AO22X1 U1316(.IN1(N883),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(N872),.Q(N889));
  AO22X1 U1317(.IN1(N866),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(N855),.Q(N872));
  AO22X1 U1318(.IN1(N849),.IN2(n215),.IN3(n1211),.IN4(N838),.Q(N855));
  AO22X1 U1319(.IN1(N832),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(N821),.Q(N838));
  AO22X1 U1320(.IN1(N815),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(N804),.Q(N821));
  AO22X1 U1321(.IN1(N798),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(N787),.Q(N804));
  AO22X1 U1322(.IN1(N781),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(N770),.Q(N787));
  AO22X1 U1323(.IN1(N764),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(N753),.Q(N770));
  AO22X1 U1324(.IN1(N747),.IN2(n204),.IN3(n1213),.IN4(N736),.Q(N753));
  AO22X1 U1325(.IN1(N730),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(N719),.Q(N736));
  AO22X1 U1326(.IN1(N713),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(N702),.Q(N719));
  AO22X1 U1327(.IN1(N696),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(N685),.Q(N702));
  AO22X1 U1328(.IN1(N679),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N668),.Q(N685));
  AO22X1 U1329(.IN1(N662),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(N651),.Q(N668));
  AO22X1 U1330(.IN1(N645),.IN2(n177),.IN3(n1289),.IN4(N634),.Q(N651));
  AO22X1 U1331(.IN1(n1380),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(N617),.Q(N634));
  AO22X1 U1332(.IN1(N611),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(N600),.Q(N617));
  AO22X1 U1333(.IN1(N594),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(N583),.Q(N600));
  AO22X1 U1334(.IN1(N577),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(N566),.Q(N583));
  AO22X1 U1335(.IN1(N560),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N549),.Q(N566));
  AO22X1 U1336(.IN1(N543),.IN2(n164),.IN3(n1217),.IN4(N532),.Q(N549));
  AO22X1 U1337(.IN1(N526),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(N515),.Q(N532));
  AO22X1 U1338(.IN1(N509),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(N498),.Q(N515));
  AO22X1 U1339(.IN1(N492),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N481),.Q(N498));
  AO22X1 U1340(.IN1(N475),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(N464),.Q(N481));
  AO22X1 U1341(.IN1(N458),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(N447),.Q(N464));
  AO22X1 U1342(.IN1(N441),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(N430),.Q(N447));
  AO22X1 U1343(.IN1(N424),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N413),.Q(N430));
  AO22X1 U1344(.IN1(N407),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(N396),.Q(N413));
  AO22X1 U1345(.IN1(N390),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(N379),.Q(N396));
  AO22X1 U1346(.IN1(N373),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N362),.Q(N379));
  AO22X1 U1347(.IN1(N356),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(N346),.Q(N362));
  AO22X1 U1348(.IN1(N341),.IN2(n123),.IN3(n1230),.IN4(N332),.Q(N346));
  XNOR2X1 U1349(.IN1(n122),.IN2(n988),.Q(N332));
  XNOR2X1 U1351(.IN1(n118),.IN2(s_fract_48_i[46:46]),.Q(n745));
  post_norm_mul_DW01_inc_0_inj add_233(.A({n1197,s_expo2b[7:0]}),.SUM({N3354,N3353,N3352,N3351,N3350,N3349,N3348,N3347,N3346}));
  post_norm_mul_DW01_inc_1_inj add_222(.A(s_frac2a[47:23]),.SUM({N3302,N3301,N3300,N3299,N3298,N3297,N3296,N3295,N3294,N3293,N3292,N3291,N3290,N3289,N3288,N3287,N3286,N3285,N3284,N3283,N3282,N3281,N3280,N3279,N3278}));
  post_norm_mul_DW01_sub_1_inj sub_154(.A(s_zeros),.B(s_exp_10a[5:0]),.CI(1'b0),.DIFF({N3024,N3023,N3022,N3021,N3020,N3019}));
  post_norm_mul_DW01_sub_2_inj sub_141(.A(s_exp_10a),.B({1'b0,1'b0,1'b0,1'b0,s_zeros}),.CI(1'b0),.DIFF(s_exp_10b));
  HADDX1 desc1139(.A0(\add_105_I47_L14036_C136/carry[2] ),.B0(N2334),.C1(\add_105_I47_L14036_C136/carry[3] ),.SO(N2344));
  HADDX1 desc1140(.A0(\add_105_I14_L14036_C136/carry[4] ),.B0(N1808),.C1(\add_105_I14_L14036_C136/carry[5] ),.SO(N1818));
  HADDX1 desc1141(.A0(\add_105_I9_L14036_C136/carry[4] ),.B0(N1728),.C1(\add_105_I9_L14036_C136/carry[5] ),.SO(N1738));
  HADDX1 desc1142(.A0(\add_105_I8_L14036_C136/carry[3] ),.B0(N1711),.C1(\add_105_I8_L14036_C136/carry[4] ),.SO(N1721));
  HADDX1 desc1143(.A0(N1695),.B0(\add_105_I7_L14036_C136/carry[3] ),.C1(\add_105_I7_L14036_C136/carry[4] ),.SO(N1705));
  HADDX1 desc1144(.A0(N1679),.B0(\add_105_I6_L14036_C136/carry[2] ),.C1(\add_105_I6_L14036_C136/carry[3] ),.SO(N1688));
  HADDX1 desc1145(.A0(N1026),.B0(N1025),.C1(\add_90_I46_L14036_C132/carry[2] ),.SO(N1037));
  HADDX1 desc1146(.A0(\add_90_I46_L14036_C132/carry[3] ),.B0(N1028),.C1(\add_90_I46_L14036_C132/carry[4] ),.SO(N1039));
  HADDX1 desc1147(.A0(\add_90_I44_L14036_C132/carry[2] ),.B0(N993),.C1(\add_90_I44_L14036_C132/carry[3] ),.SO(N1004));
  HADDX1 desc1148(.A0(N976),.B0(\add_90_I43_L14036_C132/carry[2] ),.C1(\add_90_I43_L14036_C132/carry[3] ),.SO(N987));
  HADDX1 desc1149(.A0(N978),.B0(\add_90_I43_L14036_C132/carry[4] ),.C1(\add_90_I43_L14036_C132/carry[5] ),.SO(N989));
  HADDX1 desc1150(.A0(\add_90_I41_L14036_C132/carry[3] ),.B0(N943),.C1(\add_90_I41_L14036_C132/carry[4] ),.SO(N954));
  HADDX1 desc1151(.A0(\add_90_I40_L14036_C132/carry[2] ),.B0(N925),.C1(\add_90_I40_L14036_C132/carry[3] ),.SO(N936));
  HADDX1 desc1152(.A0(\add_90_I36_L14036_C132/carry[4] ),.B0(N859),.C1(\add_90_I36_L14036_C132/carry[5] ),.SO(N870));
  HADDX1 desc1153(.A0(\add_90_I33_L14036_C132/carry[3] ),.B0(N807),.C1(\add_90_I33_L14036_C132/carry[4] ),.SO(N818));
  HADDX1 desc1154(.A0(\add_90_I32_L14036_C132/carry[4] ),.B0(N791),.C1(\add_90_I32_L14036_C132/carry[5] ),.SO(N802));
  HADDX1 desc1155(.A0(\add_90_I29_L14036_C132/carry[2] ),.B0(N738),.C1(\add_90_I29_L14036_C132/carry[3] ),.SO(N749));
  HADDX1 desc1156(.A0(\add_90_I27_L14036_C132/carry[2] ),.B0(N704),.C1(\add_90_I27_L14036_C132/carry[3] ),.SO(N715));
  HADDX1 desc1157(.A0(\add_90_I19_L14036_C132/carry[3] ),.B0(N569),.C1(\add_90_I19_L14036_C132/carry[4] ),.SO(N580));
  HADDX1 desc1158(.A0(\add_90_I17_L14036_C132/carry[2] ),.B0(N534),.C1(\add_90_I17_L14036_C132/carry[3] ),.SO(N545));
  HADDX1 desc1159(.A0(N535),.B0(\add_90_I17_L14036_C132/carry[3] ),.C1(\add_90_I17_L14036_C132/carry[4] ),.SO(N546));
  HADDX1 desc1160(.A0(\add_90_I10_L14036_C132/carry[4] ),.B0(N417),.C1(\add_90_I10_L14036_C132/carry[5] ),.SO(N428));
  HADDX1 desc1161(.A0(\add_90_I8_L14036_C132/carry[2] ),.B0(N381),.C1(\add_90_I8_L14036_C132/carry[3] ),.SO(N392));
  HADDX1 desc1162(.A0(N333),.B0(N332),.C1(\add_90_I5_L14036_C132/carry[2] ),.SO(N342));
  FADDX1 desc1163(.A(N2993),.B(n1294),.CI(\sub_0_root_add_0_root_add_148/carry[1] ),.CO(\sub_0_root_add_0_root_add_148/carry[2] ),.S(N3000));
  DFFX2 desc1164(.D(fract_48_i[42:42]),.CLK(clk_i),.Q(s_fract_48_i[42:42]),.QN(n123));
  DFFX2 desc1165(.D(fract_48_i[36:36]),.CLK(clk_i),.Q(s_fract_48_i[36:36]),.QN(n152));
  DFFX2 desc1166(.D(fract_48_i[30:30]),.CLK(clk_i),.Q(s_fract_48_i[30:30]),.QN(n164));
  DFFX2 desc1167(.D(fract_48_i[24:24]),.CLK(clk_i),.Q(s_fract_48_i[24:24]),.QN(n177));
  DFFX2 desc1168(.D(fract_48_i[18:18]),.CLK(clk_i),.Q(s_fract_48_i[18:18]),.QN(n204));
  DFFX2 desc1169(.D(fract_48_i[6:6]),.CLK(clk_i),.Q(s_fract_48_i[6:6]),.QN(n226));
  DFFX2 desc1170(.D(fract_48_i[5:5]),.CLK(clk_i),.Q(s_fract_48_i[5:5]),.QN(n227));
  DFFX1 desc1171(.D(fract_48_i[1:1]),.CLK(clk_i),.Q(s_fract_48_i[1:1]),.QN(n1206));
  DFFX1 desc1172(.D(N3083),.CLK(clk_i),.Q(s_shr2[2:2]),.QN(n71));
  DFFX2 desc1173(.D(fract_48_i[2:2]),.CLK(clk_i),.Q(s_fract_48_i[2:2]),.QN(n232));
  DFFX1 desc1174(.D(fract_48_i[12:12]),.CLK(clk_i),.Q(s_fract_48_i[12:12]),.QN(n215));
  DFFX2 desc1175(.D(fract_48_i[44:44]),.CLK(clk_i),.Q(s_fract_48_i[44:44]),.QN(n119));
  DELLN1X2 U4(.INP(N2297),.Z(n1));
  XNOR2X1 U5(.IN1(n962),.IN2(\add_105_I45_L14036_C136/carry[5] ),.Q(N2315));
  AOI222X1 U6(.IN1(n383),.IN2(n314),.IN3(n1231),.IN4(n178),.IN5(n384),.IN6(n2),.QN(n115));
  HADDX2 U7(.A0(\add_105_I29_L14036_C136/carry[4] ),.B0(N2048),.C1(\add_105_I29_L14036_C136/carry[5] ),.SO(N2058));
  AO22X1 U8(.IN1(N2313),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n314),.Q(n2));
  HADDX1 U9(.A0(\add_105_I45_L14036_C136/carry[3] ),.B0(N2303),.C1(\add_105_I45_L14036_C136/carry[4] ),.SO(N2313));
  AO22X1 U10(.IN1(n1),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n178),.Q(n314));
  DELLN1X2 U11(.INP(N2281),.Z(n3));
  HADDX2 U12(.A0(\add_105_I40_L14036_C136/carry[3] ),.B0(N2223),.C1(\add_105_I40_L14036_C136/carry[4] ),.SO(N2233));
  DELLN1X2 U13(.INP(N2298),.Z(n4));
  XNOR2X1 U14(.IN1(n880),.IN2(\add_105_I31_L14036_C136/carry[5] ),.Q(N2091));
  AOI222X1 U15(.IN1(n853),.IN2(n368),.IN3(n872),.IN4(n1216),.IN5(n816),.IN6(n369),.QN(n411));
  DELLN1X2 U16(.INP(N1688),.Z(n5));
  AO22X1 U17(.IN1(N2311),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n896),.Q(n8));
  HADDX2 U18(.A0(\add_105_I19_L14036_C136/carry[4] ),.B0(N1888),.C1(\add_105_I19_L14036_C136/carry[5] ),.SO(N1898));
  HADDX2 U19(.A0(\add_105_I32_L14036_C136/carry[3] ),.B0(N2095),.C1(\add_105_I32_L14036_C136/carry[4] ),.SO(N2105));
  HADDX2 U20(.A0(\add_105_I27_L14036_C136/carry[4] ),.B0(N2016),.C1(\add_105_I27_L14036_C136/carry[5] ),.SO(N2026));
  HADDX2 U21(.A0(\add_105_I16_L14036_C136/carry[3] ),.B0(N1839),.C1(\add_105_I16_L14036_C136/carry[4] ),.SO(N1849));
  DELLN2X2 U22(.INP(N1689),.Z(n9));
  DELLN2X2 U23(.INP(N2331),.Z(n10));
  AO22X2 U24(.IN1(N2329),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n2),.Q(n11));
  AO22X1 U25(.IN1(N2331),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n29),.Q(N2337));
  AO22X1 U26(.IN1(n10),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n29),.Q(n31));
  XNOR2X1 U27(.IN1(n12),.IN2(\add_105_I46_L14036_C136/carry[5] ),.Q(N2331));
  AOI22X1 U28(.IN1(N2315),.IN2(n47),.IN3(s_fract_48_i[44:44]),.IN4(n48),.QN(n12));
  DELLN1X2 U29(.INP(N1899),.Z(n13));
  DELLN1X2 U30(.INP(N2155),.Z(n14));
  DELLN1X2 U31(.INP(N2011),.Z(n15));
  AO22X2 U32(.IN1(N1850),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n207),.Q(n16));
  HADDX1 U33(.A0(\add_105_I16_L14036_C136/carry[4] ),.B0(N1840),.C1(\add_105_I16_L14036_C136/carry[5] ),.SO(N1850));
  AO22X1 U34(.IN1(N2121),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n817),.Q(n17));
  HADDX2 U35(.A0(\add_105_I9_L14036_C136/carry[2] ),.B0(N1726),.C1(\add_105_I9_L14036_C136/carry[3] ),.SO(N1736));
  XNOR2X1 U36(.IN1(\add_105_I26_L14036_C136/carry[5] ),.IN2(n18),.Q(N2011));
  AOI22X1 U37(.IN1(N1995),.IN2(n177),.IN3(n1289),.IN4(N1985),.QN(n18));
  DELLN1X2 U38(.INP(N2123),.Z(n19));
  DELLN1X2 U39(.INP(N2107),.Z(n20));
  DELLN1X2 U40(.INP(N2267),.Z(n21));
  XNOR2X2 U41(.IN1(n508),.IN2(\add_105_I42_L14036_C136/carry[5] ),.Q(N2267));
  DELLN2X2 U42(.INP(N1739),.Z(n22));
  DELLN2X2 U43(.INP(N1851),.Z(n23));
  DELLN2X2 U44(.INP(N1931),.Z(n24));
  AO22X1 U45(.IN1(N2187),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n1073),.Q(N2193));
  DELLN2X2 U46(.INP(N2139),.Z(n25));
  XNOR2X2 U47(.IN1(n866),.IN2(\add_105_I37_L14036_C136/carry[5] ),.Q(N2187));
  AO22X2 U48(.IN1(N1914),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n996),.Q(n26));
  AO22X2 U49(.IN1(N1912),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1050),.Q(n27));
  AO22X2 U50(.IN1(n210),.IN2(N1849),.IN3(s_fract_48_i[15:15]),.IN4(n924),.Q(n28));
  AO22X1 U51(.IN1(N2315),.IN2(n47),.IN3(s_fract_48_i[44:44]),.IN4(n48),.Q(n29));
  HADDX2 U52(.A0(\add_105_I13_L14036_C136/carry[4] ),.B0(N1792),.C1(\add_105_I13_L14036_C136/carry[5] ),.SO(N1802));
  HADDX2 U53(.A0(\add_105_I29_L14036_C136/carry[2] ),.B0(N2046),.C1(\add_105_I29_L14036_C136/carry[3] ),.SO(N2056));
  HADDX2 U54(.A0(\add_105_I26_L14036_C136/carry[3] ),.B0(N1999),.C1(\add_105_I26_L14036_C136/carry[4] ),.SO(N2009));
  HADDX2 U55(.A0(\add_105_I11_L14036_C136/carry[4] ),.B0(N1760),.C1(\add_105_I11_L14036_C136/carry[5] ),.SO(N1770));
  AO22X2 U56(.IN1(N2009),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1071),.Q(n30));
  AO22X2 U57(.IN1(n152),.IN2(N2186),.IN3(s_fract_48_i[36:36]),.IN4(n1131),.Q(n32));
  HADDX1 U58(.A0(\add_105_I37_L14036_C136/carry[4] ),.B0(N2176),.C1(\add_105_I37_L14036_C136/carry[5] ),.SO(N2186));
  AO22X2 U59(.IN1(N2074),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n807),.Q(n33));
  HADDX1 U60(.A0(\add_105_I30_L14036_C136/carry[4] ),.B0(N2064),.C1(\add_105_I30_L14036_C136/carry[5] ),.SO(N2074));
  AO22X1 U61(.IN1(N2058),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n645),.Q(n807));
  HADDX2 U62(.A0(\add_105_I11_L14036_C136/carry[3] ),.B0(N1759),.C1(\add_105_I11_L14036_C136/carry[4] ),.SO(N1769));
  AO22X1 U63(.IN1(N1752),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n230),.Q(n34));
  HADDX2 U64(.A0(\add_105_I14_L14036_C136/carry[3] ),.B0(N1807),.C1(\add_105_I14_L14036_C136/carry[4] ),.SO(N1817));
  AOI22X2 U65(.IN1(N2326),.IN2(n118),.IN3(s_fract_48_i[45:45]),.IN4(N2316),.QN(n35));
  AO22X2 U66(.IN1(N2310),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(N2300),.Q(N2316));
  AOI221X1 U67(.IN1(n347),.IN2(N1884),.IN3(n520),.IN4(n429),.IN5(n521),.QN(n80));
  HADDX1 U68(.A0(\add_90_I46_L14036_C132/carry[2] ),.B0(N1027),.C1(\add_90_I46_L14036_C132/carry[3] ),.SO(N1038));
  AOI222X2 U69(.IN1(n624),.IN2(N1038),.IN3(n625),.IN4(N1010),.IN5(n626),.IN6(N1027),.QN(n86));
  AOI221X1 U70(.IN1(n588),.IN2(n1081),.IN3(n724),.IN4(n696),.IN5(n725),.QN(n82));
  OAI221X1 U71(.IN1(n751),.IN2(n38),.IN3(n36),.IN4(n37),.IN5(n39),.QN(n685));
  INVX32 U72(.INP(n577),.ZN(n36));
  INVX32 U73(.INP(n1120),.ZN(n37));
  AND4X1 U74(.IN1(n691),.IN2(n690),.IN3(n692),.IN4(n693),.Q(n38));
  AOI22X1 U75(.IN1(n578),.IN2(n850),.IN3(n635),.IN4(n911),.QN(n39));
  AO22X1 U76(.IN1(N612),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1068),.Q(N618));
  DELLN1X2 U77(.INP(N975),.Z(n40));
  HADDX2 U78(.A0(N2284),.B0(N2285),.C1(\add_105_I44_L14036_C136/carry[2] ),.SO(N2295));
  AO22X1 U79(.IN1(N2295),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n895),.Q(N2301));
  HADDX2 U80(.A0(N1772),.B0(N1773),.C1(\add_105_I12_L14036_C136/carry[2] ),.SO(N1783));
  AO22X1 U81(.IN1(N2343),.IN2(n69),.IN3(n1205),.IN4(n42),.Q(n41));
  HADDX2 U82(.A0(\add_105_I30_L14036_C136/carry[2] ),.B0(n191),.C1(\add_105_I30_L14036_C136/carry[3] ),.SO(N2072));
  AO22X1 U83(.IN1(N1751),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n852),.Q(N1757));
  AO22X1 U84(.IN1(N1751),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n852),.Q(n153));
  AO22X1 U85(.IN1(N1783),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1091),.Q(N1789));
  AO22X1 U86(.IN1(N1783),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1091),.Q(n155));
  HADDX2 U87(.A0(\add_105_I46_L14036_C136/carry[2] ),.B0(N2318),.C1(\add_105_I46_L14036_C136/carry[3] ),.SO(N2328));
  AO22X1 U88(.IN1(N1831),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n620),.Q(N1837));
  AO22X1 U89(.IN1(N1943),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n243),.Q(N1949));
  AO22X1 U90(.IN1(N1943),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n243),.Q(n168));
  HADDX2 U91(.A0(N2268),.B0(N2269),.C1(\add_105_I43_L14036_C136/carry[2] ),.SO(N2279));
  HADDX2 U92(.A0(N1820),.B0(N1821),.C1(\add_105_I15_L14036_C136/carry[2] ),.SO(N1831));
  HADDX2 U93(.A0(N2348),.B0(N2349),.C1(\add_105_I48_L14036_C136/carry[2] ),.SO(N2359));
  HADDX1 U94(.A0(\add_105_I48_L14036_C136/carry[2] ),.B0(N2350),.C1(\add_105_I48_L14036_C136/carry[3] ),.SO(N2360));
  AO22X1 U95(.IN1(N2327),.IN2(n118),.IN3(s_fract_48_i[45:45]),.IN4(n8),.Q(N2333));
  HADDX2 U96(.A0(N2316),.B0(N2317),.C1(\add_105_I46_L14036_C136/carry[2] ),.SO(N2327));
  HADDX2 U97(.A0(\add_105_I45_L14036_C136/carry[2] ),.B0(N2302),.C1(\add_105_I45_L14036_C136/carry[3] ),.SO(N2312));
  HADDX2 U98(.A0(\add_105_I43_L14036_C136/carry[3] ),.B0(N2271),.C1(\add_105_I43_L14036_C136/carry[4] ),.SO(N2281));
  HADDX2 U99(.A0(\add_105_I46_L14036_C136/carry[3] ),.B0(N2319),.C1(\add_105_I46_L14036_C136/carry[4] ),.SO(N2329));
  HADDX2 U100(.A0(\add_105_I47_L14036_C136/carry[3] ),.B0(N2335),.C1(\add_105_I47_L14036_C136/carry[4] ),.SO(N2345));
  AO22X1 U101(.IN1(N2329),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n2),.Q(N2335));
  HADDX2 U102(.A0(\add_105_I28_L14036_C136/carry[2] ),.B0(N2030),.C1(\add_105_I28_L14036_C136/carry[3] ),.SO(N2040));
  DELLN1X2 U103(.INP(N2333),.Z(n42));
  AO22X1 U104(.IN1(N2312),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n148),.Q(n43));
  AOI221X1 U105(.IN1(n1454),.IN2(n62),.IN3(n434),.IN4(n1453),.IN5(n435),.QN(n116));
  HADDX2 U106(.A0(N994),.B0(\add_90_I44_L14036_C132/carry[3] ),.C1(\add_90_I44_L14036_C132/carry[4] ),.SO(N1005));
  HADDX2 U109(.A0(\add_90_I37_L14036_C132/carry[4] ),.B0(N876),.C1(\add_90_I37_L14036_C132/carry[5] ),.SO(N887));
  AO22X1 U110(.IN1(N562),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n908),.Q(n451));
  AO22X1 U111(.IN1(N988),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1008),.Q(n193));
  AO22X1 U112(.IN1(N988),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1008),.Q(N994));
  HADDX2 U113(.A0(\add_90_I13_L14036_C132/carry[3] ),.B0(N467),.C1(\add_90_I13_L14036_C132/carry[4] ),.SO(N478));
  HADDX2 U114(.A0(N430),.B0(N431),.C1(\add_90_I11_L14036_C132/carry[2] ),.SO(N442));
  HADDX2 U115(.A0(N498),.B0(N499),.C1(\add_90_I15_L14036_C132/carry[2] ),.SO(N510));
  HADDX2 U116(.A0(\add_90_I19_L14036_C132/carry[4] ),.B0(N570),.C1(\add_90_I19_L14036_C132/carry[5] ),.SO(N581));
  HADDX2 U117(.A0(\add_90_I20_L14036_C132/carry[4] ),.B0(N587),.C1(\add_90_I20_L14036_C132/carry[5] ),.SO(N598));
  HADDX1 U118(.A0(\add_90_I42_L14036_C132/carry[2] ),.B0(N959),.C1(\add_90_I42_L14036_C132/carry[3] ),.SO(N970));
  NAND3X1 U119(.IN1(n69),.IN2(n68),.IN3(n557),.QN(n558));
  HADDX2 U120(.A0(\add_90_I34_L14036_C132/carry[4] ),.B0(N825),.C1(\add_90_I34_L14036_C132/carry[5] ),.SO(N836));
  HADDX2 U121(.A0(\add_90_I38_L14036_C132/carry[4] ),.B0(n886),.C1(\add_90_I38_L14036_C132/carry[5] ),.SO(N904));
  HADDX2 U122(.A0(\add_90_I27_L14036_C132/carry[4] ),.B0(N706),.C1(\add_90_I27_L14036_C132/carry[5] ),.SO(N717));
  HADDX2 U123(.A0(\add_90_I17_L14036_C132/carry[4] ),.B0(N536),.C1(\add_90_I17_L14036_C132/carry[5] ),.SO(N547));
  HADDX2 U124(.A0(\add_90_I42_L14036_C132/carry[3] ),.B0(N960),.C1(\add_90_I42_L14036_C132/carry[4] ),.SO(N971));
  HADDX2 U125(.A0(N977),.B0(\add_90_I43_L14036_C132/carry[3] ),.C1(\add_90_I43_L14036_C132/carry[4] ),.SO(N988));
  HADDX2 U126(.A0(\add_90_I29_L14036_C132/carry[3] ),.B0(N739),.C1(\add_90_I29_L14036_C132/carry[4] ),.SO(N750));
  HADDX1 U127(.A0(N1011),.B0(\add_90_I45_L14036_C132/carry[3] ),.C1(\add_90_I45_L14036_C132/carry[4] ),.SO(N1022));
  HADDX2 U128(.A0(\add_90_I32_L14036_C132/carry[3] ),.B0(N790),.C1(\add_90_I32_L14036_C132/carry[4] ),.SO(N801));
  HADDX2 U129(.A0(\add_90_I35_L14036_C132/carry[3] ),.B0(N841),.C1(\add_90_I35_L14036_C132/carry[4] ),.SO(N852));
  HADDX2 U130(.A0(\add_90_I39_L14036_C132/carry[3] ),.B0(N909),.C1(\add_90_I39_L14036_C132/carry[4] ),.SO(N920));
  DELLN1X2 U131(.INP(N822),.Z(n44));
  DELLN1X2 U132(.INP(N856),.Z(n45));
  AOI222X2 U133(.IN1(n610),.IN2(n44),.IN3(n609),.IN4(n804),.IN5(n608),.IN6(n902),.QN(n85));
  HADDX2 U134(.A0(N855),.B0(N856),.C1(\add_90_I36_L14036_C132/carry[2] ),.SO(N867));
  HADDX2 U135(.A0(\add_90_I45_L14036_C132/carry[2] ),.B0(N1010),.C1(\add_90_I45_L14036_C132/carry[3] ),.SO(N1021));
  AO22X1 U136(.IN1(N1021),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(N1010),.Q(N1027));
  XNOR2X2 U137(.IN1(n684),.IN2(\add_90_I35_L14036_C132/carry[5] ),.Q(N854));
  HADDX2 U138(.A0(\add_90_I22_L14036_C132/carry[4] ),.B0(N621),.C1(\add_90_I22_L14036_C132/carry[5] ),.SO(N632));
  HADDX2 U139(.A0(\add_90_I18_L14036_C132/carry[4] ),.B0(N553),.C1(\add_90_I18_L14036_C132/carry[5] ),.SO(N564));
  HADDX2 U140(.A0(\add_90_I15_L14036_C132/carry[3] ),.B0(N501),.C1(\add_90_I15_L14036_C132/carry[4] ),.SO(N512));
  HADDX2 U141(.A0(\add_90_I25_L14036_C132/carry[4] ),.B0(N672),.C1(\add_90_I25_L14036_C132/carry[5] ),.SO(N683));
  HADDX2 U142(.A0(\add_90_I40_L14036_C132/carry[4] ),.B0(N927),.C1(\add_90_I40_L14036_C132/carry[5] ),.SO(N938));
  HADDX2 U143(.A0(\add_90_I42_L14036_C132/carry[4] ),.B0(N961),.C1(\add_90_I42_L14036_C132/carry[5] ),.SO(N972));
  HADDX2 U144(.A0(\add_90_I16_L14036_C132/carry[4] ),.B0(N519),.C1(\add_90_I16_L14036_C132/carry[5] ),.SO(N530));
  HADDX2 U145(.A0(\add_90_I44_L14036_C132/carry[4] ),.B0(N995),.C1(\add_90_I44_L14036_C132/carry[5] ),.SO(N1006));
  HADDX2 U146(.A0(\add_90_I12_L14036_C132/carry[3] ),.B0(N450),.C1(\add_90_I12_L14036_C132/carry[4] ),.SO(N461));
  HADDX2 U147(.A0(\add_90_I12_L14036_C132/carry[2] ),.B0(N449),.C1(\add_90_I12_L14036_C132/carry[3] ),.SO(N460));
  HADDX2 U148(.A0(\add_90_I13_L14036_C132/carry[4] ),.B0(N468),.C1(\add_90_I13_L14036_C132/carry[5] ),.SO(N479));
  HADDX2 U149(.A0(\add_90_I12_L14036_C132/carry[4] ),.B0(N451),.C1(\add_90_I12_L14036_C132/carry[5] ),.SO(N462));
  HADDX2 U150(.A0(\add_90_I15_L14036_C132/carry[4] ),.B0(N502),.C1(\add_90_I15_L14036_C132/carry[5] ),.SO(N513));
  HADDX2 U151(.A0(\add_90_I29_L14036_C132/carry[4] ),.B0(N740),.C1(\add_90_I29_L14036_C132/carry[5] ),.SO(N751));
  AOI222X2 U152(.IN1(N417),.IN2(n575),.IN3(n577),.IN4(n64),.IN5(n574),.IN6(n914),.QN(n1190));
  XOR2X2 U153(.IN1(\add_90_I45_L14036_C132/carry[5] ),.IN2(N1013),.Q(N1024));
  XOR2X2 U154(.IN1(\add_90_I44_L14036_C132/carry[5] ),.IN2(N996),.Q(N1007));
  AOI22X1 U155(.IN1(n171),.IN2(N582),.IN3(s_fract_48_i[28:28]),.IN4(n884),.QN(n46));
  XNOR2X1 U156(.IN1(\add_90_I20_L14036_C132/carry[5] ),.IN2(n46),.Q(N599));
  HADDX2 U157(.A0(N365),.B0(\add_90_I7_L14036_C132/carry[3] ),.C1(\add_90_I7_L14036_C132/carry[4] ),.SO(N376));
  XNOR2X2 U158(.IN1(n745),.IN2(n119),.Q(n803));
  HADDX2 U159(.A0(\add_105_I39_L14036_C136/carry[3] ),.B0(N2207),.C1(\add_105_I39_L14036_C136/carry[4] ),.SO(N2217));
  HADDX2 U160(.A0(\add_105_I41_L14036_C136/carry[3] ),.B0(N2239),.C1(\add_105_I41_L14036_C136/carry[4] ),.SO(N2249));
  AO22X2 U161(.IN1(N1817),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1142),.Q(n810));
  INVX0 U162(.INP(s_fract_48_i[44:44]),.ZN(n47));
  XOR2X2 U163(.IN1(n802),.IN2(n801),.Q(N333));
  HADDX2 U164(.A0(\add_105_I22_L14036_C136/carry[2] ),.B0(N1934),.C1(\add_105_I22_L14036_C136/carry[3] ),.SO(N1944));
  HADDX2 U165(.A0(\add_105_I22_L14036_C136/carry[4] ),.B0(N1936),.C1(\add_105_I22_L14036_C136/carry[5] ),.SO(N1946));
  AO22X2 U166(.IN1(N1867),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n919),.Q(N1873));
  AO22X2 U167(.IN1(n24),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1029),.Q(N1937));
  AO22X2 U168(.IN1(N1947),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(N1937),.Q(N1953));
  XNOR2X2 U169(.IN1(n873),.IN2(\add_105_I23_L14036_C136/carry[5] ),.Q(N1963));
  AO22X2 U170(.IN1(N1979),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n943),.Q(N1985));
  AO22X2 U171(.IN1(N2027),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1089),.Q(N2033));
  AO22X2 U172(.IN1(N2056),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n205),.Q(N2062));
  AO22X2 U173(.IN1(N2075),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n1052),.Q(N2081));
  AO22X2 U174(.IN1(n19),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n1065),.Q(N2129));
  AO22X2 U175(.IN1(N2120),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n819),.Q(N2126));
  AO22X2 U176(.IN1(N2153),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n909),.Q(N2159));
  AO22X2 U177(.IN1(N2185),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n742),.Q(N2191));
  AO22X2 U178(.IN1(N2184),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n723),.Q(N2190));
  AO22X2 U179(.IN1(N2216),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n823),.Q(N2222));
  AO22X2 U180(.IN1(N2264),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n917),.Q(N2270));
  AO22X2 U181(.IN1(N2299),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n52),.Q(n48));
  AO22X2 U182(.IN1(N1913),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1060),.Q(n49));
  DELLN1X2 U183(.INP(N1833),.Z(n50));
  HADDX2 U184(.A0(N1724),.B0(N1725),.C1(\add_105_I9_L14036_C136/carry[2] ),.SO(N1735));
  HADDX2 U185(.A0(\add_105_I15_L14036_C136/carry[2] ),.B0(N1822),.C1(\add_105_I15_L14036_C136/carry[3] ),.SO(N1832));
  HADDX2 U186(.A0(\add_105_I16_L14036_C136/carry[2] ),.B0(N1838),.C1(\add_105_I16_L14036_C136/carry[3] ),.SO(N1848));
  HADDX2 U187(.A0(\add_105_I10_L14036_C136/carry[2] ),.B0(N1742),.C1(\add_105_I10_L14036_C136/carry[3] ),.SO(N1752));
  AO22X1 U188(.IN1(N2058),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n645),.Q(N2064));
  HADDX1 U189(.A0(\add_105_I10_L14036_C136/carry[4] ),.B0(N1744),.C1(\add_105_I10_L14036_C136/carry[5] ),.SO(N1754));
  AO22X1 U190(.IN1(N1738),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n945),.Q(N1744));
  AO22X1 U191(.IN1(N2025),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n30),.Q(N2031));
  AO22X1 U192(.IN1(N1770),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n912),.Q(N1776));
  AO22X1 U193(.IN1(N427),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1066),.Q(N433));
  AO22X1 U194(.IN1(N2263),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n107),.Q(N2269));
  AO22X1 U195(.IN1(N2232),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(N2222),.Q(n106));
  AO22X1 U196(.IN1(n152),.IN2(N2186),.IN3(s_fract_48_i[36:36]),.IN4(n1131),.Q(N2192));
  AO22X1 U197(.IN1(N2072),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N2062),.Q(n132));
  AO22X1 U198(.IN1(N2026),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n183),.Q(N2032));
  AO22X1 U199(.IN1(N2026),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n183),.Q(n217));
  AO22X1 U200(.IN1(N1769),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n1102),.Q(N1775));
  AO22X1 U201(.IN1(N444),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n830),.Q(N450));
  AO22X1 U202(.IN1(N1769),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n1102),.Q(n203));
  AO22X1 U203(.IN1(N1722),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n898),.Q(N1728));
  AO22X1 U204(.IN1(N480),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n841),.Q(n861));
  AO22X1 U205(.IN1(N2216),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n823),.Q(n192));
  AO22X1 U206(.IN1(N886),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n169),.Q(N892));
  AO22X1 U207(.IN1(N922),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n818),.Q(n1009));
  AOI222X1 U208(.IN1(n383),.IN2(n148),.IN3(n1229),.IN4(n103),.IN5(n384),.IN6(n43),.QN(n109));
  AO22X1 U209(.IN1(n134),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n32),.Q(n700));
  AO22X1 U210(.IN1(N1978),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n836),.Q(N1984));
  AO22X1 U211(.IN1(N783),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n980),.Q(N789));
  AO22X1 U212(.IN1(N1962),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n195),.Q(N1968));
  AO22X1 U213(.IN1(n131),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n816),.Q(n853));
  AO22X1 U214(.IN1(n14),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n1016),.Q(n1061));
  AO22X1 U215(.IN1(n135),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n217),.Q(n645));
  AO22X1 U216(.IN1(N1834),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n891),.Q(N1840));
  AO22X1 U217(.IN1(N1883),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(N1873),.Q(N1889));
  AO22X1 U218(.IN1(N613),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1028),.Q(n404));
  AO22X1 U219(.IN1(N682),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n1064),.Q(N688));
  AO22X1 U220(.IN1(N701),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n1000),.Q(n1018));
  AO22X1 U221(.IN1(N477),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n186),.Q(N483));
  AO22X1 U222(.IN1(N443),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n850),.Q(N449));
  AO22X1 U223(.IN1(N463),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n831),.Q(N469));
  AO22X1 U224(.IN1(N1831),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n620),.Q(n157));
  AO22X1 U225(.IN1(N1815),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n890),.Q(n620));
  AO22X1 U226(.IN1(N1736),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n955),.Q(N1742));
  AO22X1 U227(.IN1(N1721),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n61),.Q(N1727));
  AO22X1 U228(.IN1(N1771),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n888),.Q(N1777));
  AO22X1 U229(.IN1(N460),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n811),.Q(n186));
  AO22X1 U230(.IN1(N359),.IN2(n130),.IN3(N349),.IN4(s_fract_48_i[41:41]),.Q(N365));
  HADDX1 U231(.A0(N400),.B0(\add_90_I9_L14036_C132/carry[4] ),.C1(\add_90_I9_L14036_C132/carry[5] ),.SO(N411));
  AO22X1 U232(.IN1(N394),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n914),.Q(N400));
  AO22X1 U233(.IN1(n459),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n831),.Q(n841));
  AO22X1 U234(.IN1(N1771),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n888),.Q(n918));
  AO22X1 U235(.IN1(N2279),.IN2(n123),.IN3(n1229),.IN4(n1077),.Q(N2285));
  AO22X1 U236(.IN1(N2264),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n917),.Q(n167));
  AO22X1 U237(.IN1(N2279),.IN2(n123),.IN3(n1229),.IN4(n1077),.Q(n895));
  AO22X1 U238(.IN1(N2199),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n199),.Q(N2205));
  AO22X1 U239(.IN1(N2233),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n200),.Q(n184));
  AO22X1 U240(.IN1(N2249),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n184),.Q(n828));
  AO22X1 U241(.IN1(n133),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n1078),.Q(n1047));
  AO22X1 U242(.IN1(N2187),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n1073),.Q(n977));
  AO22X1 U243(.IN1(N2203),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n977),.Q(n1019));
  HADDX1 U244(.A0(N1029),.B0(\add_90_I46_L14036_C132/carry[4] ),.C1(\add_90_I46_L14036_C132/carry[5] ),.SO(N1040));
  AO22X1 U245(.IN1(N887),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n929),.Q(n886));
  AO22X1 U246(.IN1(N888),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n936),.Q(N894));
  AO22X1 U247(.IN1(N2007),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n417),.Q(N2013));
  AO22X1 U248(.IN1(n867),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N2061),.Q(n915));
  AO22X1 U249(.IN1(n20),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1080),.Q(n1065));
  AO22X1 U250(.IN1(N681),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n976),.Q(N687));
  AO22X1 U251(.IN1(N817),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n357),.Q(N823));
  AO22X1 U252(.IN1(N800),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n835),.Q(n357));
  AO22X1 U253(.IN1(N801),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1083),.Q(N807));
  AO22X1 U254(.IN1(N886),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n169),.Q(n180));
  AO22X1 U255(.IN1(N887),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n929),.Q(N893));
  AO22X1 U256(.IN1(N803),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1051),.Q(n1005));
  AO22X1 U257(.IN1(N2008),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1082),.Q(n642));
  AO22X1 U258(.IN1(N2024),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n642),.Q(n972));
  AOI222X1 U259(.IN1(n369),.IN2(n819),.IN3(n1217),.IN4(n487),.IN5(n368),.IN6(N2126),.QN(n111));
  AO22X1 U260(.IN1(N1944),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n809),.Q(n188));
  AO22X1 U261(.IN1(N2025),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n30),.Q(n213));
  AO22X1 U262(.IN1(N1946),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n175),.Q(n195));
  AO22X1 U263(.IN1(N2059),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n995),.Q(n1052));
  AO22X1 U264(.IN1(N2043),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(N2033),.Q(n995));
  AO22X1 U265(.IN1(N612),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1068),.Q(n994));
  AO22X1 U266(.IN1(N630),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n404),.Q(n433));
  AO22X1 U267(.IN1(N835),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n382),.Q(n613));
  AO22X1 U268(.IN1(N818),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n432),.Q(n382));
  AO22X1 U269(.IN1(N495),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n1069),.Q(N501));
  HADDX1 U270(.A0(N638),.B0(\add_90_I23_L14036_C132/carry[4] ),.C1(\add_90_I23_L14036_C132/carry[5] ),.SO(N649));
  AO22X1 U271(.IN1(N768),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1063),.Q(n633));
  AO22X1 U272(.IN1(N718),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1018),.Q(N724));
  AO22X1 U273(.IN1(n470),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1084),.Q(n982));
  AO22X1 U274(.IN1(N1817),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1142),.Q(N1823));
  AO22X1 U275(.IN1(N1929),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n49),.Q(n658));
  AO22X1 U276(.IN1(N1866),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n16),.Q(N1872));
  AO22X1 U277(.IN1(N1930),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n26),.Q(n175));
  AOI222X1 U278(.IN1(n358),.IN2(n183),.IN3(n1289),.IN4(n1023),.IN5(n359),.IN6(n217),.QN(n129));
  AO22X1 U279(.IN1(N563),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n350),.Q(N569));
  AO22X1 U280(.IN1(N682),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n1064),.Q(n356));
  AO22X1 U281(.IN1(N699),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n356),.Q(n956));
  AO22X1 U282(.IN1(N614),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1110),.Q(n984));
  AO22X1 U283(.IN1(N666),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n59),.Q(n671));
  AO22X1 U284(.IN1(N564),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n572),.Q(n209));
  AO22X1 U285(.IN1(N513),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n1119),.Q(N519));
  AO22X1 U286(.IN1(N462),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n827),.Q(N468));
  AO22X1 U287(.IN1(N1832),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n833),.Q(n179));
  AO22X1 U288(.IN1(N1705),.IN2(n226),.IN3(n1227),.IN4(n1013),.Q(N1711));
  AO22X1 U289(.IN1(N1882),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n672),.Q(n187));
  AOI22X1 U290(.IN1(N1802),.IN2(n215),.IN3(n1211),.IN4(n1040),.QN(n1046));
  AO22X1 U291(.IN1(N1818),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1092),.Q(n891));
  AO22X1 U292(.IN1(N1770),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n912),.Q(n951));
  AO22X1 U293(.IN1(N527),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1074),.Q(n1081));
  AO22X1 U294(.IN1(N494),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n894),.Q(n202));
  AO22X1 U295(.IN1(N393),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n58),.Q(N399));
  AO22X1 U296(.IN1(N580),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n806),.Q(n486));
  AOI22X1 U297(.IN1(N597),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n486),.QN(n871));
  AO22X1 U298(.IN1(N444),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n830),.Q(n1007));
  AO22X1 U299(.IN1(N598),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1094),.Q(n983));
  AOI22X1 U300(.IN1(N581),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n209),.QN(n881));
  AO22X1 U301(.IN1(n458),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n937),.Q(n831));
  AO22X1 U302(.IN1(N412),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n907),.Q(n1032));
  AOI222X1 U303(.IN1(n344),.IN2(n620),.IN3(n1211),.IN4(n890),.IN5(n343),.IN6(n157),.QN(n100));
  AO22X1 U304(.IN1(n952),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1001),.Q(n955));
  AO22X1 U305(.IN1(N1721),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n61),.Q(n939));
  AO22X1 U306(.IN1(N1738),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n945),.Q(n176));
  AO22X1 U307(.IN1(N408),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n815),.Q(n1100));
  AO22X1 U308(.IN1(N426),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n735),.Q(N432));
  AO22X1 U309(.IN1(N393),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n58),.Q(n904));
  AO22X1 U310(.IN1(N410),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n904),.Q(n1066));
  AO22X1 U311(.IN1(N359),.IN2(n130),.IN3(N349),.IN4(s_fract_48_i[41:41]),.Q(n876));
  INVX0 U312(.INP(n1032),.ZN(n969));
  INVX0 U313(.INP(n1196),.ZN(n967));
  AOI22X1 U314(.IN1(n337),.IN2(n918),.IN3(n338),.IN4(n888),.QN(n1123));
  HADDX1 U315(.A0(\add_105_I47_L14036_C136/carry[4] ),.B0(N2336),.C1(\add_105_I47_L14036_C136/carry[5] ),.SO(N2346));
  AOI22X1 U316(.IN1(n21),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n926),.QN(n51));
  OAI22X2 U317(.IN1(n1139),.IN2(n1231),.IN3(n123),.IN4(n51),.QN(n52));
  AOI22X1 U318(.IN1(N1787),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n918),.QN(n57));
  AO22X1 U319(.IN1(N376),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n876),.Q(n58));
  AO22X2 U320(.IN1(N649),.IN2(n177),.IN3(n1289),.IN4(n1097),.Q(n59));
  AO22X1 U321(.IN1(N1705),.IN2(n226),.IN3(n1227),.IN4(n1013),.Q(n61));
  AO22X1 U322(.IN1(N2073),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n1086),.Q(n62));
  AO22X2 U323(.IN1(n4),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n990),.Q(n63));
  AO22X2 U324(.IN1(N394),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n914),.Q(n64));
  AO22X2 U325(.IN1(N375),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n911),.Q(n65));
  AO22X1 U326(.IN1(N785),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n633),.Q(n66));
  AO22X1 U327(.IN1(N972),.IN2(n227),.IN3(n1220),.IN4(n1115),.Q(n67));
  AO22X2 U328(.IN1(N1005),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n193),.Q(n70));
  AND2X1 U329(.IN1(n80),.IN2(n81),.Q(n515));
  AOI222X2 U330(.IN1(n344),.IN2(N1820),.IN3(n1211),.IN4(N1804),.IN5(n343),.IN6(N1836),.QN(n81));
  NAND2X0 U331(.IN1(n82),.IN2(n83),.QN(n721));
  AOI222X2 U332(.IN1(n586),.IN2(n1074),.IN3(n585),.IN4(n981),.IN5(n584),.IN6(n839),.QN(n83));
  AOI222X2 U333(.IN1(n624),.IN2(N1037),.IN3(n625),.IN4(N1009),.IN5(n626),.IN6(N1026),.QN(n1191));
  HADDX1 U334(.A0(N346),.B0(N347),.C1(\add_90_I6_L14036_C132/carry[2] ),.SO(N357));
  HADDX1 U335(.A0(N906),.B0(N907),.C1(\add_90_I39_L14036_C132/carry[2] ),.SO(N918));
  AO22X1 U336(.IN1(N901),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n216),.Q(N907));
  AO22X1 U337(.IN1(N374),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1104),.Q(n825));
  AO22X1 U338(.IN1(N374),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1104),.Q(N380));
  AO22X1 U339(.IN1(N442),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n821),.Q(n646));
  AO22X1 U340(.IN1(N442),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n821),.Q(N448));
  AO22X1 U341(.IN1(N476),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n713),.Q(N482));
  AO22X1 U342(.IN1(N476),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n713),.Q(n839));
  AO22X1 U343(.IN1(N680),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n507),.Q(n875));
  AO22X1 U377(.IN1(N680),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n507),.Q(N686));
  AO22X1 U378(.IN1(N697),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n875),.Q(n842));
  AO22X1 U386(.IN1(N697),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n875),.Q(N703));
  AO22X1 U388(.IN1(N714),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1003),.Q(n105));
  AO22X1 U390(.IN1(N714),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1003),.Q(N720));
  HADDX2 U392(.A0(N974),.B0(N975),.C1(\add_90_I43_L14036_C132/carry[2] ),.SO(N986));
  AOI222X1 U393(.IN1(n622),.IN2(n40),.IN3(n1225),.IN4(N958),.IN5(n623),.IN6(N992),.QN(n1192));
  AO22X1 U398(.IN1(N969),.IN2(n227),.IN3(n1221),.IN4(N958),.Q(N975));
  AO22X1 U400(.IN1(N1020),.IN2(n232),.IN3(s_fract_48_i[2:2]),.IN4(N1009),.Q(N1026));
  AND2X1 U402(.IN1(n84),.IN2(n85),.Q(n732));
  AOI221X2 U404(.IN1(n612),.IN2(n878),.IN3(n709),.IN4(n736),.IN5(n737),.QN(n84));
  AND2X1 U405(.IN1(n86),.IN2(n87),.Q(n710));
  AOI222X2 U451(.IN1(n622),.IN2(n934),.IN3(n1226),.IN4(n1090),.IN5(n623),.IN6(n1101),.QN(n87));
  AND2X1 U453(.IN1(n88),.IN2(n89),.Q(n697));
  AOI221X2 U455(.IN1(n1465),.IN2(n958),.IN3(n1464),.IN4(n701),.IN5(n702),.QN(n88));
  AOI222X1 U456(.IN1(n598),.IN2(n874),.IN3(n599),.IN4(n500),.IN5(n600),.IN6(n1004),.QN(n89));
  NAND3X1 U457(.IN1(n738),.IN2(n739),.IN3(n740),.QN(n736));
  AOI221X1 U506(.IN1(n1465),.IN2(n1070),.IN3(n673),.IN4(n1464),.IN5(n674),.QN(n92));
  HADDX2 U532(.A0(\add_90_I37_L14036_C132/carry[2] ),.B0(N874),.C1(\add_90_I37_L14036_C132/carry[3] ),.SO(N885));
  AO22X1 U536(.IN1(N767),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n989),.Q(n634));
  AO22X1 U537(.IN1(N869),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n840),.Q(n169));
  AO22X1 U538(.IN1(N869),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n840),.Q(N875));
  AO22X1 U539(.IN1(N459),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n863),.Q(N465));
  AO22X1 U543(.IN1(N868),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n864),.Q(N874));
  HADDX2 U544(.A0(N787),.B0(N788),.C1(\add_90_I32_L14036_C132/carry[2] ),.SO(N799));
  AO22X1 U545(.IN1(N782),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n1043),.Q(N788));
  AO22X1 U546(.IN1(N698),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n1004),.Q(N704));
  AO22X1 U551(.IN1(N698),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n1004),.Q(n500));
  AOI22X1 U552(.IN1(N919),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n239),.QN(n159));
  HADDX1 U554(.A0(\add_90_I14_L14036_C132/carry[2] ),.B0(N483),.C1(\add_90_I14_L14036_C132/carry[3] ),.SO(N494));
  HADDX1 U555(.A0(\add_90_I33_L14036_C132/carry[2] ),.B0(N806),.C1(\add_90_I33_L14036_C132/carry[3] ),.SO(N817));
  AO22X1 U556(.IN1(N800),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n835),.Q(N806));
  HADDX2 U564(.A0(\add_90_I41_L14036_C132/carry[2] ),.B0(N942),.C1(\add_90_I41_L14036_C132/carry[3] ),.SO(N953));
  AO22X1 U568(.IN1(N799),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n902),.Q(n804));
  AO22X1 U569(.IN1(N799),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n902),.Q(N805));
  AO22X1 U572(.IN1(N765),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n997),.Q(n1043));
  AO22X1 U573(.IN1(N765),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n997),.Q(N771));
  AO22X1 U577(.IN1(N425),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1100),.Q(N431));
  HADDX2 U578(.A0(N2300),.B0(N2301),.C1(\add_105_I45_L14036_C136/carry[2] ),.SO(N2311));
  AOI222X1 U579(.IN1(n1336),.IN2(N2359),.IN3(n385),.IN4(n42),.IN5(n386),.IN6(n41),.QN(n95));
  AND2X1 U591(.IN1(n90),.IN2(n91),.Q(n681));
  AOI222X1 U592(.IN1(n624),.IN2(N1039),.IN3(n625),.IN4(n70),.IN5(n626),.IN6(N1028),.QN(n90));
  AOI222X2 U595(.IN1(n622),.IN2(n1008),.IN3(n1224),.IN4(n860),.IN5(n623),.IN6(n193),.QN(n91));
  HADDX2 U596(.A0(N2332),.B0(N2333),.C1(\add_105_I47_L14036_C136/carry[2] ),.SO(N2343));
  AND2X1 U600(.IN1(n92),.IN2(n93),.Q(n669));
  AOI222X2 U601(.IN1(n598),.IN2(n1067),.IN3(n599),.IN4(n956),.IN5(n600),.IN6(n356),.QN(n93));
  AOI221X1 U602(.IN1(n347),.IN2(n925),.IN3(n489),.IN4(n429),.IN5(n490),.QN(n99));
  AOI22X1 U603(.IN1(N1789),.IN2(n1501),.IN3(n1500),.IN4(n94),.QN(n485));
  NAND2X0 U604(.IN1(n100),.IN2(n99),.QN(n94));
  AND2X1 U605(.IN1(n95),.IN2(n96),.Q(n506));
  AOI222X1 U607(.IN1(n383),.IN2(n896),.IN3(n1230),.IN4(n895),.IN5(n384),.IN6(n8),.QN(n96));
  AND2X1 U608(.IN1(n97),.IN2(n98),.Q(n497));
  AOI221X2 U616(.IN1(n372),.IN2(n699),.IN3(n442),.IN4(n501),.IN5(n502),.QN(n97));
  AOI222X2 U617(.IN1(n369),.IN2(n813),.IN3(n1217),.IN4(n965),.IN5(n368),.IN6(n978),.QN(n98));
  AO22X1 U619(.IN1(N479),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n938),.Q(N485));
  AO22X1 U620(.IN1(N391),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n825),.Q(N397));
  AO22X1 U622(.IN1(N663),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1020),.Q(n507));
  AO22X1 U623(.IN1(N376),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n876),.Q(N382));
  AO22X1 U625(.IN1(N785),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n633),.Q(N791));
  HADDX2 U631(.A0(\add_90_I41_L14036_C132/carry[4] ),.B0(N944),.C1(\add_90_I41_L14036_C132/carry[5] ),.SO(N955));
  AO22X1 U632(.IN1(N819),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n381),.Q(N825));
  AO22X1 U633(.IN1(N819),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n381),.Q(n478));
  OAI221X1 U634(.IN1(n643),.IN2(n592),.IN3(n1062),.IN4(n593),.IN5(n644),.QN(n102));
  HADDX2 U636(.A0(\add_90_I36_L14036_C132/carry[2] ),.B0(N857),.C1(\add_90_I36_L14036_C132/carry[3] ),.SO(N868));
  HADDX2 U641(.A0(N549),.B0(N550),.C1(\add_90_I18_L14036_C132/carry[2] ),.SO(N561));
  AO22X1 U642(.IN1(N561),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n921),.Q(n834));
  AO22X1 U644(.IN1(N561),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n921),.Q(N567));
  HADDX1 U647(.A0(\add_90_I31_L14036_C132/carry[3] ),.B0(N773),.C1(\add_90_I31_L14036_C132/carry[4] ),.SO(N784));
  AO22X1 U648(.IN1(N767),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n989),.Q(N773));
  AO22X1 U653(.IN1(N853),.IN2(n215),.IN3(n1210),.IN4(n1088),.Q(N859));
  HADDX1 U657(.A0(N842),.B0(\add_90_I35_L14036_C132/carry[4] ),.C1(\add_90_I35_L14036_C132/carry[5] ),.SO(N853));
  OAI21X1 U658(.IN1(n101),.IN2(n102),.IN3(n696),.QN(n637));
  OAI222X1 U680(.IN1(n881),.IN2(n630),.IN3(n1319),.IN4(n631),.IN5(n1039),.IN6(n632),.QN(n101));
  HADDX1 U692(.A0(\add_90_I34_L14036_C132/carry[3] ),.B0(N824),.C1(\add_90_I34_L14036_C132/carry[4] ),.SO(N835));
  AO22X1 U698(.IN1(N818),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n432),.Q(N824));
  HADDX2 U699(.A0(N872),.B0(N873),.C1(\add_90_I37_L14036_C132/carry[2] ),.SO(N884));
  HADDX2 U700(.A0(\add_90_I38_L14036_C132/carry[2] ),.B0(N891),.C1(\add_90_I38_L14036_C132/carry[3] ),.SO(N902));
  HADDX2 U701(.A0(\add_90_I39_L14036_C132/carry[4] ),.B0(N910),.C1(\add_90_I39_L14036_C132/carry[5] ),.SO(N921));
  HADDX2 U702(.A0(N413),.B0(N414),.C1(\add_90_I10_L14036_C132/carry[2] ),.SO(N425));
  HADDX2 U704(.A0(N583),.B0(N584),.C1(\add_90_I20_L14036_C132/carry[2] ),.SO(N595));
  AO22X1 U705(.IN1(N409),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n1120),.Q(N415));
  AO22X1 U706(.IN1(N904),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n1095),.Q(N910));
  HADDX1 U707(.A0(\add_90_I22_L14036_C132/carry[3] ),.B0(N620),.C1(\add_90_I22_L14036_C132/carry[4] ),.SO(N631));
  AO22X1 U709(.IN1(N614),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1110),.Q(N620));
  HADDX2 U710(.A0(N532),.B0(N533),.C1(\add_90_I17_L14036_C132/carry[2] ),.SO(N544));
  HADDX2 U711(.A0(\add_90_I23_L14036_C132/carry[3] ),.B0(N637),.C1(\add_90_I23_L14036_C132/carry[4] ),.SO(N648));
  AO22X1 U712(.IN1(N631),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n984),.Q(N637));
  AO22X1 U713(.IN1(N494),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n894),.Q(N500));
  AO22X1 U714(.IN1(N817),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n357),.Q(n336));
  AO22X1 U716(.IN1(N699),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n356),.Q(N705));
  AO22X1 U718(.IN1(N835),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n382),.Q(N841));
  AO22X1 U720(.IN1(N528),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n931),.Q(N534));
  AO22X1 U722(.IN1(N630),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n404),.Q(N636));
  HADDX1 U723(.A0(\add_90_I22_L14036_C132/carry[2] ),.B0(N619),.C1(\add_90_I22_L14036_C132/carry[3] ),.SO(N630));
  AO22X1 U724(.IN1(N562),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n908),.Q(N568));
  AO22X1 U725(.IN1(N613),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1028),.Q(N619));
  HADDX2 U726(.A0(\add_90_I21_L14036_C132/carry[2] ),.B0(N602),.C1(\add_90_I21_L14036_C132/carry[3] ),.SO(N613));
  AO22X1 U728(.IN1(N2280),.IN2(n123),.IN3(n1231),.IN4(N2270),.Q(n103));
  AO22X1 U729(.IN1(N2231),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n479),.Q(n104));
  AOI22X1 U730(.IN1(N921),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n1124),.QN(n1053));
  AO22X1 U731(.IN1(N921),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n1124),.Q(N927));
  HADDX2 U732(.A0(\add_90_I33_L14036_C132/carry[4] ),.B0(N808),.C1(\add_90_I33_L14036_C132/carry[5] ),.SO(N819));
  HADDX2 U734(.A0(N515),.B0(N516),.C1(\add_90_I16_L14036_C132/carry[2] ),.SO(N527));
  AO22X1 U735(.IN1(N802),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n66),.Q(n381));
  AO22X1 U736(.IN1(N802),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n66),.Q(N808));
  AOI22X1 U737(.IN1(N938),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1109),.QN(n1099));
  AO22X2 U738(.IN1(N1003),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(N992),.Q(N1009));
  HADDX2 U740(.A0(N957),.B0(N958),.C1(\add_90_I42_L14036_C132/carry[2] ),.SO(N969));
  AO22X1 U741(.IN1(N461),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1007),.Q(N467));
  AO22X1 U742(.IN1(N580),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n806),.Q(N586));
  AO22X1 U743(.IN1(N938),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1109),.Q(N944));
  HADDX2 U746(.A0(N991),.B0(N992),.C1(\add_90_I44_L14036_C132/carry[2] ),.SO(N1003));
  HADDX2 U747(.A0(N1008),.B0(N1009),.C1(\add_90_I45_L14036_C132/carry[2] ),.SO(N1020));
  AO22X1 U748(.IN1(N410),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n904),.Q(N416));
  HADDX1 U749(.A0(\add_90_I9_L14036_C132/carry[3] ),.B0(N399),.C1(\add_90_I9_L14036_C132/carry[4] ),.SO(N410));
  AO22X1 U750(.IN1(N581),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n209),.Q(N587));
  AO22X1 U752(.IN1(N426),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n735),.Q(n242));
  AO22X1 U753(.IN1(N460),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n811),.Q(N466));
  AO22X1 U754(.IN1(N598),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1094),.Q(N604));
  AO22X1 U755(.IN1(N511),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n202),.Q(N517));
  HADDX1 U758(.A0(\add_90_I15_L14036_C132/carry[2] ),.B0(N500),.C1(\add_90_I15_L14036_C132/carry[3] ),.SO(N511));
  HADDX2 U759(.A0(\add_90_I25_L14036_C132/carry[2] ),.B0(N670),.C1(\add_90_I25_L14036_C132/carry[3] ),.SO(N681));
  AO22X1 U760(.IN1(N564),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n572),.Q(N570));
  AO22X1 U761(.IN1(N666),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n59),.Q(N672));
  AO22X1 U764(.IN1(N936),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1055),.Q(N942));
  AO22X1 U766(.IN1(N700),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n987),.Q(N706));
  AO22X1 U770(.IN1(N768),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1063),.Q(N774));
  AO22X1 U771(.IN1(N2313),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n314),.Q(N2319));
  AO22X1 U772(.IN1(N445),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n1006),.Q(N451));
  AO22X1 U773(.IN1(N512),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n597),.Q(N518));
  HADDX2 U774(.A0(\add_105_I44_L14036_C136/carry[2] ),.B0(N2286),.C1(\add_105_I44_L14036_C136/carry[3] ),.SO(N2296));
  AO22X1 U776(.IN1(N2231),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n479),.Q(N2237));
  AO22X1 U777(.IN1(N2296),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n103),.Q(N2302));
  HADDX2 U778(.A0(\add_105_I43_L14036_C136/carry[2] ),.B0(n167),.C1(\add_105_I43_L14036_C136/carry[3] ),.SO(N2280));
  AO22X1 U779(.IN1(N2056),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n205),.Q(n191));
  AO22X1 U780(.IN1(N411),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n64),.Q(N417));
  AO22X1 U782(.IN1(N496),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n944),.Q(N502));
  AO22X1 U783(.IN1(N392),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n65),.Q(N398));
  AO22X1 U784(.IN1(N902),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n848),.Q(N908));
  AO22X1 U785(.IN1(N595),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n930),.Q(N601));
  AO22X1 U788(.IN1(N510),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n981),.Q(N516));
  AO22X1 U790(.IN1(N579),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n451),.Q(N585));
  AO22X1 U794(.IN1(N766),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n657),.Q(N772));
  AO22X2 U795(.IN1(N2247),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N2237),.Q(n107));
  HADDX2 U796(.A0(N2236),.B0(n104),.C1(\add_105_I41_L14036_C136/carry[2] ),.SO(N2247));
  AO22X1 U797(.IN1(N2247),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N2237),.Q(N2253));
  AO22X1 U798(.IN1(N2040),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n972),.Q(N2046));
  AND2X1 U800(.IN1(n108),.IN2(n109),.Q(n477));
  AOI222X1 U801(.IN1(n1336),.IN2(N2360),.IN3(n385),.IN4(n892),.IN5(n386),.IN6(N2350),.QN(n108));
  AND2X1 U802(.IN1(n110),.IN2(n111),.Q(n468));
  AOI221X2 U803(.IN1(n372),.IN2(n723),.IN3(n442),.IN4(n472),.IN5(n473),.QN(n110));
  AND2X1 U804(.IN1(n112),.IN2(n113),.Q(n643));
  AOI221X2 U806(.IN1(n1465),.IN2(n1121),.IN3(n1464),.IN4(n647),.IN5(n648),.QN(n112));
  AOI222X1 U807(.IN1(n598),.IN2(n1072),.IN3(n599),.IN4(n992),.IN5(n600),.IN6(n987),.QN(n113));
  AOI221X1 U808(.IN1(n347),.IN2(n887),.IN3(n460),.IN4(n429),.IN5(n461),.QN(n124));
  AND2X1 U809(.IN1(n114),.IN2(n115),.Q(n443));
  AOI222X1 U812(.IN1(n1336),.IN2(N2361),.IN3(n385),.IN4(n11),.IN5(n386),.IN6(N2351),.QN(n114));
  AND2X1 U813(.IN1(n116),.IN2(n117),.Q(n430));
  AOI222X2 U814(.IN1(n358),.IN2(n30),.IN3(n1289),.IN4(n1071),.IN5(n359),.IN6(n213),.QN(n117));
  AND2X1 U815(.IN1(n120),.IN2(n121),.Q(n655));
  AOI222X2 U818(.IN1(N1040),.IN2(n624),.IN3(n625),.IN4(n1126),.IN5(n626),.IN6(n1048),.QN(n120));
  AOI222X2 U819(.IN1(n622),.IN2(n67),.IN3(n1225),.IN4(n1115),.IN5(n623),.IN6(n165),.QN(n121));
  AO22X1 U820(.IN1(N833),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n44),.Q(N839));
  AO22X1 U821(.IN1(N867),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n45),.Q(N873));
  AND2X1 U822(.IN1(n124),.IN2(n125),.Q(n457));
  AOI222X2 U824(.IN1(n344),.IN2(n833),.IN3(n1210),.IN4(n1143),.IN5(n343),.IN6(n179),.QN(n125));
  HADDX1 U825(.A0(N2352),.B0(\add_105_I48_L14036_C136/carry[4] ),.C1(\add_105_I48_L14036_C136/carry[5] ),.SO(N2362));
  AO22X1 U826(.IN1(N358),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n838),.Q(N364));
  HADDX1 U830(.A0(\add_90_I45_L14036_C132/carry[4] ),.B0(N1012),.C1(\add_90_I45_L14036_C132/carry[5] ),.SO(N1023));
  AO22X1 U831(.IN1(N1004),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n1101),.Q(N1010));
  HADDX2 U832(.A0(N923),.B0(N924),.C1(\add_90_I40_L14036_C132/carry[2] ),.SO(N935));
  AND2X1 U833(.IN1(n126),.IN2(n127),.Q(n414));
  AOI222X2 U837(.IN1(n1336),.IN2(N2362),.IN3(n385),.IN4(n991),.IN5(n386),.IN6(n903),.QN(n126));
  AOI222X2 U838(.IN1(n383),.IN2(n63),.IN3(n1229),.IN4(n990),.IN5(n384),.IN6(n950),.QN(n127));
  AND2X1 U842(.IN1(n128),.IN2(n129),.Q(n402));
  AOI221X2 U844(.IN1(n1454),.IN2(n33),.IN3(n1453),.IN4(n406),.IN5(n407),.QN(n128));
  AOI22X1 U845(.IN1(N633),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n982),.QN(n194));
  AO22X1 U846(.IN1(N718),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1018),.Q(n855));
  AO22X1 U848(.IN1(N1735),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n953),.Q(N1741));
  AO22X1 U849(.IN1(N2119),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n813),.Q(N2125));
  INVX0 U850(.INP(n573),.ZN(n1127));
  INVX0 U851(.INP(n574),.ZN(n968));
  AO221X1 U854(.IN1(n575),.IN2(n735),.IN3(n574),.IN4(n65),.IN5(n687),.Q(n686));
  AOI222X1 U855(.IN1(n825),.IN2(n574),.IN3(n815),.IN4(n577),.IN5(n1100),.IN6(n575),.QN(n719));
  AOI222X2 U856(.IN1(N379),.IN2(n574),.IN3(N396),.IN4(n577),.IN5(N413),.IN6(n575),.QN(n747));
  INVX0 U857(.INP(n575),.ZN(n970));
  INVX0 U858(.INP(n592),.ZN(n329));
  INVX0 U860(.INP(n351),.ZN(n1116));
  AO22X1 U862(.IN1(N2138),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n853),.Q(n1125));
  AO22X1 U866(.IN1(N2138),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n853),.Q(N2144));
  DELLN1X2 U867(.INP(N2122),.Z(n131));
  AO22X1 U868(.IN1(N2122),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n816),.Q(N2128));
  DELLN1X2 U869(.INP(N2234),.Z(n133));
  DELLN1X2 U870(.INP(N2202),.Z(n134));
  DELLN1X2 U872(.INP(N2042),.Z(n135));
  DELLN1X2 U873(.INP(N2282),.Z(n136));
  DELLN1X2 U874(.INP(N2218),.Z(n138));
  DELLN1X2 U875(.INP(N2154),.Z(n139));
  DELLN1X2 U878(.INP(N2170),.Z(n140));
  DELLN1X2 U879(.INP(N2090),.Z(n141));
  DELLN1X2 U880(.INP(N2106),.Z(n142));
  XNOR2X1 U881(.IN1(\add_90_I46_L14036_C132/carry[5] ),.IN2(n143),.Q(N1041));
  AOI22X1 U884(.IN1(N1024),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(n901),.QN(n143));
  HADDX2 U885(.A0(N383),.B0(\add_90_I8_L14036_C132/carry[4] ),.C1(\add_90_I8_L14036_C132/carry[5] ),.SO(N394));
  AO22X1 U886(.IN1(N377),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N366),.Q(N383));
  AOI22X1 U887(.IN1(N377),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N366),.QN(n241));
  DELLN2X2 U888(.INP(N343),.Z(n147));
  AO22X2 U890(.IN1(N2296),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n103),.Q(n148));
  AO22X1 U891(.IN1(N2106),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n872),.Q(N2112));
  AO22X1 U892(.IN1(n142),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n872),.Q(n816));
  HADDX2 U893(.A0(\add_105_I32_L14036_C136/carry[4] ),.B0(N2096),.C1(\add_105_I32_L14036_C136/carry[5] ),.SO(N2106));
  HADDX2 U896(.A0(\add_105_I21_L14036_C136/carry[4] ),.B0(N1920),.C1(\add_105_I21_L14036_C136/carry[5] ),.SO(N1930));
  HADDX2 U898(.A0(\add_105_I43_L14036_C136/carry[4] ),.B0(N2272),.C1(\add_105_I43_L14036_C136/carry[5] ),.SO(N2282));
  HADDX2 U899(.A0(\add_105_I22_L14036_C136/carry[3] ),.B0(N1935),.C1(\add_105_I22_L14036_C136/carry[4] ),.SO(N1945));
  AO22X1 U900(.IN1(N1848),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n179),.Q(n149));
  HADDX2 U902(.A0(\add_105_I45_L14036_C136/carry[4] ),.B0(N2304),.C1(\add_105_I45_L14036_C136/carry[5] ),.SO(N2314));
  HADDX2 U903(.A0(\add_105_I9_L14036_C136/carry[3] ),.B0(N1727),.C1(\add_105_I9_L14036_C136/carry[4] ),.SO(N1737));
  OAI21X1 U904(.IN1(n150),.IN2(n151),.IN3(n709),.QN(n604));
  OAI222X1 U906(.IN1(n1314),.IN2(n627),.IN3(n1313),.IN4(n628),.IN5(n1312),.IN6(n629),.QN(n150));
  OAI221X1 U908(.IN1(n615),.IN2(n616),.IN3(n1311),.IN4(n617),.IN5(n618),.QN(n151));
  HADDX2 U909(.A0(\add_90_I11_L14036_C132/carry[4] ),.B0(N434),.C1(\add_90_I11_L14036_C132/carry[5] ),.SO(N445));
  AO22X1 U910(.IN1(N395),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n1196),.Q(N401));
  AO22X1 U911(.IN1(N480),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n841),.Q(N486));
  AO22X1 U912(.IN1(n152),.IN2(N446),.IN3(s_fract_48_i[36:36]),.IN4(n937),.Q(N452));
  DELLN1X2 U914(.INP(N650),.Z(n161));
  AO22X1 U915(.IN1(n227),.IN2(n5),.IN3(n1223),.IN4(n1132),.Q(n163));
  AO22X2 U916(.IN1(n857),.IN2(n229),.IN3(N1666),.IN4(s_fract_48_i[4:4]),.Q(n1132));
  AO22X2 U917(.IN1(N989),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n67),.Q(n165));
  DELLN1X2 U918(.INP(N907),.Z(n166));
  HADDX2 U920(.A0(\add_105_I23_L14036_C136/carry[3] ),.B0(N1951),.C1(\add_105_I23_L14036_C136/carry[4] ),.SO(N1961));
  HADDX2 U921(.A0(\add_90_I14_L14036_C132/carry[4] ),.B0(N485),.C1(\add_90_I14_L14036_C132/carry[5] ),.SO(N496));
  HADDX2 U923(.A0(N940),.B0(N941),.C1(\add_90_I41_L14036_C132/carry[2] ),.SO(N952));
  HADDX2 U924(.A0(\add_105_I28_L14036_C136/carry[3] ),.B0(N2031),.C1(\add_105_I28_L14036_C136/carry[4] ),.SO(N2041));
  HADDX2 U926(.A0(\add_90_I36_L14036_C132/carry[3] ),.B0(N858),.C1(\add_90_I36_L14036_C132/carry[4] ),.SO(N869));
  AO22X1 U927(.IN1(N1722),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n898),.Q(n945));
  HADDX1 U928(.A0(\add_105_I12_L14036_C136/carry[4] ),.B0(N1776),.C1(\add_105_I12_L14036_C136/carry[5] ),.SO(N1786));
  AO22X1 U929(.IN1(n3),.IN2(n123),.IN3(n1230),.IN4(n1033),.Q(n178));
  AO22X2 U930(.IN1(N1816),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1143),.Q(n833));
  AOI22X2 U932(.IN1(N2263),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n107),.QN(n181));
  AO22X2 U934(.IN1(N2010),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1023),.Q(n183));
  AO22X1 U938(.IN1(N2217),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n868),.Q(n200));
  AO22X1 U939(.IN1(N2041),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n213),.Q(n185));
  AO22X1 U944(.IN1(N1866),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n16),.Q(n672));
  AO22X1 U949(.IN1(N1723),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1195),.Q(N1729));
  AO22X1 U953(.IN1(N1801),.IN2(n215),.IN3(n1211),.IN4(n1014),.Q(N1807));
  HADDX1 U954(.A0(\add_105_I12_L14036_C136/carry[3] ),.B0(N1775),.C1(\add_105_I12_L14036_C136/carry[4] ),.SO(N1785));
  AO22X1 U956(.IN1(N1945),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n658),.Q(n190));
  HADDX2 U957(.A0(\add_105_I13_L14036_C136/carry[3] ),.B0(N1791),.C1(\add_105_I13_L14036_C136/carry[4] ),.SO(N1801));
  XNOR2X2 U962(.IN1(n194),.IN2(\add_90_I23_L14036_C132/carry[5] ),.Q(N650));
  AO22X1 U963(.IN1(N429),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1032),.Q(N435));
  AO22X1 U964(.IN1(N2183),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n699),.Q(n199));
  AO22X1 U965(.IN1(N2201),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N2191),.Q(n868));
  XNOR2X2 U970(.IN1(n201),.IN2(\add_105_I14_L14036_C136/carry[5] ),.Q(N1819));
  OA22X1 U971(.IN1(n1209),.IN2(n1056),.IN3(n215),.IN4(n57),.Q(n201));
  AO22X1 U973(.IN1(N477),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n186),.Q(n894));
  AO22X1 U974(.IN1(N2040),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n972),.Q(n205));
  AO22X1 U975(.IN1(N1834),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n891),.Q(n207));
  XNOR2X1 U977(.IN1(\add_90_I37_L14036_C132/carry[5] ),.IN2(n211),.Q(N888));
  AOI22X1 U978(.IN1(N871),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1044),.QN(n211));
  AO22X1 U981(.IN1(N884),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n854),.Q(n216));
  XNOR2X2 U982(.IN1(n856),.IN2(\add_105_I33_L14036_C136/carry[5] ),.Q(N2123));
  XNOR2X2 U983(.IN1(n814),.IN2(\add_105_I39_L14036_C136/carry[5] ),.Q(N2219));
  XNOR2X1 U985(.IN1(\add_90_I32_L14036_C132/carry[5] ),.IN2(n218),.Q(N803));
  AOI22X1 U986(.IN1(N786),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n1022),.QN(n218));
  AO22X2 U987(.IN1(N1978),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n836),.Q(n219));
  XNOR2X2 U994(.IN1(N1793),.IN2(\add_105_I13_L14036_C136/carry[5] ),.Q(n1056));
  AO22X1 U995(.IN1(N834),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n900),.Q(n220));
  AO22X1 U997(.IN1(n499),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n942),.Q(n818));
  DELLN1X2 U1002(.INP(N905),.Z(n499));
  AO22X1 U1006(.IN1(n130),.IN2(N2267),.IN3(s_fract_48_i[41:41]),.IN4(n926),.Q(n228));
  DELLN1X2 U1007(.INP(N1742),.Z(n230));
  XNOR2X1 U1015(.IN1(n234),.IN2(\add_90_I40_L14036_C132/carry[5] ),.Q(N939));
  AOI22X1 U1016(.IN1(N922),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n818),.QN(n234));
  AO22X1 U1019(.IN1(N731),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n105),.Q(n237));
  HADDX2 U1020(.A0(N366),.B0(\add_90_I7_L14036_C132/carry[4] ),.C1(N378),.SO(N377));
  HADDX1 U1021(.A0(N382),.B0(\add_90_I8_L14036_C132/carry[3] ),.C1(\add_90_I8_L14036_C132/carry[4] ),.SO(N393));
  DELLN1X2 U1022(.INP(N908),.Z(n239));
  AO22X1 U1028(.IN1(n221),.IN2(N1784),.IN3(s_fract_48_i[11:11]),.IN4(n843),.Q(n240));
  AO22X1 U1029(.IN1(N1927),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n885),.Q(n243));
  AO22X1 U1036(.IN1(N1944),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n809),.Q(N1950));
  AO22X1 U1037(.IN1(N2200),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N2190),.Q(N2206));
  AO22X1 U1038(.IN1(N2200),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N2190),.Q(n823));
  AO22X1 U1043(.IN1(N1961),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n190),.Q(N1967));
  XNOR2X1 U1044(.IN1(n245),.IN2(\add_90_I39_L14036_C132/carry[5] ),.Q(N922));
  AOI22X1 U1045(.IN1(N905),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n942),.QN(n245));
  AO22X1 U1053(.IN1(N2024),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n642),.Q(N2030));
  DELLN2X2 U1054(.INP(N990),.Z(n313));
  AO22X1 U1055(.IN1(N2184),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n723),.Q(n689));
  HADDX2 U1056(.A0(\add_105_I44_L14036_C136/carry[3] ),.B0(N2287),.C1(\add_105_I44_L14036_C136/carry[4] ),.SO(N2297));
  AO22X1 U1060(.IN1(N2168),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n960),.Q(N2174));
  AO22X1 U1061(.IN1(N2168),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n960),.Q(n723));
  AOI221X1 U1063(.IN1(n329),.IN2(n330),.IN3(n986),.IN4(n1451),.IN5(n335),.QN(n590));
  NAND2X0 U1098(.IN1(n1180),.IN2(n1181),.QN(n330));
  AO22X2 U1101(.IN1(n923),.IN2(n1217),.IN3(n884),.IN4(n595),.Q(n335));
  AO22X1 U1104(.IN1(N633),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n982),.Q(n986));
  NAND2X0 U1105(.IN1(n766),.IN2(n592),.QN(n593));
  AO22X1 U1107(.IN1(N2297),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n178),.Q(N2303));
  DELLN1X2 U1108(.INP(N552),.Z(n350));
  AO22X1 U1110(.IN1(N990),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1079),.Q(N996));
  AO22X1 U1111(.IN1(n313),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1079),.Q(n893));
  DELLN2X2 U1112(.INP(N565),.Z(n353));
  AO22X1 U1113(.IN1(N2232),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(N2222),.Q(N2238));
  AO22X1 U1114(.IN1(N2217),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n868),.Q(N2223));
  HADDX2 U1115(.A0(\add_90_I25_L14036_C132/carry[3] ),.B0(N671),.C1(\add_90_I25_L14036_C132/carry[4] ),.SO(N682));
  HADDX2 U1117(.A0(\add_90_I32_L14036_C132/carry[2] ),.B0(N789),.C1(\add_90_I32_L14036_C132/carry[3] ),.SO(N800));
  XNOR2X1 U1118(.IN1(\add_90_I43_L14036_C132/carry[5] ),.IN2(n373),.Q(N990));
  AOI22X1 U1119(.IN1(N973),.IN2(n227),.IN3(n1223),.IN4(n974),.QN(n373));
  AO22X1 U1120(.IN1(N565),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n923),.Q(N571));
  AO22X1 U1121(.IN1(n353),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n923),.Q(n884));
  DELLN2X2 U1122(.INP(N769),.Z(n374));
  AO22X1 U1123(.IN1(N801),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1083),.Q(n432));
  XNOR2X1 U1124(.IN1(\add_105_I48_L14036_C136/carry[5] ),.IN2(n405),.Q(N2363));
  AOI22X1 U1125(.IN1(N2347),.IN2(n69),.IN3(n1205),.IN4(n31),.QN(n405));
  AO22X1 U1126(.IN1(N1881),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1140),.Q(N1887));
  AO22X1 U1128(.IN1(N1881),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1140),.Q(n1026));
  XNOR2X1 U1129(.IN1(\add_90_I18_L14036_C132/carry[5] ),.IN2(n416),.Q(N565));
  AOI22X1 U1131(.IN1(N548),.IN2(n164),.IN3(n1217),.IN4(n865),.QN(n416));
  HADDX1 U1132(.A0(\add_105_I10_L14036_C136/carry[3] ),.B0(N1743),.C1(\add_105_I10_L14036_C136/carry[4] ),.SO(N1753));
  AO22X1 U1133(.IN1(N1818),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1092),.Q(N1824));
  AO22X1 U1135(.IN1(N2136),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N2126),.Q(N2142));
  AO22X1 U1136(.IN1(N2136),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N2126),.Q(n877));
  AO22X1 U1137(.IN1(N1739),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n940),.Q(N1745));
  AO22X1 U1138(.IN1(N769),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1076),.Q(N775));
  AO22X1 U1139(.IN1(n374),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1076),.Q(n1022));
  AO22X1 U1140(.IN1(N1929),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n49),.Q(N1935));
  AO22X1 U1141(.IN1(N1991),.IN2(n177),.IN3(n1290),.IN4(n947),.Q(n417));
  AO22X1 U1143(.IN1(N2248),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n106),.Q(N2254));
  AO22X1 U1144(.IN1(N2248),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n106),.Q(n917));
  AO22X1 U1145(.IN1(N2137),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n1054),.Q(N2143));
  AO22X1 U1146(.IN1(N2137),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n1054),.Q(n909));
  AO22X1 U1147(.IN1(N2120),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n819),.Q(n812));
  AO22X1 U1150(.IN1(N2169),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(N2159),.Q(N2175));
  AO22X1 U1151(.IN1(N2169),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(N2159),.Q(n742));
  AO22X1 U1152(.IN1(N1833),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n810),.Q(N1839));
  AO22X1 U1153(.IN1(n50),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n810),.Q(n924));
  HADDX2 U1155(.A0(\add_105_I15_L14036_C136/carry[3] ),.B0(N1823),.C1(\add_105_I15_L14036_C136/carry[4] ),.SO(N1833));
  AO22X1 U1157(.IN1(N1928),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n27),.Q(N1934));
  AO22X1 U1158(.IN1(N1928),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n27),.Q(n809));
  XNOR2X1 U1159(.IN1(\add_90_I30_L14036_C132/carry[5] ),.IN2(n445),.Q(N769));
  AOI22X1 U1160(.IN1(N752),.IN2(n204),.IN3(n1214),.IN4(n824),.QN(n445));
  DELLN2X2 U1162(.INP(N1007),.Z(n446));
  AO22X1 U1164(.IN1(N1007),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n893),.Q(N1013));
  AO22X1 U1165(.IN1(n446),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n893),.Q(n901));
  AO22X1 U1166(.IN1(N1977),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n837),.Q(N1983));
  AO22X1 U1167(.IN1(N1977),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n837),.Q(n805));
  HADDX2 U1168(.A0(\add_90_I18_L14036_C132/carry[2] ),.B0(N551),.C1(\add_90_I18_L14036_C132/carry[3] ),.SO(N562));
  AO22X1 U1170(.IN1(N582),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n884),.Q(N588));
  AO22X1 U1171(.IN1(N1816),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1143),.Q(N1822));
  AO22X1 U1172(.IN1(N2104),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n487),.Q(N2110));
  AO22X1 U1175(.IN1(N2104),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n487),.Q(n819));
  AO22X1 U1176(.IN1(N684),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n1057),.Q(N690));
  AO22X1 U1177(.IN1(N684),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n1057),.Q(n1000));
  AO22X1 U1178(.IN1(N2330),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n950),.Q(N2336));
  AO22X1 U1179(.IN1(N2330),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n950),.Q(n991));
  AO22X1 U1180(.IN1(N497),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n861),.Q(N503));
  AO22X1 U1181(.IN1(N497),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n861),.Q(n889));
  AO22X1 U1182(.IN1(N2233),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n200),.Q(N2239));
  HADDX2 U1183(.A0(\add_105_I36_L14036_C136/carry[2] ),.B0(N2158),.C1(\add_105_I36_L14036_C136/carry[3] ),.SO(N2168));
  AO22X1 U1184(.IN1(N531),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n844),.Q(N537));
  AO22X1 U1185(.IN1(N531),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n844),.Q(n865));
  AO22X1 U1186(.IN1(N786),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n1022),.Q(N792));
  DELLN2X2 U1187(.INP(N446),.Z(n458));
  DELLN2X2 U1189(.INP(N463),.Z(n459));
  DELLN2X2 U1191(.INP(N616),.Z(n470));
  DELLN2X2 U1192(.INP(N820),.Z(n471));
  AO22X1 U1193(.IN1(N357),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(N347),.Q(N363));
  AO22X1 U1194(.IN1(N820),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n1005),.Q(N826));
  AO22X1 U1196(.IN1(N1768),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n916),.Q(N1774));
  HADDX2 U1197(.A0(N379),.B0(N380),.C1(\add_90_I8_L14036_C132/carry[2] ),.SO(N391));
  AO22X1 U1198(.IN1(N2215),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n846),.Q(n479));
  HADDX2 U1199(.A0(N804),.B0(N805),.C1(\add_90_I33_L14036_C132/carry[2] ),.SO(N816));
  AO22X1 U1200(.IN1(N563),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n350),.Q(n806));
  AO22X1 U1204(.IN1(N2249),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n184),.Q(N2255));
  HADDX2 U1205(.A0(\add_105_I42_L14036_C136/carry[2] ),.B0(N2254),.C1(\add_105_I42_L14036_C136/carry[3] ),.SO(N2264));
  HADDX2 U1207(.A0(N702),.B0(n842),.C1(\add_90_I27_L14036_C132/carry[2] ),.SO(N714));
  AO22X1 U1208(.IN1(N2265),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n828),.Q(N2271));
  AOI22X1 U1209(.IN1(N2265),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(n828),.QN(n959));
  HADDX2 U1211(.A0(\add_105_I42_L14036_C136/carry[3] ),.B0(N2255),.C1(\add_105_I42_L14036_C136/carry[4] ),.SO(N2265));
  AO22X1 U1212(.IN1(N2088),.IN2(n164),.IN3(n1217),.IN4(n132),.Q(n487));
  XNOR2X1 U1215(.IN1(n488),.IN2(\add_90_I33_L14036_C132/carry[5] ),.Q(N820));
  AOI22X1 U1216(.IN1(N803),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1051),.QN(n488));
  AO22X1 U1217(.IN1(N2105),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1011),.Q(N2111));
  AO22X1 U1218(.IN1(N2105),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1011),.Q(n817));
  HADDX2 U1219(.A0(\add_105_I46_L14036_C136/carry[4] ),.B0(N2320),.C1(\add_105_I46_L14036_C136/carry[5] ),.SO(N2330));
  HADDX2 U1220(.A0(N651),.B0(n851),.C1(\add_90_I24_L14036_C132/carry[2] ),.SO(N663));
  AOI22X1 U1221(.IN1(N2251),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1021),.QN(n508));
  HADDX2 U1222(.A0(\add_90_I39_L14036_C132/carry[2] ),.B0(N908),.C1(\add_90_I39_L14036_C132/carry[3] ),.SO(N919));
  AO22X1 U1223(.IN1(N2281),.IN2(n123),.IN3(n1230),.IN4(n1033),.Q(N2287));
  HADDX2 U1224(.A0(N566),.B0(N567),.C1(\add_90_I19_L14036_C132/carry[2] ),.SO(N578));
  HADDX2 U1226(.A0(\add_90_I19_L14036_C132/carry[2] ),.B0(N568),.C1(\add_90_I19_L14036_C132/carry[3] ),.SO(N579));
  HADDX2 U1227(.A0(N770),.B0(N771),.C1(\add_90_I31_L14036_C132/carry[2] ),.SO(N782));
  XNOR2X1 U1230(.IN1(n516),.IN2(\add_90_I38_L14036_C132/carry[5] ),.Q(N905));
  AOI22X1 U1231(.IN1(N888),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n936),.QN(n516));
  HADDX2 U1232(.A0(\add_90_I31_L14036_C132/carry[2] ),.B0(N772),.C1(\add_90_I31_L14036_C132/carry[3] ),.SO(N783));
  DELLN2X2 U1233(.INP(N514),.Z(n517));
  HADDX2 U1234(.A0(N617),.B0(N618),.C1(\add_90_I22_L14036_C132/carry[2] ),.SO(N629));
  DELLN1X2 U1237(.INP(N553),.Z(n572));
  AO22X1 U1238(.IN1(N514),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n889),.Q(N520));
  AO22X1 U1239(.IN1(N748),.IN2(n204),.IN3(n1214),.IN4(n237),.Q(N754));
  AO22X2 U1240(.IN1(N647),.IN2(n177),.IN3(n1289),.IN4(n433),.Q(n576));
  AO22X1 U1242(.IN1(N461),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1007),.Q(n591));
  OAI22X2 U1244(.IN1(n1056),.IN2(n1209),.IN3(n215),.IN4(n57),.QN(n594));
  XNOR2X1 U1245(.IN1(\add_90_I42_L14036_C132/carry[5] ),.IN2(n596),.Q(N973));
  AOI22X1 U1247(.IN1(N956),.IN2(n226),.IN3(n1224),.IN4(n1027),.QN(n596));
  AO22X2 U1248(.IN1(N495),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n1069),.Q(n597));
  XNOR2X1 U1249(.IN1(n614),.IN2(\add_90_I29_L14036_C132/carry[5] ),.Q(N752));
  AOI22X1 U1251(.IN1(N735),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n946),.QN(n614));
  AOI22X1 U1252(.IN1(N2299),.IN2(n122),.IN3(s_fract_48_i[43:43]),.IN4(n52),.QN(n962));
  AO22X1 U1254(.IN1(N2185),.IN2(n152),.IN3(s_fract_48_i[36:36]),.IN4(n742),.Q(n621));
  XOR2X1 U1255(.IN1(\add_105_I9_L14036_C136/carry[5] ),.IN2(N1729),.Q(N1739));
  HADDX2 U1256(.A0(\add_90_I30_L14036_C132/carry[4] ),.B0(N757),.C1(\add_90_I30_L14036_C132/carry[5] ),.SO(N768));
  AO22X1 U1257(.IN1(n22),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n940),.Q(n935));
  HADDX2 U1258(.A0(\add_90_I30_L14036_C132/carry[3] ),.B0(N756),.C1(\add_90_I30_L14036_C132/carry[4] ),.SO(N767));
  XNOR2X1 U1259(.IN1(n641),.IN2(\add_90_I36_L14036_C132/carry[5] ),.Q(N871));
  AOI22X1 U1260(.IN1(N854),.IN2(n215),.IN3(n1211),.IN4(n1002),.QN(n641));
  HADDX2 U1261(.A0(\add_105_I26_L14036_C136/carry[2] ),.B0(N1998),.C1(\add_105_I26_L14036_C136/carry[3] ),.SO(N2008));
  HADDX1 U1262(.A0(\add_105_I18_L14036_C136/carry[4] ),.B0(N1872),.C1(\add_105_I18_L14036_C136/carry[5] ),.SO(N1882));
  DELLN1X2 U1263(.INP(N755),.Z(n657));
  HADDX2 U1264(.A0(N753),.B0(N754),.C1(\add_90_I30_L14036_C132/carry[2] ),.SO(N765));
  HADDX2 U1267(.A0(\add_90_I24_L14036_C132/carry[4] ),.B0(N655),.C1(\add_90_I24_L14036_C132/carry[5] ),.SO(N666));
  HADDX2 U1269(.A0(N481),.B0(N482),.C1(\add_90_I14_L14036_C132/carry[2] ),.SO(N493));
  AO22X2 U1273(.IN1(N1976),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1059),.Q(n683));
  AOI22X1 U1275(.IN1(N837),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1012),.QN(n684));
  XNOR2X1 U1277(.IN1(\add_105_I32_L14036_C136/carry[5] ),.IN2(n688),.Q(N2107));
  AOI22X1 U1279(.IN1(N2091),.IN2(n164),.IN3(n1216),.IN4(N2081),.QN(n688));
  AO22X1 U1280(.IN1(N2167),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n829),.Q(n699));
  AO22X1 U1281(.IN1(N2153),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n909),.Q(n712));
  AO22X2 U1282(.IN1(N459),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n863),.Q(n713));
  HADDX2 U1284(.A0(N447),.B0(n646),.C1(\add_90_I12_L14036_C132/carry[2] ),.SO(N459));
  XNOR2X1 U1285(.IN1(\add_90_I41_L14036_C132/carry[5] ),.IN2(n722),.Q(N956));
  AOI22X1 U1286(.IN1(N939),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1009),.QN(n722));
  HADDX1 U1288(.A0(N348),.B0(\add_90_I6_L14036_C132/carry[2] ),.C1(\add_90_I6_L14036_C132/carry[3] ),.SO(N358));
  HADDX2 U1290(.A0(\add_105_I25_L14036_C136/carry[4] ),.B0(N1984),.C1(\add_105_I25_L14036_C136/carry[5] ),.SO(N1994));
  XNOR2X1 U1291(.IN1(\add_105_I20_L14036_C136/carry[5] ),.IN2(n734),.Q(N1915));
  AOI22X1 U1293(.IN1(N1899),.IN2(n204),.IN3(n1213),.IN4(n1025),.QN(n734));
  AO22X2 U1296(.IN1(N409),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n1120),.Q(n735));
  HADDX2 U1298(.A0(\add_90_I9_L14036_C132/carry[2] ),.B0(N398),.C1(\add_90_I9_L14036_C132/carry[3] ),.SO(N409));
  XOR2X1 U1299(.IN1(\add_90_I11_L14036_C132/carry[5] ),.IN2(N435),.Q(N446));
  DELLN1X2 U1300(.INP(N874),.Z(n743));
  HADDX2 U1301(.A0(\add_90_I18_L14036_C132/carry[3] ),.B0(N552),.C1(\add_90_I18_L14036_C132/carry[4] ),.SO(N563));
  XNOR2X1 U1303(.IN1(n808),.IN2(\add_105_I29_L14036_C136/carry[5] ),.Q(N2059));
  AOI22X1 U1304(.IN1(N2043),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(N2033),.QN(n808));
  AO22X1 U1305(.IN1(N885),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n743),.Q(N891));
  AO22X2 U1307(.IN1(N989),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n67),.Q(N995));
  DELLN1X2 U1350(.INP(N449),.Z(n811));
  AO22X1 U1352(.IN1(N2103),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n965),.Q(n813));
  AOI22X1 U1353(.IN1(N2203),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n977),.QN(n814));
  HADDX2 U1354(.A0(\add_105_I27_L14036_C136/carry[2] ),.B0(N2014),.C1(\add_105_I27_L14036_C136/carry[3] ),.SO(N2024));
  AO22X1 U1355(.IN1(N391),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n825),.Q(n815));
  HADDX2 U1356(.A0(\add_105_I37_L14036_C136/carry[2] ),.B0(N2174),.C1(\add_105_I37_L14036_C136/carry[3] ),.SO(N2184));
  HADDX2 U1357(.A0(N838),.B0(N839),.C1(\add_90_I35_L14036_C132/carry[2] ),.SO(N850));
  AO22X1 U1358(.IN1(N2139),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N2129),.Q(N2145));
  AO22X1 U1359(.IN1(n25),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(N2129),.Q(n1016));
  AO22X1 U1360(.IN1(N1006),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n165),.Q(N1012));
  AO22X1 U1361(.IN1(N2089),.IN2(n164),.IN3(n1217),.IN4(n62),.Q(n1011));
  HADDX2 U1362(.A0(N821),.B0(N822),.C1(\add_90_I34_L14036_C132/carry[2] ),.SO(N833));
  AO22X2 U1363(.IN1(N528),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n931),.Q(n820));
  HADDX2 U1364(.A0(\add_90_I16_L14036_C132/carry[2] ),.B0(N517),.C1(\add_90_I16_L14036_C132/carry[3] ),.SO(N528));
  AO22X1 U1365(.IN1(N425),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1100),.Q(n821));
  XNOR2X1 U1366(.IN1(\add_105_I34_L14036_C136/carry[5] ),.IN2(n822),.Q(N2139));
  AOI22X1 U1367(.IN1(N2123),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n1065),.QN(n822));
  AO22X1 U1368(.IN1(N2027),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n1089),.Q(n1038));
  AO22X2 U1369(.IN1(N735),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n946),.Q(n824));
  HADDX2 U1370(.A0(N362),.B0(N363),.C1(\add_90_I7_L14036_C132/carry[2] ),.SO(N374));
  XOR2X1 U1371(.IN1(\add_90_I15_L14036_C132/carry[5] ),.IN2(N503),.Q(N514));
  XNOR2X1 U1372(.IN1(\add_105_I27_L14036_C136/carry[5] ),.IN2(n826),.Q(N2027));
  AOI22X1 U1373(.IN1(N2011),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1030),.QN(n826));
  DELLN1X2 U1374(.INP(N451),.Z(n827));
  AO22X1 U1375(.IN1(N1851),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1010),.Q(N1857));
  AO22X1 U1376(.IN1(n23),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n1010),.Q(n919));
  AO22X1 U1377(.IN1(N2151),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n973),.Q(n829));
  AO22X1 U1378(.IN1(N427),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1066),.Q(n830));
  HADDX1 U1379(.A0(\add_90_I10_L14036_C132/carry[3] ),.B0(N416),.C1(\add_90_I10_L14036_C132/carry[4] ),.SO(N427));
  AO22X1 U1380(.IN1(n221),.IN2(N1787),.IN3(s_fract_48_i[11:11]),.IN4(n918),.Q(N1793));
  DELLN2X2 U1381(.INP(N2347),.Z(n832));
  DELLN1X2 U1382(.INP(N789),.Z(n835));
  DELLN1X2 U1383(.INP(N1968),.Z(n836));
  DELLN1X2 U1384(.INP(N1967),.Z(n837));
  AO22X1 U1385(.IN1(n147),.IN2(n123),.IN3(n1228),.IN4(N334),.Q(n838));
  HADDX2 U1386(.A0(N464),.B0(N465),.C1(\add_90_I13_L14036_C132/carry[2] ),.SO(N476));
  AO22X1 U1387(.IN1(N919),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n239),.Q(N925));
  DELLN1X2 U1388(.INP(N858),.Z(n840));
  HADDX2 U1389(.A0(\add_90_I30_L14036_C132/carry[2] ),.B0(N755),.C1(\add_90_I30_L14036_C132/carry[3] ),.SO(N766));
  HADDX2 U1390(.A0(\add_90_I26_L14036_C132/carry[2] ),.B0(N687),.C1(\add_90_I26_L14036_C132/carry[3] ),.SO(N698));
  AO22X1 U1391(.IN1(N903),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n180),.Q(N909));
  HADDX2 U1392(.A0(N685),.B0(N686),.C1(\add_90_I26_L14036_C132/carry[2] ),.SO(N697));
  DELLN1X2 U1393(.INP(N1774),.Z(n843));
  HADDX2 U1394(.A0(N889),.B0(N890),.C1(\add_90_I38_L14036_C132/carry[2] ),.SO(N901));
  AO22X1 U1395(.IN1(n517),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n889),.Q(n844));
  AO22X1 U1396(.IN1(n832),.IN2(n69),.IN3(n1205),.IN4(n31),.Q(n845));
  DELLN1X2 U1397(.INP(N2205),.Z(n846));
  DELLN1X2 U1398(.INP(N909),.Z(n847));
  DELLN1X2 U1399(.INP(N891),.Z(n848));
  AO22X1 U1400(.IN1(N1024),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(n901),.Q(n849));
  HADDX2 U1401(.A0(\add_90_I38_L14036_C132/carry[3] ),.B0(N892),.C1(\add_90_I38_L14036_C132/carry[4] ),.SO(N903));
  DELLN1X2 U1402(.INP(N432),.Z(n850));
  AO22X1 U1403(.IN1(N646),.IN2(n177),.IN3(n1289),.IN4(n899),.Q(n851));
  DELLN1X2 U1404(.INP(N1741),.Z(n852));
  DELLN1X2 U1405(.INP(N873),.Z(n854));
  AO22X1 U1406(.IN1(n210),.IN2(N1849),.IN3(s_fract_48_i[15:15]),.IN4(n924),.Q(N1855));
  HADDX2 U1407(.A0(N2220),.B0(N2221),.C1(\add_105_I40_L14036_C136/carry[2] ),.SO(N2231));
  AO22X1 U1408(.IN1(N647),.IN2(n177),.IN3(n1289),.IN4(n433),.Q(N653));
  HADDX2 U1409(.A0(\add_90_I23_L14036_C132/carry[2] ),.B0(N636),.C1(\add_90_I23_L14036_C132/carry[3] ),.SO(N647));
  AOI22X1 U1410(.IN1(N2107),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1080),.QN(n856));
  AO22X1 U1411(.IN1(N2010),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1023),.Q(N2016));
  AO22X1 U1412(.IN1(N2009),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1071),.Q(N2015));
  HADDX2 U1413(.A0(N2188),.B0(N2189),.C1(\add_105_I38_L14036_C136/carry[2] ),.SO(N2199));
  NAND3X1 U1414(.IN1(n504),.IN2(n503),.IN3(n505),.QN(n501));
  HADDX2 U1415(.A0(N2204),.B0(N2205),.C1(\add_105_I39_L14036_C136/carry[2] ),.SO(N2215));
  AO22X1 U1416(.IN1(N1848),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n179),.Q(N1854));
  AO22X1 U1417(.IN1(N1819),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n594),.Q(N1825));
  AO22X1 U1418(.IN1(N1819),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n594),.Q(n913));
  AO22X1 U1419(.IN1(N1752),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n230),.Q(N1758));
  DELLN2X2 U1420(.INP(N1674),.Z(n857));
  DELLN1X2 U1421(.INP(N1704),.Z(n858));
  HADDX2 U1422(.A0(N2156),.B0(N2157),.C1(\add_105_I36_L14036_C136/carry[2] ),.SO(N2167));
  HADDX2 U1423(.A0(N2172),.B0(N2173),.C1(\add_105_I37_L14036_C136/carry[2] ),.SO(N2183));
  DELLN1X2 U1424(.INP(N2135),.Z(n859));
  DELLN1X2 U1425(.INP(N960),.Z(n860));
  AO22X1 U1426(.IN1(N954),.IN2(n226),.IN3(n1226),.IN4(n1096),.Q(N960));
  AO22X1 U1427(.IN1(N2135),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n978),.Q(N2141));
  AO22X1 U1428(.IN1(n859),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n978),.Q(n973));
  XNOR2X2 U1429(.IN1(n964),.IN2(\add_105_I40_L14036_C136/carry[5] ),.Q(N2235));
  HADDX2 U1430(.A0(\add_90_I16_L14036_C132/carry[3] ),.B0(N518),.C1(\add_90_I16_L14036_C132/carry[4] ),.SO(N529));
  HADDX2 U1431(.A0(\add_105_I39_L14036_C136/carry[2] ),.B0(N2206),.C1(\add_105_I39_L14036_C136/carry[3] ),.SO(N2216));
  NAND3X1 U1432(.IN1(n475),.IN2(n474),.IN3(n476),.QN(n472));
  AO22X1 U1433(.IN1(N2055),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n932),.Q(N2061));
  AO22X1 U1434(.IN1(N2055),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n932),.Q(n920));
  DELLN1X2 U1435(.INP(N1879),.Z(n862));
  HADDX2 U1436(.A0(\add_105_I41_L14036_C136/carry[2] ),.B0(N2238),.C1(\add_105_I41_L14036_C136/carry[3] ),.SO(N2248));
  DELLN1X2 U1437(.INP(N448),.Z(n863));
  DELLN1X2 U1438(.INP(N857),.Z(n864));
  AO22X1 U1439(.IN1(N1879),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n941),.Q(N1885));
  AO22X1 U1440(.IN1(n862),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n941),.Q(n925));
  AO22X1 U1441(.IN1(N1767),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n153),.Q(N1773));
  AO22X1 U1442(.IN1(N1767),.IN2(n222),.IN3(s_fract_48_i[10:10]),.IN4(n153),.Q(n1091));
  AOI22X1 U1443(.IN1(N2171),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1061),.QN(n866));
  HADDX1 U1444(.A0(\add_105_I15_L14036_C136/carry[4] ),.B0(N1824),.C1(\add_105_I15_L14036_C136/carry[5] ),.SO(N1834));
  AO22X1 U1445(.IN1(N1835),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n913),.Q(N1841));
  AO22X1 U1446(.IN1(N1719),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n998),.Q(N1725));
  AO22X1 U1447(.IN1(N1719),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n998),.Q(n953));
  DELLN1X2 U1448(.INP(N2071),.Z(n867));
  HADDX2 U1449(.A0(\add_105_I38_L14036_C136/carry[3] ),.B0(n621),.C1(\add_105_I38_L14036_C136/carry[4] ),.SO(N2201));
  AO22X1 U1450(.IN1(N2071),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N2061),.Q(N2077));
  XNOR2X1 U1451(.IN1(\add_105_I21_L14036_C136/carry[5] ),.IN2(n869),.Q(N1931));
  AOI22X1 U1452(.IN1(N1915),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n999),.QN(n869));
  HADDX2 U1453(.A0(N1708),.B0(N1709),.C1(\add_105_I8_L14036_C136/carry[2] ),.SO(N1719));
  INVX0 U1454(.INP(n106),.ZN(n870));
  HADDX2 U1455(.A0(N2092),.B0(N2093),.C1(\add_105_I32_L14036_C136/carry[2] ),.SO(N2103));
  HADDX2 U1456(.A0(\add_105_I32_L14036_C136/carry[2] ),.B0(N2094),.C1(\add_105_I32_L14036_C136/carry[3] ),.SO(N2104));
  HADDX2 U1457(.A0(N1677),.B0(N1678),.C1(\add_105_I6_L14036_C136/carry[2] ),.SO(N1687));
  HADDX2 U1458(.A0(\add_105_I38_L14036_C136/carry[2] ),.B0(n689),.C1(\add_105_I38_L14036_C136/carry[3] ),.SO(N2200));
  HADDX2 U1459(.A0(N1852),.B0(N1853),.C1(\add_105_I17_L14036_C136/carry[2] ),.SO(N1863));
  HADDX2 U1460(.A0(\add_90_I20_L14036_C132/carry[3] ),.B0(N586),.C1(\add_90_I20_L14036_C132/carry[4] ),.SO(N597));
  AO22X1 U1461(.IN1(n141),.IN2(n164),.IN3(n1217),.IN4(n33),.Q(n872));
  HADDX2 U1462(.A0(N1916),.B0(N1917),.C1(\add_105_I21_L14036_C136/carry[2] ),.SO(N1927));
  AOI22X1 U1463(.IN1(N1947),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(N1937),.QN(n873));
  AO22X1 U1464(.IN1(N715),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n500),.Q(n874));
  HADDX2 U1465(.A0(\add_105_I19_L14036_C136/carry[3] ),.B0(N1887),.C1(\add_105_I19_L14036_C136/carry[4] ),.SO(N1897));
  HADDX2 U1466(.A0(N1804),.B0(N1805),.C1(\add_105_I14_L14036_C136/carry[2] ),.SO(N1815));
  HADDX2 U1467(.A0(\add_90_I7_L14036_C132/carry[2] ),.B0(N364),.C1(\add_90_I7_L14036_C132/carry[3] ),.SO(N375));
  HADDX2 U1468(.A0(N668),.B0(N669),.C1(\add_90_I25_L14036_C132/carry[2] ),.SO(N680));
  AO22X1 U1469(.IN1(N375),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(N364),.Q(N381));
  DELLN1X2 U1470(.INP(N839),.Z(n878));
  AO22X1 U1471(.IN1(N732),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n874),.Q(N738));
  HADDX2 U1472(.A0(\add_90_I28_L14036_C132/carry[2] ),.B0(N721),.C1(\add_90_I28_L14036_C132/carry[3] ),.SO(N732));
  AO22X1 U1473(.IN1(N1895),.IN2(n204),.IN3(n1214),.IN4(n925),.Q(n879));
  AOI22X1 U1474(.IN1(N2075),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n1052),.QN(n880));
  HADDX2 U1475(.A0(\add_90_I35_L14036_C132/carry[2] ),.B0(N840),.C1(\add_90_I35_L14036_C132/carry[3] ),.SO(N851));
  HADDX2 U1476(.A0(N1980),.B0(N1981),.C1(\add_105_I25_L14036_C136/carry[2] ),.SO(N1991));
  AOI22X2 U1477(.IN1(n864),.IN2(n1211),.IN3(n743),.IN4(n619),.QN(n711));
  HADDX2 U1478(.A0(\add_90_I37_L14036_C132/carry[3] ),.B0(N875),.C1(\add_90_I37_L14036_C132/carry[4] ),.SO(N886));
  AOI22X1 U1479(.IN1(N971),.IN2(n227),.IN3(n1220),.IN4(n860),.QN(n882));
  XNOR2X1 U1480(.IN1(\add_105_I30_L14036_C136/carry[5] ),.IN2(n883),.Q(N2075));
  AOI22X1 U1481(.IN1(N2059),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n995),.QN(n883));
  AO22X1 U1482(.IN1(N2251),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1021),.Q(n926));
  AO22X2 U1483(.IN1(N1911),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(N1901),.Q(n885));
  HADDX2 U1484(.A0(N1900),.B0(n879),.C1(\add_105_I20_L14036_C136/carry[2] ),.SO(N1911));
  AO22X2 U1485(.IN1(N1880),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1049),.Q(n887));
  AO22X1 U1486(.IN1(N1755),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n935),.Q(n888));
  XOR2X1 U1487(.IN1(\add_105_I10_L14036_C136/carry[5] ),.IN2(N1745),.Q(N1755));
  AOI22X2 U1488(.IN1(n1007),.IN2(s_fract_48_i[36:36]),.IN3(n591),.IN4(n587),.QN(n665));
  AO22X1 U1489(.IN1(N478),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n591),.Q(N484));
  AO22X1 U1490(.IN1(N1799),.IN2(n215),.IN3(n1210),.IN4(N1789),.Q(n890));
  HADDX2 U1491(.A0(N1884),.B0(N1885),.C1(\add_105_I19_L14036_C136/carry[2] ),.SO(N1895));
  HADDX2 U1492(.A0(N1868),.B0(N1869),.C1(\add_105_I18_L14036_C136/carry[2] ),.SO(N1879));
  XOR2X1 U1493(.IN1(\add_105_I16_L14036_C136/carry[5] ),.IN2(N1841),.Q(N1851));
  HADDX2 U1494(.A0(N2252),.B0(N2253),.C1(\add_105_I42_L14036_C136/carry[2] ),.SO(N2263));
  AO22X2 U1495(.IN1(N2328),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n43),.Q(n892));
  HADDX2 U1496(.A0(N2108),.B0(N2109),.C1(\add_105_I33_L14036_C136/carry[2] ),.SO(N2119));
  HADDX2 U1497(.A0(N2140),.B0(N2141),.C1(\add_105_I35_L14036_C136/carry[2] ),.SO(N2151));
  XNOR2X2 U1498(.IN1(n228),.IN2(\add_105_I43_L14036_C136/carry[5] ),.Q(n1139));
  XNOR2X1 U1499(.IN1(\add_105_I41_L14036_C136/carry[5] ),.IN2(n966),.Q(N2251));
  HADDX2 U1500(.A0(\add_90_I13_L14036_C132/carry[2] ),.B0(N466),.C1(\add_90_I13_L14036_C132/carry[3] ),.SO(N477));
  DELLN1X2 U1501(.INP(N2301),.Z(n896));
  AO22X1 U1502(.IN1(N1867),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n919),.Q(n897));
  AO22X1 U1503(.IN1(N1706),.IN2(n226),.IN3(n1226),.IN4(N1696),.Q(n898));
  AO22X1 U1504(.IN1(N629),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n994),.Q(n899));
  DELLN1X2 U1505(.INP(N823),.Z(n900));
  HADDX2 U1506(.A0(N719),.B0(N720),.C1(\add_90_I28_L14036_C132/carry[2] ),.SO(N731));
  DELLN1X2 U1507(.INP(N788),.Z(n902));
  AO22X1 U1508(.IN1(N2346),.IN2(n69),.IN3(n1205),.IN4(n991),.Q(n903));
  AO22X1 U1509(.IN1(N1979),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n943),.Q(n905));
  AO22X1 U1510(.IN1(N2074),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n807),.Q(N2080));
  INVX0 U1511(.INP(N401),.ZN(n906));
  INVX0 U1512(.INP(n906),.ZN(n907));
  DELLN1X2 U1513(.INP(N551),.Z(n908));
  AO22X1 U1514(.IN1(N428),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N417),.Q(N434));
  HADDX2 U1515(.A0(\add_105_I17_L14036_C136/carry[3] ),.B0(N1855),.C1(\add_105_I17_L14036_C136/carry[4] ),.SO(N1865));
  HADDX2 U1516(.A0(\add_105_I18_L14036_C136/carry[3] ),.B0(N1871),.C1(\add_105_I18_L14036_C136/carry[4] ),.SO(N1881));
  INVX0 U1517(.INP(N364),.ZN(n910));
  INVX0 U1518(.INP(n910),.ZN(n911));
  DELLN1X2 U1519(.INP(N1760),.Z(n912));
  INVX0 U1520(.INP(n241),.ZN(n914));
  HADDX2 U1521(.A0(N2060),.B0(n920),.C1(\add_105_I30_L14036_C136/carry[2] ),.SO(N2071));
  HADDX2 U1522(.A0(N1756),.B0(N1757),.C1(\add_105_I11_L14036_C136/carry[2] ),.SO(N1767));
  DELLN1X2 U1523(.INP(N1758),.Z(n916));
  AO22X1 U1524(.IN1(N1835),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n913),.Q(n1010));
  AOI222X2 U1525(.IN1(n658),.IN2(n389),.IN3(n1060),.IN4(n1213),.IN5(n49),.IN6(n390),.QN(n427));
  AO22X1 U1526(.IN1(N1945),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n658),.Q(N1951));
  AO22X1 U1527(.IN1(N1754),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n176),.Q(N1760));
  HADDX2 U1528(.A0(N2044),.B0(N2045),.C1(\add_105_I29_L14036_C136/carry[2] ),.SO(N2055));
  HADDX2 U1529(.A0(N1836),.B0(N1837),.C1(\add_105_I16_L14036_C136/carry[2] ),.SO(N1847));
  AND2X4 U1530(.IN1(N378),.IN2(n137),.Q(n1196));
  HADDX2 U1531(.A0(N349),.B0(\add_90_I6_L14036_C132/carry[3] ),.C1(N360),.SO(N359));
  AO22X1 U1532(.IN1(N544),.IN2(n164),.IN3(n1217),.IN4(n1081),.Q(n921));
  AO22X1 U1533(.IN1(N530),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1107),.Q(n922));
  DELLN1X2 U1534(.INP(N554),.Z(n923));
  HADDX2 U1535(.A0(N2028),.B0(N2029),.C1(\add_105_I28_L14036_C136/carry[2] ),.SO(N2039));
  AO22X1 U1536(.IN1(N2235),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n1085),.Q(n1021));
  XOR2X1 U1537(.IN1(\add_105_I12_L14036_C136/carry[5] ),.IN2(N1777),.Q(N1787));
  HADDX2 U1538(.A0(N1932),.B0(N1933),.C1(\add_105_I22_L14036_C136/carry[2] ),.SO(N1943));
  HADDX2 U1539(.A0(N2012),.B0(N2013),.C1(\add_105_I27_L14036_C136/carry[2] ),.SO(N2023));
  AO22X1 U1540(.IN1(N1832),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n833),.Q(N1838));
  HADDX2 U1541(.A0(N1996),.B0(N1997),.C1(\add_105_I26_L14036_C136/carry[2] ),.SO(N2007));
  HADDX2 U1542(.A0(\add_105_I33_L14036_C136/carry[2] ),.B0(N2110),.C1(\add_105_I33_L14036_C136/carry[3] ),.SO(N2120));
  AO22X1 U1543(.IN1(N1737),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n939),.Q(n927));
  AOI22X1 U1544(.IN1(N1801),.IN2(n215),.IN3(n1211),.IN4(n1014),.QN(n928));
  HADDX2 U1545(.A0(\add_105_I40_L14036_C136/carry[2] ),.B0(n192),.C1(\add_105_I40_L14036_C136/carry[3] ),.SO(N2232));
  AO22X1 U1546(.IN1(N870),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1035),.Q(n929));
  AO22X1 U1547(.IN1(N578),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n834),.Q(n930));
  DELLN1X2 U1548(.INP(N517),.Z(n931));
  AO22X1 U1549(.IN1(N1994),.IN2(n177),.IN3(n1290),.IN4(n219),.Q(N2000));
  AO22X1 U1550(.IN1(N2039),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n963),.Q(n932));
  AO22X1 U1551(.IN1(N2042),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n217),.Q(N2048));
  AO22X1 U1552(.IN1(N646),.IN2(n177),.IN3(n1289),.IN4(n899),.Q(N652));
  HADDX2 U1553(.A0(N634),.B0(N635),.C1(\add_90_I23_L14036_C132/carry[2] ),.SO(N646));
  INVX0 U1554(.INP(N976),.ZN(n933));
  INVX0 U1555(.INP(n933),.ZN(n934));
  AO22X1 U1556(.IN1(N920),.IN2(n224),.IN3(s_fract_48_i[8:8]),.IN4(n847),.Q(N926));
  AO22X1 U1557(.IN1(N871),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n1044),.Q(n936));
  AO22X1 U1558(.IN1(N429),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n1032),.Q(n937));
  AO22X1 U1559(.IN1(N2312),.IN2(n119),.IN3(s_fract_48_i[44:44]),.IN4(n148),.Q(N2318));
  HADDX2 U1560(.A0(\add_105_I35_L14036_C136/carry[2] ),.B0(N2142),.C1(\add_105_I35_L14036_C136/carry[3] ),.SO(N2152));
  DELLN1X2 U1561(.INP(N468),.Z(n938));
  DELLN1X2 U1562(.INP(N1729),.Z(n940));
  AOI222X2 U1563(.IN1(n243),.IN2(n389),.IN3(N1901),.IN4(n1213),.IN5(n885),.IN6(n390),.QN(n494));
  AO22X1 U1564(.IN1(N1911),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(N1901),.Q(N1917));
  AO22X1 U1565(.IN1(N1863),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n954),.Q(n941));
  DELLN1X2 U1566(.INP(N894),.Z(n942));
  AO22X1 U1567(.IN1(N649),.IN2(n177),.IN3(n1289),.IN4(n1097),.Q(N655));
  AO22X1 U1568(.IN1(N1963),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N1953),.Q(n943));
  AOI222X1 U1569(.IN1(n577),.IN2(n907),.IN3(n578),.IN4(n937),.IN5(n1387),.IN6(n579),.QN(n971));
  DELLN1X2 U1570(.INP(N485),.Z(n944));
  HADDX1 U1571(.A0(N1712),.B0(\add_105_I8_L14036_C136/carry[4] ),.C1(\add_105_I8_L14036_C136/carry[5] ),.SO(N1722));
  DELLN1X2 U1572(.INP(N724),.Z(n946));
  AO22X1 U1573(.IN1(N1975),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1041),.Q(n947));
  HADDX2 U1574(.A0(N1964),.B0(N1965),.C1(\add_105_I24_L14036_C136/carry[2] ),.SO(N1975));
  HADDX2 U1575(.A0(\add_105_I12_L14036_C136/carry[2] ),.B0(N1774),.C1(\add_105_I12_L14036_C136/carry[3] ),.SO(N1784));
  XNOR2X1 U1576(.IN1(\add_105_I36_L14036_C136/carry[5] ),.IN2(n948),.Q(N2171));
  AOI22X1 U1577(.IN1(N2155),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n1016),.QN(n948));
  XNOR2X1 U1578(.IN1(n118),.IN2(s_fract_48_i[46:46]),.Q(n949));
  AO22X1 U1579(.IN1(N2314),.IN2(n47),.IN3(s_fract_48_i[44:44]),.IN4(n63),.Q(n950));
  AO22X1 U1580(.IN1(N2314),.IN2(n47),.IN3(s_fract_48_i[44:44]),.IN4(n63),.Q(N2320));
  AO22X1 U1581(.IN1(N2121),.IN2(n160),.IN3(s_fract_48_i[32:32]),.IN4(n817),.Q(N2127));
  AO22X1 U1582(.IN1(N1880),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n1049),.Q(N1886));
  AO22X1 U1583(.IN1(N1864),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n149),.Q(N1870));
  DELLN1X2 U1584(.INP(N1720),.Z(n952));
  HADDX2 U1585(.A0(\add_105_I8_L14036_C136/carry[2] ),.B0(N1710),.C1(\add_105_I8_L14036_C136/carry[3] ),.SO(N1720));
  AO22X1 U1586(.IN1(N1847),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n157),.Q(n954));
  AO22X1 U1587(.IN1(N1914),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n996),.Q(N1920));
  HADDX2 U1588(.A0(\add_105_I20_L14036_C136/carry[4] ),.B0(N1904),.C1(\add_105_I20_L14036_C136/carry[5] ),.SO(N1914));
  AO22X1 U1589(.IN1(n221),.IN2(N1785),.IN3(s_fract_48_i[11:11]),.IN4(n203),.Q(N1791));
  AO22X1 U1590(.IN1(N1720),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1001),.Q(N1726));
  HADDX2 U1591(.A0(\add_90_I26_L14036_C132/carry[3] ),.B0(N688),.C1(\add_90_I26_L14036_C132/carry[4] ),.SO(N699));
  XNOR2X1 U1592(.IN1(\add_90_I24_L14036_C132/carry[5] ),.IN2(n957),.Q(N667));
  AOI22X1 U1593(.IN1(N650),.IN2(n177),.IN3(n1289),.IN4(n986),.QN(n957));
  DELLN1X2 U1594(.INP(N738),.Z(n958));
  HADDX2 U1595(.A0(N334),.B0(\add_90_I5_L14036_C132/carry[2] ),.C1(N344),.SO(N343));
  AO22X1 U1596(.IN1(N2152),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n877),.Q(n960));
  AO22X1 U1597(.IN1(N2202),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(n32),.Q(N2208));
  HADDX2 U1598(.A0(\add_105_I36_L14036_C136/carry[3] ),.B0(n712),.C1(\add_105_I36_L14036_C136/carry[4] ),.SO(N2169));
  DELLN1X2 U1599(.INP(N2250),.Z(n961));
  HADDX2 U1600(.A0(\add_105_I44_L14036_C136/carry[4] ),.B0(N2288),.C1(\add_105_I44_L14036_C136/carry[5] ),.SO(N2298));
  AO22X1 U1601(.IN1(N2023),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n985),.Q(n963));
  AO22X1 U1602(.IN1(N2250),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1047),.Q(n1017));
  AO22X1 U1603(.IN1(N2266),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(N2256),.Q(N2272));
  AO22X1 U1604(.IN1(n122),.IN2(N2298),.IN3(s_fract_48_i[43:43]),.IN4(n990),.Q(N2304));
  AOI22X1 U1605(.IN1(N2219),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n1019),.QN(n964));
  AO22X1 U1606(.IN1(N2087),.IN2(n164),.IN3(n1216),.IN4(n915),.Q(n965));
  HADDX2 U1607(.A0(N2076),.B0(N2077),.C1(\add_105_I31_L14036_C136/carry[2] ),.SO(N2087));
  AOI22X1 U1608(.IN1(N2235),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n1085),.QN(n966));
  HADDX2 U1609(.A0(\add_105_I29_L14036_C136/carry[3] ),.B0(N2047),.C1(\add_105_I29_L14036_C136/carry[4] ),.SO(N2057));
  OAI221X1 U1610(.IN1(n967),.IN2(n968),.IN3(n969),.IN4(n970),.IN5(n971),.QN(n1128));
  HADDX2 U1611(.A0(N2124),.B0(N2125),.C1(\add_105_I34_L14036_C136/carry[2] ),.SO(N2135));
  AO22X1 U1612(.IN1(N956),.IN2(n226),.IN3(n1224),.IN4(n1027),.Q(n974));
  AO22X1 U1613(.IN1(N939),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1009),.Q(n1027));
  AO22X1 U1614(.IN1(N1931),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n1029),.Q(n975));
  AO22X1 U1615(.IN1(N2072),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(N2062),.Q(N2078));
  XOR2X1 U1616(.IN1(\add_90_I34_L14036_C132/carry[5] ),.IN2(N826),.Q(N837));
  AO22X1 U1617(.IN1(N664),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n576),.Q(n976));
  HADDX2 U1618(.A0(\add_90_I24_L14036_C132/carry[2] ),.B0(N653),.C1(\add_90_I24_L14036_C132/carry[3] ),.SO(N664));
  HADDX2 U1619(.A0(\add_90_I40_L14036_C132/carry[3] ),.B0(N926),.C1(\add_90_I40_L14036_C132/carry[4] ),.SO(N937));
  AOI22X1 U1620(.IN1(N904),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n1095),.QN(n1058));
  AO22X1 U1621(.IN1(N2057),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n185),.Q(N2063));
  AO22X1 U1622(.IN1(N2057),.IN2(n171),.IN3(s_fract_48_i[28:28]),.IN4(n185),.Q(n1086));
  HADDX2 U1623(.A0(\add_105_I31_L14036_C136/carry[2] ),.B0(N2078),.C1(\add_105_I31_L14036_C136/carry[3] ),.SO(N2088));
  HADDX2 U1624(.A0(\add_105_I37_L14036_C136/carry[3] ),.B0(N2175),.C1(\add_105_I37_L14036_C136/carry[4] ),.SO(N2185));
  DELLN1X2 U1625(.INP(N2125),.Z(n978));
  XOR2X1 U1626(.IN1(\add_105_I19_L14036_C136/carry[5] ),.IN2(N1889),.Q(N1899));
  AO22X1 U1627(.IN1(N632),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1098),.Q(N638));
  AO22X1 U1628(.IN1(n140),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1141),.Q(n1131));
  AO22X1 U1629(.IN1(N2170),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1141),.Q(N2176));
  OAI22X1 U1630(.IN1(n1231),.IN2(n1139),.IN3(n123),.IN4(n51),.QN(N2289));
  AO22X1 U1631(.IN1(N667),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1036),.Q(n979));
  DELLN1X2 U1632(.INP(N772),.Z(n980));
  AO22X1 U1633(.IN1(N493),.IN2(n158),.IN3(s_fract_48_i[33:33]),.IN4(n839),.Q(n981));
  HADDX2 U1634(.A0(\add_90_I24_L14036_C132/carry[3] ),.B0(N654),.C1(\add_90_I24_L14036_C132/carry[4] ),.SO(N665));
  AO22X1 U1635(.IN1(N648),.IN2(n177),.IN3(n1290),.IN4(n1108),.Q(N654));
  DELLN1X2 U1636(.INP(N2013),.Z(n985));
  DELLN1X2 U1637(.INP(N689),.Z(n987));
  AO22X1 U1638(.IN1(n961),.IN2(n137),.IN3(s_fract_48_i[40:40]),.IN4(n1047),.Q(N2256));
  AO22X1 U1639(.IN1(N701),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n1000),.Q(N707));
  DELLN1X2 U1640(.INP(n803),.Z(n988));
  DELLN1X2 U1641(.INP(N756),.Z(n989));
  AO22X1 U1642(.IN1(n136),.IN2(n123),.IN3(n1229),.IN4(n1042),.Q(n990));
  AO22X1 U1643(.IN1(N752),.IN2(n204),.IN3(n1214),.IN4(n824),.Q(N758));
  AOI22X2 U1644(.IN1(n827),.IN2(s_fract_48_i[36:36]),.IN3(n938),.IN4(n587),.QN(n639));
  HADDX2 U1645(.A0(\add_90_I14_L14036_C132/carry[3] ),.B0(N484),.C1(\add_90_I14_L14036_C132/carry[4] ),.SO(N495));
  HADDX2 U1646(.A0(\add_90_I11_L14036_C132/carry[3] ),.B0(N433),.C1(\add_90_I11_L14036_C132/carry[4] ),.SO(N444));
  AO22X1 U1647(.IN1(N700),.IN2(n196),.IN3(s_fract_48_i[21:21]),.IN4(n987),.Q(n992));
  HADDX2 U1648(.A0(\add_90_I26_L14036_C132/carry[4] ),.B0(N689),.C1(\add_90_I26_L14036_C132/carry[5] ),.SO(N700));
  AO22X1 U1649(.IN1(N1687),.IN2(n227),.IN3(n1223),.IN4(n1024),.Q(n993));
  AO22X2 U1650(.IN1(N1673),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n1134),.Q(n1024));
  AO22X1 U1651(.IN1(N1753),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n927),.Q(N1759));
  HADDX2 U1652(.A0(N600),.B0(N601),.C1(\add_90_I21_L14036_C132/carry[2] ),.SO(N612));
  AO22X1 U1653(.IN1(N784),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n634),.Q(N790));
  HADDX2 U1654(.A0(\add_105_I7_L14036_C136/carry[2] ),.B0(N1694),.C1(\add_105_I7_L14036_C136/carry[3] ),.SO(N1704));
  DELLN1X2 U1655(.INP(N1904),.Z(n996));
  XOR2X2 U1656(.IN1(\add_105_I8_L14036_C136/carry[5] ),.IN2(n1195),.Q(N1723));
  HADDX2 U1657(.A0(\add_105_I31_L14036_C136/carry[3] ),.B0(N2079),.C1(\add_105_I31_L14036_C136/carry[4] ),.SO(N2089));
  DELLN1X2 U1658(.INP(N754),.Z(n997));
  AO22X1 U1659(.IN1(N1703),.IN2(n226),.IN3(n1225),.IN4(n993),.Q(n998));
  AO22X1 U1660(.IN1(n13),.IN2(n204),.IN3(n1213),.IN4(n1025),.Q(n999));
  HADDX2 U1661(.A0(\add_105_I41_L14036_C136/carry[4] ),.B0(N2240),.C1(\add_105_I41_L14036_C136/carry[5] ),.SO(N2250));
  AO22X1 U1662(.IN1(N2234),.IN2(n144),.IN3(s_fract_48_i[39:39]),.IN4(n1078),.Q(N2240));
  AO22X1 U1663(.IN1(N2091),.IN2(n164),.IN3(n1216),.IN4(N2081),.Q(N2097));
  AO22X1 U1664(.IN1(n858),.IN2(n226),.IN3(n1227),.IN4(n163),.Q(n1001));
  AO22X2 U1665(.IN1(N837),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n1012),.Q(n1002));
  AO22X1 U1666(.IN1(n471),.IN2(n212),.IN3(s_fract_48_i[14:14]),.IN4(n1005),.Q(n1012));
  DELLN1X2 U1667(.INP(N703),.Z(n1003));
  AOI222X1 U1668(.IN1(n332),.IN2(n940),.IN3(n333),.IN4(n1195),.IN5(n334),.IN6(n935),.QN(n1112));
  AO22X1 U1669(.IN1(N1755),.IN2(n223),.IN3(s_fract_48_i[9:9]),.IN4(n935),.Q(N1761));
  DELLN1X2 U1670(.INP(N687),.Z(n1004));
  HADDX2 U1671(.A0(\add_90_I11_L14036_C132/carry[2] ),.B0(n242),.C1(\add_90_I11_L14036_C132/carry[3] ),.SO(N443));
  DELLN1X2 U1672(.INP(N434),.Z(n1006));
  HADDX2 U1673(.A0(\add_105_I14_L14036_C136/carry[2] ),.B0(N1806),.C1(\add_105_I14_L14036_C136/carry[3] ),.SO(N1816));
  HADDX2 U1674(.A0(\add_105_I34_L14036_C136/carry[2] ),.B0(n812),.C1(\add_105_I34_L14036_C136/carry[3] ),.SO(N2136));
  INVX0 U1675(.INP(n882),.ZN(n1008));
  HADDX2 U1676(.A0(\add_90_I34_L14036_C132/carry[2] ),.B0(n336),.C1(\add_90_I34_L14036_C132/carry[3] ),.SO(N834));
  HADDX2 U1677(.A0(N736),.B0(N737),.C1(\add_90_I29_L14036_C132/carry[2] ),.SO(N748));
  AO22X1 U1678(.IN1(n9),.IN2(n227),.IN3(N1680),.IN4(n1221),.Q(n1013));
  HADDX2 U1679(.A0(N1680),.B0(\add_105_I6_L14036_C136/carry[3] ),.C1(N1690),.SO(N1689));
  DELLN1X2 U1680(.INP(N1791),.Z(n1014));
  AO22X1 U1681(.IN1(N599),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1037),.Q(n1015));
  AO22X1 U1682(.IN1(N599),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1037),.Q(N605));
  HADDX2 U1683(.A0(\add_105_I42_L14036_C136/carry[4] ),.B0(n1017),.C1(\add_105_I42_L14036_C136/carry[5] ),.SO(N2266));
  DELLN1X2 U1684(.INP(N652),.Z(n1020));
  DELLN1X2 U1685(.INP(N2000),.Z(n1023));
  AO22X2 U1686(.IN1(N1883),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(N1873),.Q(n1025));
  HADDX2 U1687(.A0(\add_105_I40_L14036_C136/carry[4] ),.B0(N2224),.C1(\add_105_I40_L14036_C136/carry[5] ),.SO(N2234));
  AO22X1 U1688(.IN1(N2218),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n700),.Q(N2224));
  AO22X1 U1689(.IN1(N1912),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1050),.Q(N1918));
  AO22X1 U1690(.IN1(N1897),.IN2(n204),.IN3(n1214),.IN4(n1026),.Q(N1903));
  AO22X1 U1691(.IN1(N596),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n1031),.Q(n1028));
  HADDX2 U1692(.A0(\add_90_I20_L14036_C132/carry[2] ),.B0(N585),.C1(\add_90_I20_L14036_C132/carry[3] ),.SO(N596));
  AO22X2 U1693(.IN1(N1915),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n999),.Q(n1029));
  HADDX2 U1694(.A0(\add_105_I17_L14036_C136/carry[2] ),.B0(N1854),.C1(\add_105_I17_L14036_C136/carry[3] ),.SO(N1864));
  AO22X1 U1695(.IN1(N1913),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1060),.Q(N1919));
  AO22X1 U1696(.IN1(N1995),.IN2(n177),.IN3(n1289),.IN4(N1985),.Q(n1030));
  DELLN1X2 U1697(.INP(N585),.Z(n1031));
  AO22X1 U1698(.IN1(N2073),.IN2(n170),.IN3(s_fract_48_i[29:29]),.IN4(n1086),.Q(N2079));
  HADDX2 U1699(.A0(\add_105_I30_L14036_C136/carry[3] ),.B0(N2063),.C1(\add_105_I30_L14036_C136/carry[4] ),.SO(N2073));
  AO22X1 U1700(.IN1(N1799),.IN2(n215),.IN3(n1210),.IN4(N1789),.Q(N1805));
  HADDX2 U1701(.A0(N1788),.B0(n155),.C1(\add_105_I13_L14036_C136/carry[2] ),.SO(N1799));
  AO22X1 U1702(.IN1(N1800),.IN2(n215),.IN3(n1211),.IN4(n240),.Q(N1806));
  HADDX2 U1703(.A0(\add_105_I13_L14036_C136/carry[2] ),.B0(N1790),.C1(\add_105_I13_L14036_C136/carry[3] ),.SO(N1800));
  AOI222X2 U1704(.IN1(n1336),.IN2(N2363),.IN3(n385),.IN4(n31),.IN5(n386),.IN6(n845),.QN(n1187));
  INVX0 U1705(.INP(n959),.ZN(n1033));
  AO22X1 U1706(.IN1(N2089),.IN2(n164),.IN3(n1217),.IN4(n62),.Q(N2095));
  AOI22X2 U1707(.IN1(N2266),.IN2(n130),.IN3(s_fract_48_i[41:41]),.IN4(N2256),.QN(n1034));
  AO22X1 U1708(.IN1(N853),.IN2(n215),.IN3(n1210),.IN4(n1088),.Q(n1035));
  AO22X2 U1709(.IN1(n161),.IN2(n177),.IN3(n1289),.IN4(n986),.Q(n1036));
  AO22X1 U1710(.IN1(N2041),.IN2(n172),.IN3(s_fract_48_i[27:27]),.IN4(n213),.Q(N2047));
  DELLN1X2 U1711(.INP(N588),.Z(n1037));
  AOI22X1 U1712(.IN1(N615),.IN2(n173),.IN3(s_fract_48_i[26:26]),.IN4(n983),.QN(n1039));
  DELLN1X2 U1713(.INP(N1792),.Z(n1040));
  AO22X1 U1714(.IN1(N1786),.IN2(n221),.IN3(s_fract_48_i[11:11]),.IN4(n951),.Q(N1792));
  AO22X1 U1715(.IN1(N1959),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(N1949),.Q(n1041));
  HADDX2 U1716(.A0(N1948),.B0(n168),.C1(\add_105_I23_L14036_C136/carry[2] ),.SO(N1959));
  INVX0 U1717(.INP(n1034),.ZN(n1042));
  DELLN1X2 U1718(.INP(N860),.Z(n1044));
  XOR2X1 U1719(.IN1(\add_105_I44_L14036_C136/carry[5] ),.IN2(N2289),.Q(N2299));
  AO22X1 U1720(.IN1(N1865),.IN2(n208),.IN3(s_fract_48_i[16:16]),.IN4(n28),.Q(N1871));
  AOI22X1 U1721(.IN1(N631),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n984),.QN(n1045));
  HADDX2 U1722(.A0(N1692),.B0(N1693),.C1(\add_105_I7_L14036_C136/carry[2] ),.SO(N1703));
  AOI22X1 U1723(.IN1(n852),.IN2(n334),.IN3(n993),.IN4(n1223),.QN(n482));
  AO22X1 U1724(.IN1(n138),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n700),.Q(n1078));
  AO22X1 U1725(.IN1(N1023),.IN2(n1136),.IN3(s_fract_48_i[2:2]),.IN4(n1126),.Q(n1048));
  DELLN1X2 U1726(.INP(N1870),.Z(n1049));
  DELLN1X2 U1727(.INP(N1902),.Z(n1050));
  AO22X1 U1728(.IN1(N1850),.IN2(n210),.IN3(s_fract_48_i[15:15]),.IN4(n207),.Q(N1856));
  HADDX2 U1729(.A0(\add_90_I31_L14036_C132/carry[4] ),.B0(N774),.C1(\add_90_I31_L14036_C132/carry[5] ),.SO(N785));
  DELLN1X2 U1730(.INP(N792),.Z(n1051));
  DELLN1X2 U1731(.INP(N2127),.Z(n1054));
  INVX0 U1732(.INP(n159),.ZN(n1055));
  NBUFFX4 U1733(.INP(s_fract_48_i[12:12]),.Z(n1209));
  DELLN1X2 U1734(.INP(N673),.Z(n1057));
  DELLN1X2 U1735(.INP(N1966),.Z(n1059));
  DELLN1X2 U1736(.INP(N1903),.Z(n1060));
  HADDX2 U1737(.A0(\add_105_I39_L14036_C136/carry[4] ),.B0(N2208),.C1(\add_105_I39_L14036_C136/carry[5] ),.SO(N2218));
  AOI22X1 U1738(.IN1(N632),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1098),.QN(n1062));
  DELLN1X2 U1739(.INP(N757),.Z(n1063));
  DELLN1X2 U1740(.INP(N671),.Z(n1064));
  AO22X1 U1741(.IN1(N1976),.IN2(n182),.IN3(s_fract_48_i[23:23]),.IN4(n1059),.Q(N1982));
  HADDX2 U1742(.A0(\add_105_I23_L14036_C136/carry[2] ),.B0(N1950),.C1(\add_105_I23_L14036_C136/carry[3] ),.SO(N1960));
  AO22X1 U1743(.IN1(N1993),.IN2(n177),.IN3(n1290),.IN4(n805),.Q(N1999));
  XOR2X2 U1744(.IN1(\add_90_I10_L14036_C132/carry[5] ),.IN2(N418),.Q(N429));
  HADDX2 U1745(.A0(\add_90_I10_L14036_C132/carry[2] ),.B0(N415),.C1(\add_90_I10_L14036_C132/carry[3] ),.SO(N426));
  DELLN1X2 U1746(.INP(N722),.Z(n1067));
  AOI22X2 U1747(.IN1(n16),.IN2(n345),.IN3(n672),.IN4(n346),.QN(n398));
  AO22X1 U1748(.IN1(N1882),.IN2(n206),.IN3(s_fract_48_i[17:17]),.IN4(n672),.Q(N1888));
  DELLN1X2 U1749(.INP(N601),.Z(n1068));
  DELLN1X2 U1750(.INP(N484),.Z(n1069));
  HADDX2 U1751(.A0(N1740),.B0(N1741),.C1(\add_105_I10_L14036_C136/carry[2] ),.SO(N1751));
  AO22X2 U1752(.IN1(N733),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1067),.Q(n1070));
  HADDX2 U1753(.A0(\add_90_I28_L14036_C132/carry[3] ),.B0(N722),.C1(\add_90_I28_L14036_C132/carry[4] ),.SO(N733));
  DELLN1X2 U1754(.INP(N1999),.Z(n1071));
  AOI222X2 U1755(.IN1(N2222),.IN2(n387),.IN3(N2190),.IN4(s_fract_48_i[36:36]),.IN5(n823),.IN6(n388),.QN(n476));
  DELLN1X2 U1756(.INP(N723),.Z(n1072));
  AO22X1 U1757(.IN1(N734),.IN2(n198),.IN3(s_fract_48_i[19:19]),.IN4(n1072),.Q(N740));
  HADDX2 U1758(.A0(\add_90_I28_L14036_C132/carry[4] ),.B0(N723),.C1(\add_90_I28_L14036_C132/carry[5] ),.SO(N734));
  AO22X2 U1759(.IN1(n603),.IN2(n671),.IN3(n1290),.IN4(n59),.Q(n648));
  AO22X1 U1760(.IN1(N683),.IN2(n189),.IN3(s_fract_48_i[22:22]),.IN4(n671),.Q(N689));
  AO22X1 U1761(.IN1(N2171),.IN2(n154),.IN3(s_fract_48_i[35:35]),.IN4(n1061),.Q(n1073));
  AO22X1 U1762(.IN1(N2328),.IN2(n1130),.IN3(s_fract_48_i[45:45]),.IN4(n43),.Q(N2334));
  DELLN1X2 U1763(.INP(N516),.Z(n1074));
  DELLN1X2 U1764(.INP(N654),.Z(n1075));
  DELLN1X2 U1765(.INP(N758),.Z(n1076));
  INVX0 U1766(.INP(n181),.ZN(n1077));
  DELLN1X2 U1767(.INP(N979),.Z(n1079));
  DELLN1X2 U1768(.INP(N2097),.Z(n1080));
  DELLN1X2 U1769(.INP(N1998),.Z(n1082));
  AOI222X2 U1770(.IN1(n972),.IN2(n359),.IN3(n1082),.IN4(n1289),.IN5(n642),.IN6(n358),.QN(n466));
  AO22X1 U1771(.IN1(N2008),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1082),.Q(N2014));
  DELLN1X2 U1772(.INP(N790),.Z(n1083));
  DELLN1X2 U1773(.INP(N605),.Z(n1084));
  AO22X1 U1774(.IN1(N2219),.IN2(n145),.IN3(s_fract_48_i[38:38]),.IN4(n1019),.Q(n1085));
  AO22X1 U1775(.IN1(N529),.IN2(n162),.IN3(s_fract_48_i[31:31]),.IN4(n1106),.Q(n1087));
  AO22X1 U1776(.IN1(N836),.IN2(n214),.IN3(s_fract_48_i[13:13]),.IN4(n478),.Q(n1088));
  AO22X1 U1777(.IN1(n15),.IN2(n174),.IN3(s_fract_48_i[25:25]),.IN4(n1030),.Q(n1089));
  DELLN1X2 U1778(.INP(N959),.Z(n1090));
  AOI222X2 U1779(.IN1(n200),.IN2(n387),.IN3(N2191),.IN4(s_fract_48_i[36:36]),.IN5(n868),.IN6(n388),.QN(n440));
  AO22X1 U1780(.IN1(N2201),.IN2(n146),.IN3(s_fract_48_i[37:37]),.IN4(N2191),.Q(N2207));
  INVX0 U1781(.INP(n1046),.ZN(n1092));
  DELLN1X2 U1782(.INP(N942),.Z(n1093));
  INVX0 U1783(.INP(n881),.ZN(n1094));
  DELLN1X2 U1784(.INP(N893),.Z(n1095));
  AO22X1 U1785(.IN1(N937),.IN2(n225),.IN3(s_fract_48_i[7:7]),.IN4(n1103),.Q(n1096));
  INVX0 U1786(.INP(n1062),.ZN(n1097));
  AOI222X2 U1787(.IN1(n624),.IN2(N1041),.IN3(n625),.IN4(n901),.IN5(n626),.IN6(n849),.QN(n1182));
  INVX0 U1788(.INP(n1039),.ZN(n1098));
  HADDX2 U1789(.A0(N396),.B0(N397),.C1(\add_90_I9_L14036_C132/carry[2] ),.SO(N408));
  DELLN1X2 U1790(.INP(N993),.Z(n1101));
  AO22X2 U1791(.IN1(N987),.IN2(n229),.IN3(s_fract_48_i[4:4]),.IN4(n934),.Q(N993));
  DELLN1X2 U1792(.INP(N1759),.Z(n1102));
  DELLN1X2 U1793(.INP(N926),.Z(n1103));
  XOR2X2 U1794(.IN1(\add_90_I8_L14036_C132/carry[5] ),.IN2(n1196),.Q(N395));
  DELLN1X2 U1795(.INP(N363),.Z(n1104));
  INVX0 U1796(.INP(n1099),.ZN(n1105));
  DELLN1X2 U1797(.INP(N518),.Z(n1106));
  DELLN1X2 U1798(.INP(N519),.Z(n1107));
  INVX0 U1799(.INP(n1045),.ZN(n1108));
  AO22X1 U1800(.IN1(N1005),.IN2(n231),.IN3(s_fract_48_i[3:3]),.IN4(n193),.Q(N1011));
  INVX0 U1801(.INP(n1053),.ZN(n1109));
  INVX0 U1802(.INP(n871),.ZN(n1110));
  HADDX2 U1803(.A0(\add_105_I38_L14036_C136/carry[4] ),.B0(N2192),.C1(\add_105_I38_L14036_C136/carry[5] ),.SO(N2202));
  AOI21X1 U1804(.IN1(n1112),.IN2(n1111),.IN3(n1513),.QN(N2979));
  OA221X1 U1805(.IN1(n450),.IN2(n57),.IN3(n449),.IN4(n1122),.IN5(n1123),.Q(n1111));
  OAI21X1 U1806(.IN1(n1113),.IN2(n1114),.IN3(n442),.QN(n364));
  AO222X1 U1807(.IN1(n1085),.IN2(n387),.IN3(n977),.IN4(s_fract_48_i[36:36]),.IN5(n1019),.IN6(n388),.Q(n1113));
  OAI221X1 U1808(.IN1(n376),.IN2(n375),.IN3(n51),.IN4(n377),.IN5(n378),.QN(n1114));
  DELLN1X2 U1809(.INP(N961),.Z(n1115));
  XNOR2X2 U1810(.IN1(n568),.IN2(n232),.Q(n571));
  XOR2X1 U1811(.IN1(\add_105_I47_L14036_C136/carry[5] ),.IN2(N2337),.Q(N2347));
  AOI221X1 U1812(.IN1(n1116),.IN2(n1117),.IN3(N1985),.IN4(n1466),.IN5(n1118),.QN(n349));
  NAND2X0 U1813(.IN1(n1185),.IN2(n1184),.QN(n1117));
  OAI22X2 U1814(.IN1(n1323),.IN2(n354),.IN3(n1322),.IN4(n355),.QN(n1118));
  NAND2X0 U1815(.IN1(n531),.IN2(n351),.QN(n352));
  DELLN1X2 U1816(.INP(N502),.Z(n1119));
  DELLN1X2 U1817(.INP(N398),.Z(n1120));
  DELLN1X2 U1818(.INP(N740),.Z(n1121));
  AND4X1 U1819(.IN1(n340),.IN2(n339),.IN3(n341),.IN4(n342),.Q(n1122));
  NAND2X0 U1820(.IN1(n562),.IN2(n449),.QN(n450));
  HADDX2 U1821(.A0(N1696),.B0(\add_105_I7_L14036_C136/carry[4] ),.C1(N1707),.SO(N1706));
  HADDX2 U1822(.A0(N1666),.B0(\add_105_I5_L14036_C136/carry[2] ),.C1(N1675),.SO(N1674));
  INVX0 U1823(.INP(n1058),.ZN(n1124));
  HADDX2 U1824(.A0(\add_90_I21_L14036_C132/carry[4] ),.B0(N604),.C1(\add_90_I21_L14036_C132/carry[5] ),.SO(N615));
  AO22X1 U1825(.IN1(N1930),.IN2(n197),.IN3(s_fract_48_i[20:20]),.IN4(n26),.Q(N1936));
  DELLN1X2 U1826(.INP(N1012),.Z(n1126));
  HADDX2 U1827(.A0(\add_90_I27_L14036_C132/carry[3] ),.B0(N705),.C1(\add_90_I27_L14036_C132/carry[4] ),.SO(N716));
  AND2X1 U1828(.IN1(n1128),.IN2(n1127),.Q(N1637));
  HADDX2 U1829(.A0(\add_90_I21_L14036_C132/carry[3] ),.B0(N603),.C1(\add_90_I21_L14036_C132/carry[4] ),.SO(N614));
  INVX0 U1830(.INP(n118),.ZN(n1129));
  INVX0 U1831(.INP(n1129),.ZN(n1130));
  NOR2X0 U1832(.IN1(n988),.IN2(s_fract_48_i[43:43]),.QN(n1133));
  HADDX2 U1833(.A0(N1664),.B0(N1665),.C1(\add_105_I5_L14036_C136/carry[2] ),.SO(N1673));
  XNOR2X2 U1834(.IN1(n1138),.IN2(n231),.Q(N1664));
  DELLN1X2 U1835(.INP(N1665),.Z(n1134));
  INVX0 U1836(.INP(n1206),.ZN(n1135));
  INVX0 U1837(.INP(s_fract_48_i[2:2]),.ZN(n1136));
  XNOR2X1 U1838(.IN1(n233),.IN2(s_fract_48_i[1:1]),.Q(n1137));
  XNOR2X1 U1839(.IN1(n232),.IN2(n1137),.Q(n1138));
  NBUFFX4 U1840(.INP(s_fract_48_i[42:42]),.Z(n1231));
  NBUFFX4 U1841(.INP(s_fract_48_i[42:42]),.Z(n1228));
  DELLN1X2 U1842(.INP(N1871),.Z(n1140));
  AO22X1 U1843(.IN1(n139),.IN2(n156),.IN3(s_fract_48_i[34:34]),.IN4(n1125),.Q(n1141));
  INVX0 U1844(.INP(n928),.ZN(n1142));
  DELLN1X2 U1845(.INP(N1806),.Z(n1143));
  HADDX2 U1846(.A0(\add_105_I20_L14036_C136/carry[2] ),.B0(N1902),.C1(\add_105_I20_L14036_C136/carry[3] ),.SO(N1912));
  HADDX2 U1847(.A0(\add_105_I17_L14036_C136/carry[4] ),.B0(N1856),.C1(\add_105_I17_L14036_C136/carry[5] ),.SO(N1866));
  HADDX2 U1848(.A0(\add_105_I19_L14036_C136/carry[2] ),.B0(N1886),.C1(\add_105_I19_L14036_C136/carry[3] ),.SO(N1896));
  HADDX2 U1849(.A0(\add_105_I28_L14036_C136/carry[4] ),.B0(N2032),.C1(\add_105_I28_L14036_C136/carry[5] ),.SO(N2042));
  HADDX2 U1850(.A0(\add_105_I21_L14036_C136/carry[3] ),.B0(N1919),.C1(\add_105_I21_L14036_C136/carry[4] ),.SO(N1929));
  HADDX2 U1851(.A0(\add_105_I21_L14036_C136/carry[2] ),.B0(N1918),.C1(\add_105_I21_L14036_C136/carry[3] ),.SO(N1928));
  HADDX2 U1852(.A0(\add_105_I11_L14036_C136/carry[2] ),.B0(n34),.C1(\add_105_I11_L14036_C136/carry[3] ),.SO(N1768));
  HADDX2 U1853(.A0(\add_105_I18_L14036_C136/carry[2] ),.B0(N1870),.C1(\add_105_I18_L14036_C136/carry[3] ),.SO(N1880));
  HADDX2 U1854(.A0(\add_105_I26_L14036_C136/carry[4] ),.B0(N2000),.C1(\add_105_I26_L14036_C136/carry[5] ),.SO(N2010));
  HADDX2 U1855(.A0(\add_105_I24_L14036_C136/carry[4] ),.B0(N1968),.C1(\add_105_I24_L14036_C136/carry[5] ),.SO(N1978));
  NAND2X0 U1856(.IN1(n559),.IN2(n376),.QN(n377));
  AOI221X2 U1857(.IN1(n1465),.IN2(n824),.IN3(n1464),.IN4(n601),.IN5(n602),.QN(n1180));
  NAND2X0 U1858(.IN1(n787),.IN2(n616),.QN(n617));
  NAND2X0 U1859(.IN1(n551),.IN2(n560),.QN(n379));
  NAND2X0 U1860(.IN1(n788),.IN2(n786),.QN(n628));
  NBUFFX2 U1861(.INP(s_shr2[5:5]),.Z(n1285));
  NAND3X0 U1862(.IN1(n1144),.IN2(n1145),.IN3(n1146),.QN(n312));
  NAND3X0 U1863(.IN1(n1147),.IN2(n1148),.IN3(n1149),.QN(n310));
  NAND2X1 U1864(.IN1(n1150),.IN2(n1151),.QN(n311));
  NBUFFX2 U1865(.INP(s_shl2[5:5]),.Z(n1277));
  NAND3X0 U1866(.IN1(n1152),.IN2(n1153),.IN3(n1154),.QN(n285));
  NAND3X0 U1867(.IN1(n1155),.IN2(n1156),.IN3(n1157),.QN(n275));
  NAND3X0 U1868(.IN1(n1158),.IN2(n1159),.IN3(n1160),.QN(n277));
  NAND3X0 U1869(.IN1(n1161),.IN2(n1162),.IN3(n1163),.QN(n267));
  NAND3X0 U1870(.IN1(n1164),.IN2(n1165),.IN3(n1166),.QN(n284));
  NAND3X0 U1871(.IN1(n1167),.IN2(n1168),.IN3(n1169),.QN(n283));
  NAND3X0 U1872(.IN1(n1170),.IN2(n1171),.IN3(n1172),.QN(n274));
  NAND3X0 U1873(.IN1(n1173),.IN2(n1174),.IN3(n1175),.QN(n273));
  NAND2X1 U1874(.IN1(n1176),.IN2(n1177),.QN(n286));
  NAND2X1 U1875(.IN1(n1178),.IN2(n1179),.QN(n276));
  NBUFFX2 U1876(.INP(s_shr2[5:5]),.Z(n1283));
  NBUFFX2 U1877(.INP(s_shl2[5:5]),.Z(n1276));
  NBUFFX2 U1878(.INP(s_shl2[5:5]),.Z(n1275));
  NBUFFX2 U1879(.INP(s_shr2[5:5]),.Z(n1284));
  INVX0 U1880(.INP(n1718),.ZN(n1341));
  INVX0 U1881(.INP(n1686),.ZN(n1352));
  INVX0 U1882(.INP(n1726),.ZN(n1351));
  INVX0 U1883(.INP(n1734),.ZN(n1345));
  INVX0 U1884(.INP(n1702),.ZN(n1347));
  INVX0 U1885(.INP(n1742),.ZN(n1349));
  INVX0 U1886(.INP(n1748),.ZN(n1339));
  DELLN1X2 U1887(.INP(s_fract_48_i[12:12]),.Z(n1210));
  DELLN1X2 U1888(.INP(s_fract_48_i[12:12]),.Z(n1211));
  DELLN1X2 U1889(.INP(s_fract_48_i[30:30]),.Z(n1217));
  DELLN1X2 U1890(.INP(s_fract_48_i[30:30]),.Z(n1216));
  DELLN1X2 U1891(.INP(s_fract_48_i[18:18]),.Z(n1214));
  DELLN1X2 U1892(.INP(s_fract_48_i[18:18]),.Z(n1213));
  NBUFFX2 U1893(.INP(s_fract_48_i[18:18]),.Z(n1212));
  NBUFFX2 U1894(.INP(s_fract_48_i[30:30]),.Z(n1215));
  INVX0 U1895(.INP(n352),.ZN(n1466));
  INVX0 U1896(.INP(n715),.ZN(n1465));
  INVX0 U1897(.INP(n593),.ZN(n1451));
  NOR2X0 U1898(.IN1(n316),.IN2(n1330),.QN(n319));
  INVX0 U1899(.INP(n322),.ZN(n1330));
  NOR2X0 U1900(.IN1(n1329),.IN2(s_exp_10b[8:8]),.QN(n318));
  INVX0 U1901(.INP(n319),.ZN(n1329));
  INVX0 U1902(.INP(n448),.ZN(n1454));
  NOR2X0 U1903(.IN1(n250),.IN2(n1515),.QN(n263));
  INVX0 U1904(.INP(n450),.ZN(n1501));
  INVX0 U1905(.INP(n1708),.ZN(n1340));
  NAND2X0 U1906(.IN1(n1553),.IN2(n1235),.QN(n1629));
  INVX0 U1907(.INP(n1990),.ZN(n1492));
  INVX0 U1908(.INP(n1971),.ZN(n1498));
  NOR2X0 U1909(.IN1(n1689),.IN2(n1279),.QN(n1718));
  NOR2X0 U1910(.IN1(n1626),.IN2(n1279),.QN(n1686));
  NOR2X0 U1911(.IN1(n1690),.IN2(n1279),.QN(n1726));
  NOR2X0 U1912(.IN1(n1691),.IN2(n1279),.QN(n1734));
  NOR2X0 U1913(.IN1(n1688),.IN2(n1279),.QN(n1702));
  NOR2X0 U1914(.IN1(n1692),.IN2(n1280),.QN(n1742));
  NOR2X0 U1915(.IN1(n1704),.IN2(n1280),.QN(n1748));
  NOR2X0 U1916(.IN1(n316),.IN2(n322),.QN(n321));
  NAND2X0 U1917(.IN1(n1648),.IN2(n1232),.QN(n1704));
  INVX0 U1918(.INP(n1711),.ZN(n1348));
  INVX0 U1919(.INP(n1707),.ZN(n1346));
  INVX0 U1920(.INP(n1709),.ZN(n1350));
  INVX0 U1921(.INP(n1710),.ZN(n1344));
  INVX0 U1922(.INP(n1706),.ZN(n1342));
  INVX0 U1923(.INP(n1754),.ZN(n1353));
  INVX0 U1924(.INP(n1653),.ZN(n1405));
  INVX0 U1925(.INP(n1628),.ZN(n1390));
  INVX0 U1926(.INP(n1600),.ZN(n1386));
  NOR2X0 U1927(.IN1(n1677),.IN2(n1279),.QN(n1687));
  INVX0 U1928(.INP(n1929),.ZN(n1426));
  INVX0 U1929(.INP(n1938),.ZN(n1422));
  INVX0 U1930(.INP(n1947),.ZN(n1418));
  INVX0 U1931(.INP(n1956),.ZN(n1414));
  INVX0 U1932(.INP(n1777),.ZN(n1504));
  INVX0 U1933(.INP(n2000),.ZN(n1489));
  INVX0 U1934(.INP(n1980),.ZN(n1495));
  INVX0 U1935(.INP(n265),.ZN(n1335));
  INVX0 U1936(.INP(n1780),.ZN(n1509));
  INVX0 U1937(.INP(n1762),.ZN(n1503));
  INVX0 U1938(.INP(n1685),.ZN(n1337));
  INVX0 U1939(.INP(n1969),.ZN(n1459));
  INVX0 U1940(.INP(n1978),.ZN(n1457));
  INVX0 U1941(.INP(n1988),.ZN(n1452));
  INVX0 U1942(.INP(n1998),.ZN(n1448));
  NAND2X0 U1943(.IN1(n347),.IN2(n1026),.QN(n424));
  NAND2X0 U1944(.IN1(n372),.IN2(n1073),.QN(n365));
  NAND2X0 U1945(.IN1(n347),.IN2(n1025),.QN(n340));
  NAND2X0 U1946(.IN1(n612),.IN2(n1002),.QN(n605));
  AOI222X1 U1947(.IN1(n598),.IN2(n946),.IN3(n599),.IN4(n1018),.IN5(n600),.IN6(n1000),.QN(n1181));
  AND2X1 U1948(.IN1(n1182),.IN2(n1183),.Q(n615));
  AOI222X1 U1949(.IN1(n622),.IN2(n1079),.IN3(n1224),.IN4(n974),.IN5(n623),.IN6(n893),.QN(n1183));
  AOI221X2 U1950(.IN1(n1454),.IN2(N2081),.IN3(n1453),.IN4(n360),.IN5(n361),.QN(n1184));
  AOI222X1 U1951(.IN1(n358),.IN2(n1089),.IN3(n1289),.IN4(n1030),.IN5(n359),.IN6(N2033),.QN(n1185));
  HADDX1 U1952(.A0(N2351),.B0(\add_105_I48_L14036_C136/carry[3] ),.C1(\add_105_I48_L14036_C136/carry[4] ),.SO(N2361));
  INVX0 U1953(.INP(n942),.ZN(n1314));
  OAI22X1 U1954(.IN1(n1513),.IN2(n1186),.IN3(n452),.IN4(n331),.QN(N2976));
  AND4X1 U1955(.IN1(n453),.IN2(n456),.IN3(n455),.IN4(n454),.Q(n1186));
  INVX0 U1956(.INP(n331),.ZN(n1513));
  INVX0 U1957(.INP(n1037),.ZN(n1317));
  AND2X1 U1958(.IN1(n1187),.IN2(n1188),.Q(n375));
  AOI222X1 U1959(.IN1(n383),.IN2(n48),.IN3(n1228),.IN4(n52),.IN5(n384),.IN6(n29),.QN(n1188));
  OA21X1 U1960(.IN1(n418),.IN2(n419),.IN3(n331),.Q(N2977));
  NAND2X0 U1961(.IN1(n347),.IN2(n187),.QN(n397));
  NAND2X0 U1962(.IN1(n588),.IN2(n922),.QN(n638));
  NOR2X0 U1963(.IN1(n553),.IN2(n554),.QN(n552));
  INVX0 U1964(.INP(N2348),.ZN(N2358));
  NOR2X0 U1965(.IN1(n539),.IN2(n540),.QN(n534));
  AOI222X1 U1966(.IN1(n1078),.IN2(n387),.IN3(n32),.IN4(s_fract_48_i[36:36]),.IN5(n700),.IN6(n388),.QN(n412));
  INVX0 U1967(.INP(n1095),.ZN(n1318));
  AOI21X1 U1968(.IN1(n1189),.IN2(n1190),.IN3(n573),.QN(N1636));
  AOI222X1 U1969(.IN1(n578),.IN2(n1006),.IN3(n635),.IN4(N366),.IN5(n1387),.IN6(n636),.QN(n1189));
  NAND2X0 U1970(.IN1(n612),.IN2(n613),.QN(n676));
  AND2X1 U1971(.IN1(n1191),.IN2(n1192),.Q(n741));
  AO22X1 U1972(.IN1(n611),.IN2(n1043),.IN3(n1214),.IN4(n997),.Q(n737));
  INVX0 U1973(.INP(n180),.ZN(n1361));
  INVX0 U1974(.INP(n486),.ZN(n1363));
  OA21X1 U1975(.IN1(n659),.IN2(n660),.IN3(n661),.Q(N1635));
  NAND2X0 U1976(.IN1(n1451),.IN2(N634),.QN(n762));
  NAND2X0 U1977(.IN1(n612),.IN2(n220),.QN(n704));
  NAND2X0 U1978(.IN1(n588),.IN2(n820),.QN(n691));
  NOR2X0 U1979(.IN1(n775),.IN2(n776),.QN(n771));
  NOR2X0 U1980(.IN1(n791),.IN2(n792),.QN(n790));
  INVX0 U1981(.INP(N1025),.ZN(N1036));
  INVX0 U1982(.INP(n848),.ZN(n1366));
  INVX0 U1983(.INP(n1031),.ZN(n1370));
  OA21X1 U1984(.IN1(n685),.IN2(n686),.IN3(n661),.Q(N1634));
  INVX0 U1985(.INP(N2270),.ZN(n1397));
  INVX0 U1986(.INP(n926),.ZN(n1320));
  INVX0 U1987(.INP(n1027),.ZN(n1311));
  INVX0 U1988(.INP(n107),.ZN(n1404));
  INVX0 U1989(.INP(n1009),.ZN(n1312));
  INVX0 U1990(.INP(n1047),.ZN(n1325));
  INVX0 U1991(.INP(N941),.ZN(n1371));
  INVX0 U1992(.INP(n184),.ZN(n1409));
  INVX0 U1993(.INP(n1021),.ZN(n1321));
  INVX0 U1994(.INP(n1096),.ZN(n1358));
  INVX0 U1995(.INP(N2237),.ZN(n1410));
  INVX0 U1996(.INP(n1093),.ZN(n1364));
  INVX0 U1997(.INP(N924),.ZN(n1372));
  INVX0 U1998(.INP(n818),.ZN(n1313));
  INVX0 U1999(.INP(n1103),.ZN(n1359));
  INVX0 U2000(.INP(N906),.ZN(n1379));
  INVX0 U2001(.INP(n166),.ZN(n1373));
  INVX0 U2002(.INP(n847),.ZN(n1360));
  INVX0 U2003(.INP(n239),.ZN(n1365));
  INVX0 U2004(.INP(n216),.ZN(n1374));
  INVX0 U2005(.INP(n915),.ZN(n1456));
  INVX0 U2006(.INP(n237),.ZN(n1375));
  NAND2X0 U2007(.IN1(n1466),.IN2(N1980),.QN(n525));
  INVX0 U2008(.INP(n805),.ZN(n1467));
  INVX0 U2009(.INP(n943),.ZN(n1322));
  INVX0 U2010(.INP(N1949),.ZN(n1476));
  INVX0 U2011(.INP(n1041),.ZN(n1471));
  INVX0 U2012(.INP(N1953),.ZN(n1323));
  INVX0 U2013(.INP(n188),.ZN(n1475));
  INVX0 U2014(.INP(n1059),.ZN(n1470));
  INVX0 U2015(.INP(n982),.ZN(n1315));
  INVX0 U2016(.INP(N1964),.ZN(n1472));
  INVX0 U2017(.INP(n190),.ZN(n1474));
  INVX0 U2018(.INP(n1084),.ZN(n1316));
  INVX0 U2019(.INP(n433),.ZN(n1367));
  INVX0 U2020(.INP(n994),.ZN(n1376));
  INVX0 U2021(.INP(N617),.ZN(n1380));
  INVX0 U2022(.INP(n983),.ZN(n1319));
  INVX0 U2023(.INP(n984),.ZN(n1362));
  INVX0 U2024(.INP(n404),.ZN(n1368));
  INVX0 U2025(.INP(n1068),.ZN(n1377));
  INVX0 U2026(.INP(n1028),.ZN(n1369));
  INVX0 U2027(.INP(n930),.ZN(n1378));
  NAND2X0 U2028(.IN1(n588),.IN2(n865),.QN(n581));
  NOR2X0 U2029(.IN1(n1481),.IN2(n709),.QN(n612));
  INVX0 U2030(.INP(n779),.ZN(n1481));
  INVX0 U2031(.INP(n778),.ZN(n1482));
  INVX0 U2032(.INP(n777),.ZN(n1483));
  INVX0 U2033(.INP(n782),.ZN(n1484));
  NAND2X0 U2034(.IN1(n588),.IN2(n1087),.QN(n664));
  NOR2X0 U2035(.IN1(n1439),.IN2(n442),.QN(n372));
  INVX0 U2036(.INP(n545),.ZN(n1443));
  INVX0 U2037(.INP(n546),.ZN(n1439));
  INVX0 U2038(.INP(n541),.ZN(n1447));
  INVX0 U2039(.INP(n542),.ZN(n1450));
  NOR2X0 U2040(.IN1(n1428),.IN2(n696),.QN(n588));
  INVX0 U2041(.INP(n756),.ZN(n1429));
  INVX0 U2042(.INP(n755),.ZN(n1430));
  INVX0 U2043(.INP(n757),.ZN(n1428));
  INVX0 U2044(.INP(n760),.ZN(n1431));
  INVX0 U2045(.INP(n709),.ZN(n1480));
  NOR2X0 U2046(.IN1(n1482),.IN2(n779),.QN(n610));
  NOR2X0 U2047(.IN1(n1443),.IN2(n546),.QN(n371));
  INVX0 U2048(.INP(n696),.ZN(n1427));
  INVX0 U2049(.INP(n442),.ZN(n1435));
  NOR2X0 U2050(.IN1(n1488),.IN2(n429),.QN(n347));
  INVX0 U2051(.INP(n523),.ZN(n1488));
  INVX0 U2052(.INP(n522),.ZN(n1491));
  INVX0 U2053(.INP(n518),.ZN(n1494));
  INVX0 U2054(.INP(n519),.ZN(n1497));
  NOR2X0 U2055(.IN1(n1483),.IN2(n778),.QN(n609));
  NOR2X0 U2056(.IN1(n1429),.IN2(n757),.QN(n586));
  NOR2X0 U2057(.IN1(n1447),.IN2(n545),.QN(n370));
  NOR2X0 U2058(.IN1(n795),.IN2(n624),.QN(n626));
  NOR2X0 U2059(.IN1(n1491),.IN2(n523),.QN(n346));
  INVX0 U2060(.INP(n429),.ZN(n1486));
  NOR2X0 U2061(.IN1(n556),.IN2(n557),.QN(n385));
  NOR2X0 U2062(.IN1(n1430),.IN2(n756),.QN(n585));
  NOR2X0 U2063(.IN1(n1450),.IN2(n541),.QN(n368));
  NOR2X0 U2064(.IN1(n1484),.IN2(n777),.QN(n608));
  INVX0 U2065(.INP(n558),.ZN(n1336));
  NAND2X1 U2066(.IN1(n774),.IN2(n714),.QN(n715));
  NOR2X0 U2067(.IN1(n323),.IN2(s_exp_10b[9:9]),.QN(n322));
  NOR2X0 U2068(.IN1(n793),.IN2(n794),.QN(n623));
  NOR2X0 U2069(.IN1(n1494),.IN2(n522),.QN(n345));
  NAND2X1 U2070(.IN1(n537),.IN2(n447),.QN(n448));
  INVX0 U2071(.INP(n714),.ZN(n1464));
  INVX0 U2072(.INP(N3347),.ZN(n1332));
  NAND2X0 U2073(.IN1(N3349),.IN2(N3348),.QN(n298));
  NAND2X0 U2074(.IN1(n1335),.IN2(n258),.QN(n250));
  NOR2X0 U2075(.IN1(n782),.IN2(n1212),.QN(n611));
  NOR2X0 U2076(.IN1(n796),.IN2(n774),.QN(n598));
  NOR2X0 U2077(.IN1(n536),.IN2(n537),.QN(n362));
  NOR2X0 U2078(.IN1(n1431),.IN2(n755),.QN(n584));
  INVX0 U2079(.INP(n447),.ZN(n1453));
  INVX0 U2080(.INP(n1197),.ZN(n1331));
  NOR2X0 U2081(.IN1(n542),.IN2(n1215),.QN(n369));
  NOR2X0 U2082(.IN1(n555),.IN2(n1228),.QN(n383));
  NOR2X0 U2083(.IN1(n1221),.IN2(n1224),.QN(n565));
  NOR2X0 U2084(.IN1(n1497),.IN2(n518),.QN(n343));
  NOR2X0 U2085(.IN1(n550),.IN2(n551),.QN(n387));
  INVX0 U2086(.INP(n752),.ZN(n1388));
  INVX0 U2087(.INP(n751),.ZN(n1387));
  NOR2X0 U2088(.IN1(n1663),.IN2(n1279),.QN(n1708));
  NBUFFX4 U2089(.INP(n71),.Z(n1235));
  NOR2X0 U2090(.IN1(n760),.IN2(s_fract_48_i[36:36]),.QN(n587));
  NOR2X0 U2091(.IN1(n1856),.IN2(n1272),.QN(n1990));
  NOR2X0 U2092(.IN1(n1845),.IN2(n1272),.QN(n1971));
  NOR2X0 U2093(.IN1(n798),.IN2(n750),.QN(n575));
  NOR2X0 U2094(.IN1(n563),.IN2(n562),.QN(n337));
  INVX0 U2095(.INP(n449),.ZN(n1500));
  NOR2X0 U2096(.IN1(n1285),.IN2(n1340),.QN(N3137));
  NOR2X0 U2097(.IN1(n1277),.IN2(n1492),.QN(N3155));
  NOR2X0 U2098(.IN1(n1277),.IN2(n1498),.QN(N3153));
  NOR2X0 U2099(.IN1(n1683),.IN2(n1279),.QN(n1711));
  NOR2X0 U2100(.IN1(n1660),.IN2(n1279),.QN(n1707));
  NOR2X0 U2101(.IN1(n1666),.IN2(n1279),.QN(n1709));
  NOR2X0 U2102(.IN1(n1680),.IN2(n1279),.QN(n1710));
  NOR2X0 U2103(.IN1(n1657),.IN2(n1279),.QN(n1706));
  NBUFFX4 U2104(.INP(n72),.Z(n1241));
  NBUFFX4 U2105(.INP(n72),.Z(n1240));
  NOR2X0 U2106(.IN1(n1705),.IN2(n1280),.QN(n1754));
  NBUFFX4 U2107(.INP(n71),.Z(n1236));
  AO21X1 U2108(.IN1(n326),.IN2(n327),.IN3(s_exp_10a[9:9]),.Q(n316));
  NOR2X0 U2109(.IN1(n773),.IN2(n797),.QN(n600));
  NOR2X0 U2110(.IN1(n561),.IN2(n538),.QN(n359));
  NAND2X1 U2111(.IN1(n529),.IN2(n530),.QN(n354));
  NAND2X0 U2112(.IN1(n1540),.IN2(n1237),.QN(n1584));
  INVX0 U2113(.INP(n299),.ZN(n1257));
  INVX0 U2114(.INP(n1614),.ZN(n1394));
  INVX0 U2115(.INP(n1633),.ZN(n1385));
  INVX0 U2116(.INP(n1638),.ZN(n1383));
  INVX0 U2117(.INP(n1643),.ZN(n1356));
  NAND2X1 U2118(.IN1(n767),.IN2(n765),.QN(n631));
  XNOR2X1 U2119(.IN1(n1285),.IN2(n1193),.Q(N3243));
  NAND2X0 U2120(.IN1(\add_197/carry[4] ),.IN2(n1280),.QN(n1193));
  INVX0 U2121(.INP(n1746),.ZN(n1411));
  INVX0 U2122(.INP(n1752),.ZN(n1406));
  INVX0 U2123(.INP(n1732),.ZN(n1419));
  INVX0 U2124(.INP(n1716),.ZN(n1432));
  INVX0 U2125(.INP(n1724),.ZN(n1423));
  INVX0 U2126(.INP(n1740),.ZN(n1415));
  INVX0 U2127(.INP(n1700),.ZN(n1436));
  INVX0 U2128(.INP(n1679),.ZN(n1382));
  INVX0 U2129(.INP(n1656),.ZN(n1398));
  INVX0 U2130(.INP(n1676),.ZN(n1440));
  INVX0 U2131(.INP(n1662),.ZN(n1389));
  INVX0 U2132(.INP(n1625),.ZN(n1444));
  INVX0 U2133(.INP(n1665),.ZN(n1384));
  INVX0 U2134(.INP(n1659),.ZN(n1393));
  INVX0 U2135(.INP(n1572),.ZN(n1357));
  INVX0 U2136(.INP(n1948),.ZN(n1396));
  INVX0 U2137(.INP(n1926),.ZN(n1412));
  NOR2X0 U2138(.IN1(n1285),.IN2(n1349),.QN(N3132));
  NOR2X0 U2139(.IN1(n1285),.IN2(n1348),.QN(N3140));
  INVX0 U2140(.INP(n1963),.ZN(n1391));
  NOR2X0 U2141(.IN1(n1285),.IN2(n1346),.QN(N3136));
  NOR2X0 U2142(.IN1(n1285),.IN2(n1350),.QN(N3138));
  INVX0 U2143(.INP(n1945),.ZN(n1400));
  NOR2X0 U2144(.IN1(n1285),.IN2(n1353),.QN(N3134));
  NOR2X0 U2145(.IN1(n1285),.IN2(n1344),.QN(N3139));
  INVX0 U2146(.INP(n1954),.ZN(n1395));
  NOR2X0 U2147(.IN1(n1285),.IN2(n1342),.QN(N3135));
  INVX0 U2148(.INP(n1902),.ZN(n1424));
  NOR2X0 U2149(.IN1(n1284),.IN2(n1341),.QN(N3129));
  INVX0 U2150(.INP(n1878),.ZN(n1441));
  NOR2X0 U2151(.IN1(n1284),.IN2(n1352),.QN(N3126));
  INVX0 U2152(.INP(n1910),.ZN(n1420));
  NOR2X0 U2153(.IN1(n1284),.IN2(n1351),.QN(N3130));
  INVX0 U2154(.INP(n1918),.ZN(n1416));
  NOR2X0 U2155(.IN1(n1284),.IN2(n1345),.QN(N3131));
  NOR2X0 U2156(.IN1(n1275),.IN2(n1857),.QN(N3171));
  NOR2X0 U2157(.IN1(n1284),.IN2(n1681),.QN(N3123));
  NOR2X0 U2158(.IN1(n1276),.IN2(n1836),.QN(N3167));
  NOR2X0 U2159(.IN1(n1283),.IN2(n1658),.QN(N3119));
  INVX0 U2160(.INP(n1894),.ZN(n1433));
  NOR2X0 U2161(.IN1(n1284),.IN2(n1347),.QN(N3128));
  NOR2X0 U2162(.IN1(n1276),.IN2(n1815),.QN(N3163));
  NOR2X0 U2163(.IN1(n1283),.IN2(n1642),.QN(N3115));
  NOR2X0 U2164(.IN1(n1276),.IN2(n1795),.QN(N3159));
  NOR2X0 U2165(.IN1(n1283),.IN2(n1613),.QN(N3111));
  NOR2X0 U2166(.IN1(n1275),.IN2(n1846),.QN(N3169));
  NOR2X0 U2167(.IN1(n1284),.IN2(n1664),.QN(N3121));
  NOR2X0 U2168(.IN1(n1277),.IN2(n1786),.QN(N3157));
  NOR2X0 U2169(.IN1(n1283),.IN2(n1338),.QN(N3109));
  INVX0 U2170(.INP(n1936),.ZN(n1407));
  NOR2X0 U2171(.IN1(n1284),.IN2(n1339),.QN(N3133));
  NOR2X0 U2172(.IN1(n1276),.IN2(n1805),.QN(N3161));
  NOR2X0 U2173(.IN1(n1283),.IN2(n1632),.QN(N3113));
  NOR2X0 U2174(.IN1(n1276),.IN2(n1790),.QN(N3158));
  NOR2X0 U2175(.IN1(n1283),.IN2(n1608),.QN(N3110));
  NOR2X0 U2176(.IN1(n1275),.IN2(n1851),.QN(N3170));
  NOR2X0 U2177(.IN1(n1284),.IN2(n1667),.QN(N3122));
  NOR2X0 U2178(.IN1(n1276),.IN2(n1825),.QN(N3165));
  NOR2X0 U2179(.IN1(n1283),.IN2(n1651),.QN(N3117));
  NOR2X0 U2180(.IN1(n1276),.IN2(n1810),.QN(N3162));
  NOR2X0 U2181(.IN1(n1283),.IN2(n1637),.QN(N3114));
  NOR2X0 U2182(.IN1(n1276),.IN2(n1831),.QN(N3166));
  NOR2X0 U2183(.IN1(n1283),.IN2(n1655),.QN(N3118));
  NOR2X0 U2184(.IN1(n1276),.IN2(n1819),.QN(N3164));
  NOR2X0 U2185(.IN1(n1283),.IN2(n1647),.QN(N3116));
  NOR2X0 U2186(.IN1(n1276),.IN2(n1841),.QN(N3168));
  NOR2X0 U2187(.IN1(n1283),.IN2(n1661),.QN(N3120));
  NOR2X0 U2188(.IN1(n1276),.IN2(n1799),.QN(N3160));
  NOR2X0 U2189(.IN1(n1283),.IN2(n1618),.QN(N3112));
  INVX0 U2190(.INP(n1599),.ZN(n1338));
  INVX0 U2191(.INP(N3240),.ZN(n1310));
  NBUFFX4 U2192(.INP(n77),.Z(n1233));
  NBUFFX4 U2193(.INP(n73),.Z(n1238));
  NBUFFX4 U2194(.INP(n77),.Z(n1232));
  NBUFFX4 U2195(.INP(n73),.Z(n1237));
  NBUFFX2 U2196(.INP(n73),.Z(n1239));
  NOR2X0 U2197(.IN1(n519),.IN2(n1209),.QN(n344));
  NOR2X0 U2198(.IN1(n1861),.IN2(n1272),.QN(n2000));
  NOR2X0 U2199(.IN1(n1850),.IN2(n1272),.QN(n1980));
  NOR2X0 U2200(.IN1(n1388),.IN2(n799),.QN(n574));
  NOR2X0 U2201(.IN1(n566),.IN2(n564),.QN(n334));
  NOR2X0 U2202(.IN1(n528),.IN2(n529),.QN(n389));
  INVX0 U2203(.INP(n299),.ZN(n1259));
  INVX0 U2204(.INP(n299),.ZN(n1258));
  INVX0 U2205(.INP(n1609),.ZN(n1399));
  NAND2X1 U2206(.IN1(n1598),.IN2(n79),.QN(n1685));
  INVX0 U2207(.INP(n1895),.ZN(n1438));
  INVX0 U2208(.INP(n1903),.ZN(n1434));
  INVX0 U2209(.INP(n1765),.ZN(n1505));
  INVX0 U2210(.INP(n1682),.ZN(n1355));
  INVX0 U2211(.INP(n1758),.ZN(n1510));
  NAND2X1 U2212(.IN1(n1772),.IN2(n53),.QN(n1789));
  NAND2X0 U2213(.IN1(n1778),.IN2(n56),.QN(n1798));
  INVX0 U2214(.INP(n1930),.ZN(n1408));
  INVX0 U2215(.INP(n1939),.ZN(n1401));
  NAND2X1 U2216(.IN1(n254),.IN2(n252),.QN(n265));
  NOR2X0 U2217(.IN1(n1284),.IN2(n1343),.QN(N3127));
  INVX0 U2218(.INP(n1886),.ZN(n1437));
  INVX0 U2219(.INP(n1687),.ZN(n1343));
  NOR2X0 U2220(.IN1(n1284),.IN2(n1685),.QN(N3125));
  INVX0 U2221(.INP(n1870),.ZN(n1445));
  NOR2X0 U2222(.IN1(n1275),.IN2(n1862),.QN(N3172));
  NOR2X0 U2223(.IN1(n1284),.IN2(n1684),.QN(N3124));
  NOR2X0 U2224(.IN1(n1275),.IN2(n2002),.QN(N3145));
  NOR2X0 U2225(.IN1(n1277),.IN2(n1489),.QN(N3156));
  NOR2X0 U2226(.IN1(n1277),.IN2(n1495),.QN(N3154));
  NOR2X0 U2227(.IN1(n1276),.IN2(n1876),.QN(N3142));
  NOR2X0 U2228(.IN1(n1277),.IN2(n1868),.QN(N3141));
  NOR2X0 U2229(.IN1(n1275),.IN2(n1884),.QN(N3143));
  NOR2X0 U2230(.IN1(n1275),.IN2(n1927),.QN(N3144));
  NOR2X0 U2231(.IN1(n1275),.IN2(n2003),.QN(N3146));
  NOR2X0 U2232(.IN1(n1275),.IN2(n2004),.QN(N3147));
  NOR2X0 U2233(.IN1(n1277),.IN2(n1952),.QN(N3151));
  NOR2X0 U2234(.IN1(n1277),.IN2(n1961),.QN(N3152));
  NOR2X0 U2235(.IN1(n1275),.IN2(n2005),.QN(N3148));
  NOR2X0 U2236(.IN1(n1275),.IN2(n2007),.QN(N3150));
  NOR2X0 U2237(.IN1(n1275),.IN2(n2006),.QN(N3149));
  INVX0 U2238(.INP(n1967),.ZN(n1425));
  INVX0 U2239(.INP(n1976),.ZN(n1421));
  INVX0 U2240(.INP(n1986),.ZN(n1417));
  INVX0 U2241(.INP(n1996),.ZN(n1413));
  INVX0 U2242(.INP(n1768),.ZN(n1507));
  INVX0 U2243(.INP(n1771),.ZN(n1511));
  INVX0 U2244(.INP(n260),.ZN(n1334));
  NOR2X0 U2245(.IN1(n261),.IN2(n262),.QN(n251));
  OA21X1 U2246(.IN1(n1333),.IN2(n254),.IN3(n255),.Q(n253));
  NBUFFX2 U2247(.INP(n72),.Z(n1242));
  NBUFFX2 U2248(.INP(n1204),.Z(n1247));
  INVX0 U2249(.INP(s_exp_10a[0:0]),.ZN(n1293));
  INVX0 U2250(.INP(n1957),.ZN(n1392));
  XOR2X1 U2251(.IN1(s_exp_10a[6:6]),.IN2(n1194),.Q(N3005));
  NAND2X1 U2252(.IN1(\sub_0_root_add_0_root_add_148/carry[5] ),.IN2(n1298),.QN(n1194));
  NBUFFX2 U2253(.INP(n1204),.Z(n1253));
  NBUFFX2 U2254(.INP(n1204),.Z(n1252));
  NBUFFX2 U2255(.INP(n1204),.Z(n1251));
  NBUFFX2 U2256(.INP(n1204),.Z(n1250));
  NBUFFX2 U2257(.INP(n1204),.Z(n1249));
  NBUFFX2 U2258(.INP(n1204),.Z(n1248));
  NOR2X0 U2259(.IN1(n687),.IN2(n752),.QN(n635));
  NBUFFX2 U2260(.INP(n1204),.Z(n1254));
  INVX0 U2261(.INP(s_exp_10a[2:2]),.ZN(n1295));
  INVX0 U2262(.INP(s_exp_10a[4:4]),.ZN(n1297));
  INVX0 U2263(.INP(s_exp_10a[3:3]),.ZN(n1296));
  INVX0 U2264(.INP(s_exp_10a[5:5]),.ZN(n1298));
  INVX0 U2265(.INP(n257),.ZN(n1515));
  NOR2X0 U2266(.IN1(n565),.IN2(n1220),.QN(n333));
  NBUFFX2 U2267(.INP(n77),.Z(n1234));
  INVX0 U2268(.INP(n259),.ZN(n1333));
  INVX0 U2269(.INP(N583),.ZN(N594));
  INVX0 U2270(.INP(N1932),.ZN(N1942));
  INVX0 U2271(.INP(N889),.ZN(N900));
  INVX0 U2272(.INP(N2220),.ZN(N2230));
  INVX0 U2273(.INP(N719),.ZN(N730));
  INVX0 U2274(.INP(N923),.ZN(N934));
  INVX0 U2275(.INP(N1772),.ZN(N1782));
  INVX0 U2276(.INP(N2060),.ZN(N2070));
  INVX0 U2277(.INP(N2236),.ZN(N2246));
  INVX0 U2278(.INP(N2252),.ZN(N2262));
  INVX0 U2279(.INP(N566),.ZN(N577));
  INVX0 U2280(.INP(N872),.ZN(N883));
  INVX0 U2281(.INP(N600),.ZN(N611));
  INVX0 U2282(.INP(N1948),.ZN(N1958));
  INVX0 U2283(.INP(N1996),.ZN(N2006));
  INVX0 U2284(.INP(N2188),.ZN(N2198));
  INVX0 U2285(.INP(N413),.ZN(N424));
  INVX0 U2286(.INP(N2012),.ZN(N2022));
  INVX0 U2287(.INP(N991),.ZN(N1002));
  INVX0 U2288(.INP(N2028),.ZN(N2038));
  INVX0 U2289(.INP(N685),.ZN(N696));
  INVX0 U2290(.INP(N2300),.ZN(N2310));
  INVX0 U2291(.INP(N481),.ZN(N492));
  INVX0 U2292(.INP(N787),.ZN(N798));
  INVX0 U2293(.INP(N1820),.ZN(N1830));
  INVX0 U2294(.INP(N770),.ZN(N781));
  INVX0 U2295(.INP(N2108),.ZN(N2118));
  INVX0 U2296(.INP(N2316),.ZN(N2326));
  INVX0 U2297(.INP(N2268),.ZN(N2278));
  INVX0 U2298(.INP(N1788),.ZN(N1798));
  INVX0 U2299(.INP(N2076),.ZN(N2086));
  INVX0 U2300(.INP(N940),.ZN(N951));
  INVX0 U2301(.INP(N1708),.ZN(N1718));
  INVX0 U2302(.INP(N549),.ZN(N560));
  INVX0 U2303(.INP(N855),.ZN(N866));
  INVX0 U2304(.INP(N651),.ZN(N662));
  INVX0 U2305(.INP(N974),.ZN(N985));
  INVX0 U2306(.INP(N396),.ZN(N407));
  INVX0 U2307(.INP(N702),.ZN(N713));
  INVX0 U2308(.INP(N1836),.ZN(N1846));
  INVX0 U2309(.INP(N2124),.ZN(N2134));
  INVX0 U2310(.INP(N1980),.ZN(N1990));
  INVX0 U2311(.INP(N634),.ZN(N645));
  INVX0 U2312(.INP(N1884),.ZN(N1894));
  INVX0 U2313(.INP(N2172),.ZN(N2182));
  INVX0 U2314(.INP(N430),.ZN(N441));
  INVX0 U2315(.INP(N736),.ZN(N747));
  INVX0 U2316(.INP(N2284),.ZN(N2294));
  INVX0 U2317(.INP(N2156),.ZN(N2166));
  INVX0 U2318(.INP(N515),.ZN(N526));
  INVX0 U2319(.INP(N821),.ZN(N832));
  INVX0 U2320(.INP(N1756),.ZN(N1766));
  INVX0 U2321(.INP(N2044),.ZN(N2054));
  INVX0 U2322(.INP(N498),.ZN(N509));
  INVX0 U2323(.INP(N2092),.ZN(N2102));
  INVX0 U2324(.INP(N804),.ZN(N815));
  INVX0 U2325(.INP(N447),.ZN(N458));
  INVX0 U2326(.INP(N2204),.ZN(N2214));
  INVX0 U2327(.INP(N1852),.ZN(N1862));
  INVX0 U2328(.INP(N753),.ZN(N764));
  INVX0 U2329(.INP(N2140),.ZN(N2150));
  INVX0 U2330(.INP(N1916),.ZN(N1926));
  INVX0 U2331(.INP(N668),.ZN(N679));
  INVX0 U2332(.INP(N957),.ZN(N968));
  INVX0 U2333(.INP(N1724),.ZN(N1734));
  INVX0 U2334(.INP(N1692),.ZN(N1702));
  INVX0 U2335(.INP(N532),.ZN(N543));
  INVX0 U2336(.INP(N838),.ZN(N849));
  INVX0 U2337(.INP(N1008),.ZN(N1019));
  AND2X1 U2338(.IN1(N1707),.IN2(n226),.Q(n1195));
  INVX0 U2339(.INP(N1804),.ZN(N1814));
  INVX0 U2340(.INP(N362),.ZN(N373));
  INVX0 U2341(.INP(N379),.ZN(N390));
  INVX0 U2342(.INP(N1900),.ZN(N1910));
  INVX0 U2343(.INP(N464),.ZN(N475));
  INVX0 U2344(.INP(N1868),.ZN(N1878));
  INVX0 U2345(.INP(N1740),.ZN(N1750));
  INVX0 U2346(.INP(N1677),.ZN(N1686));
  INVX0 U2347(.INP(N346),.ZN(N356));
  INVX0 U2348(.INP(N332),.ZN(N341));
  INVX0 U2349(.INP(N1664),.ZN(N1672));
  NAND2X0 U2350(.IN1(n719),.IN2(n720),.QN(n717));
  NOR2X0 U2351(.IN1(N2993),.IN2(n1205),.QN(n744));
  NAND2X0 U2352(.IN1(n747),.IN2(n748),.QN(n746));
  INVX0 U2353(.INP(s_fract_48_i[24:24]),.ZN(n1291));
  NOR2X0 U2354(.IN1(n1481),.IN2(s_fract_48_i[13:13]),.QN(n709));
  NOR2X0 U2355(.IN1(n1482),.IN2(s_fract_48_i[14:14]),.QN(n779));
  NOR2X0 U2356(.IN1(n1483),.IN2(s_fract_48_i[15:15]),.QN(n778));
  NOR2X0 U2357(.IN1(n1484),.IN2(s_fract_48_i[16:16]),.QN(n777));
  NOR2X0 U2358(.IN1(s_fract_48_i[17:17]),.IN2(n1212),.QN(n782));
  NOR2X0 U2359(.IN1(n1439),.IN2(s_fract_48_i[35:35]),.QN(n442));
  NOR2X0 U2360(.IN1(n1447),.IN2(s_fract_48_i[33:33]),.QN(n545));
  NOR2X0 U2361(.IN1(n1443),.IN2(s_fract_48_i[34:34]),.QN(n546));
  NOR2X0 U2362(.IN1(n1450),.IN2(s_fract_48_i[32:32]),.QN(n541));
  NOR2X0 U2363(.IN1(n1215),.IN2(s_fract_48_i[31:31]),.QN(n542));
  NOR2X0 U2364(.IN1(n1428),.IN2(s_fract_48_i[31:31]),.QN(n696));
  NOR2X0 U2365(.IN1(n1430),.IN2(s_fract_48_i[33:33]),.QN(n756));
  NOR2X0 U2366(.IN1(n1431),.IN2(s_fract_48_i[34:34]),.QN(n755));
  NOR2X0 U2367(.IN1(n1429),.IN2(s_fract_48_i[32:32]),.QN(n757));
  NOR2X0 U2368(.IN1(s_fract_48_i[35:35]),.IN2(s_fract_48_i[36:36]),.QN(n760));
  NOR2X0 U2369(.IN1(n1488),.IN2(s_fract_48_i[17:17]),.QN(n429));
  NOR2X0 U2370(.IN1(n1491),.IN2(s_fract_48_i[16:16]),.QN(n523));
  NOR2X0 U2371(.IN1(n1494),.IN2(s_fract_48_i[15:15]),.QN(n522));
  NOR2X0 U2372(.IN1(n1497),.IN2(s_fract_48_i[14:14]),.QN(n518));
  NOR2X0 U2373(.IN1(n1209),.IN2(s_fract_48_i[13:13]),.QN(n519));
  NOR2X0 U2374(.IN1(n550),.IN2(s_fract_48_i[38:38]),.QN(n551));
  NOR2X0 U2375(.IN1(n786),.IN2(s_fract_48_i[8:8]),.QN(n787));
  NOR2X0 U2376(.IN1(n789),.IN2(s_fract_48_i[10:10]),.QN(n788));
  NOR2X0 U2377(.IN1(n560),.IN2(s_fract_48_i[40:40]),.QN(n559));
  NOR2X0 U2378(.IN1(n793),.IN2(s_fract_48_i[4:4]),.QN(n794));
  NAND2X0 U2379(.IN1(n787),.IN2(n225),.QN(n616));
  NAND2X0 U2380(.IN1(n559),.IN2(n130),.QN(n376));
  NAND2X0 U2381(.IN1(n551),.IN2(n144),.QN(n560));
  NAND2X0 U2382(.IN1(n788),.IN2(n223),.QN(n786));
  NAND2X0 U2383(.IN1(n152),.IN2(n146),.QN(n550));
  NAND2X0 U2384(.IN1(n227),.IN2(n226),.QN(n793));
  NAND2X0 U2385(.IN1(n794),.IN2(n231),.QN(n795));
  NAND2X0 U2386(.IN1(n221),.IN2(n215),.QN(n789));
  NOR2X0 U2387(.IN1(n796),.IN2(s_fract_48_i[20:20]),.QN(n774));
  NOR2X0 U2388(.IN1(n528),.IN2(s_fract_48_i[20:20]),.QN(n529));
  NOR2X0 U2389(.IN1(n765),.IN2(s_fract_48_i[26:26]),.QN(n766));
  NOR2X0 U2390(.IN1(n530),.IN2(s_fract_48_i[22:22]),.QN(n531));
  NOR2X0 U2391(.IN1(n768),.IN2(s_fract_48_i[28:28]),.QN(n767));
  NOR2X0 U2392(.IN1(n773),.IN2(s_fract_48_i[22:22]),.QN(n797));
  NAND2X0 U2393(.IN1(n531),.IN2(n182),.QN(n351));
  NOR2X0 U2394(.IN1(n1229),.IN2(s_fract_48_i[43:43]),.QN(n555));
  NAND2X0 U2395(.IN1(n766),.IN2(n174),.QN(n592));
  NAND2X0 U2396(.IN1(n767),.IN2(n172),.QN(n765));
  NAND2X0 U2397(.IN1(n529),.IN2(n196),.QN(n530));
  NAND2X0 U2398(.IN1(n797),.IN2(n196),.QN(n796));
  NAND2X0 U2399(.IN1(n204),.IN2(n198),.QN(n528));
  NAND2X0 U2400(.IN1(n774),.IN2(n198),.QN(n714));
  NOR2X0 U2401(.IN1(n556),.IN2(s_fract_48_i[45:45]),.QN(n557));
  NAND2X0 U2402(.IN1(n555),.IN2(n47),.QN(n556));
  NAND2X0 U2403(.IN1(n182),.IN2(n177),.QN(n773));
  NAND2X0 U2404(.IN1(n170),.IN2(n164),.QN(n768));
  NOR2X0 U2405(.IN1(n536),.IN2(s_fract_48_i[28:28]),.QN(n537));
  NOR2X0 U2406(.IN1(n561),.IN2(s_fract_48_i[26:26]),.QN(n538));
  NAND2X0 U2407(.IN1(n537),.IN2(n170),.QN(n447));
  NAND2X0 U2408(.IN1(n538),.IN2(n172),.QN(n536));
  NAND2X0 U2409(.IN1(n177),.IN2(n174),.QN(n561));
  AND2X1 U2410(.IN1(n263),.IN2(s_frac_rnd[24:24]),.Q(n246));
  NOR2X0 U2411(.IN1(s_expo1[7:7]),.IN2(\sub_192_aco/carry[7] ),.QN(n1197));
  NOR2X0 U2412(.IN1(n563),.IN2(s_fract_48_i[10:10]),.QN(n562));
  NOR2X0 U2413(.IN1(n566),.IN2(s_fract_48_i[8:8]),.QN(n564));
  NOR2X0 U2414(.IN1(n798),.IN2(s_fract_48_i[38:38]),.QN(n750));
  NOR2X0 U2415(.IN1(n1388),.IN2(s_fract_48_i[40:40]),.QN(n799));
  NAND2X0 U2416(.IN1(n562),.IN2(n221),.QN(n449));
  NOR2X0 U2417(.IN1(n687),.IN2(s_fract_48_i[41:41]),.QN(n752));
  NAND2X0 U2418(.IN1(n799),.IN2(n144),.QN(n798));
  NAND2X0 U2419(.IN1(n564),.IN2(n223),.QN(n563));
  NAND2X0 U2420(.IN1(n565),.IN2(n225),.QN(n566));
  NAND2X0 U2421(.IN1(n123),.IN2(n122),.QN(n687));
  AND2X1 U2422(.IN1(n263),.IN2(n244),.Q(n1218));
  AND2X1 U2423(.IN1(n263),.IN2(n244),.Q(n247));
  AND2X1 U2424(.IN1(n263),.IN2(n244),.Q(n1219));
  NAND2X0 U2425(.IN1(n750),.IN2(n146),.QN(n751));
  INVX0 U2426(.INP(n1763),.ZN(n1499));
  XOR2X1 U2427(.IN1(n1198),.IN2(n1199),.Q(s_exp_10a[9:9]));
  NAND2X0 U2428(.IN1(s_exp_10_i[8:8]),.IN2(\add_140/carry[8] ),.QN(n1199));
  INVX0 U2429(.INP(s_shr2[4:4]),.ZN(n1282));
  NAND2X0 U2430(.IN1(N2993),.IN2(n1240),.QN(n1573));
  OA21X1 U2431(.IN1(n287),.IN2(n300),.IN3(n301),.Q(n299));
  OA21X1 U2432(.IN1(s_output_o[31:31]),.IN2(n304),.IN3(n305),.Q(n300));
  INVX0 U2433(.INP(n1587),.ZN(n1354));
  AND4X1 U2434(.IN1(n1200),.IN2(n1201),.IN3(n1202),.IN4(n1203),.Q(n306));
  NOR2X0 U2435(.IN1(s_frac2a[0:0]),.IN2(N3244),.QN(n1200));
  INVX0 U2436(.INP(n1576),.ZN(n1381));
  MUX21X1 U2437(.IN1(n1207),.IN2(s_fract_48_i[0:0]),.S(n1260),.Q(n1772));
  INVX0 U2438(.INP(n1760),.ZN(n1514));
  MUX21X1 U2439(.IN1(s_fract_48_i[2:2]),.IN2(n1207),.S(n1260),.Q(n1760));
  INVX0 U2440(.INP(n1756),.ZN(n1506));
  INVX0 U2441(.INP(n1757),.ZN(n1508));
  INVX0 U2442(.INP(n1759),.ZN(n1512));
  MUX21X1 U2443(.IN1(s_fract_48_i[2:2]),.IN2(n1207),.S(n1240),.Q(n1621));
  NAND2X0 U2444(.IN1(s_fract_48_i[0:0]),.IN2(n76),.QN(n1761));
  MUX21X1 U2445(.IN1(n1207),.IN2(s_fract_48_i[0:0]),.S(n1241),.Q(n1516));
  OR4X1 U2446(.IN1(s_shr2[2:2]),.IN2(s_shr2[1:1]),.IN3(s_shr2[0:0]),.IN4(n315),.Q(n1204));
  INVX0 U2447(.INP(s_fract_48_i[13:13]),.ZN(n1496));
  INVX0 U2448(.INP(s_fract_48_i[14:14]),.ZN(n1493));
  INVX0 U2449(.INP(s_fract_48_i[15:15]),.ZN(n1490));
  INVX0 U2450(.INP(s_exp_10a[1:1]),.ZN(n1294));
  INVX0 U2451(.INP(s_fract_48_i[33:33]),.ZN(n1442));
  NBUFFX4 U2452(.INP(s_shl2[4:4]),.Z(n1272));
  INVX0 U2453(.INP(s_fract_48_i[26:26]),.ZN(n1462));
  INVX0 U2454(.INP(s_fract_48_i[28:28]),.ZN(n1460));
  INVX0 U2455(.INP(s_fract_48_i[31:31]),.ZN(n1449));
  INVX0 U2456(.INP(s_fract_48_i[32:32]),.ZN(n1446));
  INVX0 U2457(.INP(s_fract_48_i[16:16]),.ZN(n1487));
  INVX0 U2458(.INP(s_fract_48_i[20:20]),.ZN(n1478));
  INVX0 U2459(.INP(s_fract_48_i[22:22]),.ZN(n1473));
  INVX0 U2460(.INP(s_fract_48_i[17:17]),.ZN(n1485));
  INVX0 U2461(.INP(s_fract_48_i[25:25]),.ZN(n1463));
  INVX0 U2462(.INP(s_fract_48_i[27:27]),.ZN(n1461));
  INVX0 U2463(.INP(s_fract_48_i[29:29]),.ZN(n1458));
  INVX0 U2464(.INP(s_fract_48_i[19:19]),.ZN(n1479));
  INVX0 U2465(.INP(s_fract_48_i[21:21]),.ZN(n1477));
  INVX0 U2466(.INP(s_fract_48_i[23:23]),.ZN(n1468));
  NBUFFX2 U2467(.INP(s_shl2[3:3]),.Z(n1268));
  NBUFFX2 U2468(.INP(s_shr2[5:5]),.Z(n1286));
  NOR2X0 U2469(.IN1(n452),.IN2(s_fract_48_i[4:4]),.QN(n331));
  NAND2X0 U2470(.IN1(n567),.IN2(n231),.QN(n452));
  NBUFFX4 U2471(.INP(s_shl2[4:4]),.Z(n1273));
  NBUFFX2 U2472(.INP(s_shl2[3:3]),.Z(n1269));
  NBUFFX2 U2473(.INP(s_shl2[3:3]),.Z(n1270));
  NAND2X0 U2474(.IN1(n716),.IN2(n47),.QN(n573));
  NOR2X0 U2475(.IN1(n573),.IN2(s_fract_48_i[43:43]),.QN(n661));
  NOR2X0 U2476(.IN1(n573),.IN2(n122),.QN(n718));
  NAND2X1 U2477(.IN1(\s_rmode_i[1] ),.IN2(n236),.QN(n304));
  NBUFFX2 U2478(.INP(s_shl2[3:3]),.Z(n1271));
  NBUFFX2 U2479(.INP(s_shl2[4:4]),.Z(n1274));
  NOR2X0 U2480(.IN1(n1515),.IN2(s_frac_rnd[24:24]),.QN(n248));
  NOR2X0 U2481(.IN1(n244),.IN2(n1515),.QN(n249));
  INVX0 U2482(.INP(s_shr2[4:4]),.ZN(n1281));
  NBUFFX2 U2483(.INP(s_shl2[5:5]),.Z(n1278));
  HADDX2 U2484(.A0(\add_105_I35_L14036_C136/carry[4] ),.B0(N2144),.C1(\add_105_I35_L14036_C136/carry[5] ),.SO(N2154));
  AOI22X1 U2485(.IN1(n909),.IN2(n370),.IN3(N2159),.IN4(n371),.QN(n438));
  HADDX2 U2486(.A0(\add_105_I35_L14036_C136/carry[3] ),.B0(N2143),.C1(\add_105_I35_L14036_C136/carry[4] ),.SO(N2153));
  AOI222X2 U2487(.IN1(n1054),.IN2(n368),.IN3(n1011),.IN4(n1217),.IN5(n817),.IN6(n369),.QN(n439));
  HADDX2 U2488(.A0(\add_105_I33_L14036_C136/carry[3] ),.B0(N2111),.C1(\add_105_I33_L14036_C136/carry[4] ),.SO(N2121));
  HADDX2 U2489(.A0(\add_105_I34_L14036_C136/carry[4] ),.B0(N2128),.C1(\add_105_I34_L14036_C136/carry[5] ),.SO(N2138));
  NAND2X0 U2490(.IN1(n372),.IN2(n742),.QN(n437));
  AOI22X2 U2491(.IN1(n1125),.IN2(n370),.IN3(n1141),.IN4(n371),.QN(n410));
  HADDX2 U2492(.A0(\add_105_I36_L14036_C136/carry[4] ),.B0(N2160),.C1(\add_105_I36_L14036_C136/carry[5] ),.SO(N2170));
  HADDX2 U2493(.A0(\add_105_I33_L14036_C136/carry[4] ),.B0(N2112),.C1(\add_105_I33_L14036_C136/carry[5] ),.SO(N2122));
  INVX0 U2494(.INP(n69),.ZN(n1205));
  INVX0 U2495(.INP(n1206),.ZN(n1207));
  NOR2X0 U2496(.IN1(n1138),.IN2(s_fract_48_i[3:3]),.QN(n1208));
  INVX0 U2497(.INP(N2256),.ZN(n1324));
  INVX0 U2498(.INP(n836),.ZN(n1327));
  INVX0 U2499(.INP(n219),.ZN(n1326));
  HADDX2 U2500(.A0(\add_105_I25_L14036_C136/carry[3] ),.B0(N1983),.C1(\add_105_I25_L14036_C136/carry[4] ),.SO(N1993));
  HADDX2 U2501(.A0(\add_105_I25_L14036_C136/carry[2] ),.B0(N1982),.C1(\add_105_I25_L14036_C136/carry[3] ),.SO(N1992));
  HADDX2 U2502(.A0(\add_105_I27_L14036_C136/carry[3] ),.B0(N2015),.C1(\add_105_I27_L14036_C136/carry[4] ),.SO(N2025));
  HADDX2 U2503(.A0(\add_105_I20_L14036_C136/carry[3] ),.B0(N1903),.C1(\add_105_I20_L14036_C136/carry[4] ),.SO(N1913));
  HADDX2 U2504(.A0(\add_105_I34_L14036_C136/carry[3] ),.B0(n17),.C1(\add_105_I34_L14036_C136/carry[4] ),.SO(N2137));
  HADDX2 U2505(.A0(\add_105_I24_L14036_C136/carry[3] ),.B0(N1967),.C1(\add_105_I24_L14036_C136/carry[4] ),.SO(N1977));
  HADDX2 U2506(.A0(\add_105_I24_L14036_C136/carry[2] ),.B0(N1966),.C1(\add_105_I24_L14036_C136/carry[3] ),.SO(N1976));
  HADDX2 U2507(.A0(\add_105_I23_L14036_C136/carry[4] ),.B0(N1952),.C1(\add_105_I23_L14036_C136/carry[5] ),.SO(N1962));
  INVX0 U2508(.INP(n195),.ZN(n1328));
  HADDX2 U2509(.A0(\add_105_I31_L14036_C136/carry[4] ),.B0(N2080),.C1(\add_105_I31_L14036_C136/carry[5] ),.SO(N2090));
  INVX0 U2510(.INP(n837),.ZN(n1469));
  INVX0 U2511(.INP(n828),.ZN(n1402));
  INVX0 U2512(.INP(n240),.ZN(n1502));
  NAND2X1 U2513(.IN1(n1466),.IN2(n683),.QN(n463));
  INVX0 U2514(.INP(n132),.ZN(n1455));
  INVX0 U2515(.INP(n917),.ZN(n1403));
  NOR2X0 U2516(.IN1(s_fract_48_i[45:45]),.IN2(s_fract_48_i[46:46]),.QN(n800));
  NOR2X0 U2517(.IN1(n803),.IN2(s_fract_48_i[43:43]),.QN(n801));
  OA21X1 U2518(.IN1(n391),.IN2(n392),.IN3(n331),.Q(N2978));
  NAND2X0 U2519(.IN1(n1451),.IN2(n899),.QN(n727));
  NAND2X0 U2520(.IN1(n612),.IN2(n1088),.QN(n650));
  AO22X2 U2521(.IN1(n346),.IN2(n941),.IN3(n345),.IN4(n954),.Q(n490));
  NAND2X0 U2522(.IN1(n1466),.IN2(n947),.QN(n492));
  NAND2X0 U2523(.IN1(n372),.IN2(n1131),.QN(n409));
  NOR2X0 U2524(.IN1(n571),.IN2(s_fract_48_i[3:3]),.QN(n569));
  NOR2X0 U2525(.IN1(s_fract_48_i[0:0]),.IN2(n1135),.QN(n481));
  NBUFFX2 U2526(.INP(s_fract_48_i[5:5]),.Z(n1220));
  NBUFFX2 U2527(.INP(s_fract_48_i[5:5]),.Z(n1221));
  NBUFFX2 U2528(.INP(s_fract_48_i[5:5]),.Z(n1222));
  NBUFFX2 U2529(.INP(s_fract_48_i[5:5]),.Z(n1223));
  NBUFFX2 U2530(.INP(s_fract_48_i[6:6]),.Z(n1224));
  NBUFFX2 U2531(.INP(s_fract_48_i[6:6]),.Z(n1225));
  NBUFFX2 U2532(.INP(s_fract_48_i[6:6]),.Z(n1226));
  NBUFFX2 U2533(.INP(s_fract_48_i[6:6]),.Z(n1227));
  NBUFFX2 U2534(.INP(s_fract_48_i[42:42]),.Z(n1229));
  NBUFFX2 U2535(.INP(s_fract_48_i[42:42]),.Z(n1230));
  INVX0 U2536(.INP(n1247),.ZN(n1243));
  INVX0 U2537(.INP(n1247),.ZN(n1244));
  INVX0 U2538(.INP(n1247),.ZN(n1245));
  INVX0 U2539(.INP(n1247),.ZN(n1246));
  INVX0 U2540(.INP(n1257),.ZN(n1255));
  INVX0 U2541(.INP(n1257),.ZN(n1256));
  INVX0 U2542(.INP(n76),.ZN(n1260));
  INVX0 U2543(.INP(n76),.ZN(n1261));
  INVX0 U2544(.INP(n76),.ZN(n1262));
  INVX0 U2545(.INP(n53),.ZN(n1263));
  INVX0 U2546(.INP(n53),.ZN(n1264));
  INVX0 U2547(.INP(n53),.ZN(n1265));
  INVX0 U2548(.INP(n56),.ZN(n1266));
  INVX0 U2549(.INP(n56),.ZN(n1267));
  INVX0 U2550(.INP(n1282),.ZN(n1279));
  INVX0 U2551(.INP(n1282),.ZN(n1280));
  INVX0 U2552(.INP(s_fract_48_i[12:12]),.ZN(n1287));
  INVX0 U2553(.INP(s_fract_48_i[18:18]),.ZN(n1288));
  INVX0 U2554(.INP(n1291),.ZN(n1289));
  INVX0 U2555(.INP(n1291),.ZN(n1290));
  INVX0 U2556(.INP(s_fract_48_i[30:30]),.ZN(n1292));
  XNOR2X1 U2557(.IN1(\sub_192_aco/carry[7] ),.IN2(s_expo1[7:7]),.Q(s_expo2b[7:7]));
  OR2X1 U2558(.IN1(s_expo1[6:6]),.IN2(\sub_192_aco/carry[6] ),.Q(\sub_192_aco/carry[7] ));
  XNOR2X1 U2559(.IN1(\sub_192_aco/carry[6] ),.IN2(s_expo1[6:6]),.Q(s_expo2b[6:6]));
  OR2X1 U2560(.IN1(s_expo1[5:5]),.IN2(\sub_192_aco/carry[5] ),.Q(\sub_192_aco/carry[6] ));
  XNOR2X1 U2561(.IN1(\sub_192_aco/carry[5] ),.IN2(s_expo1[5:5]),.Q(s_expo2b[5:5]));
  OR2X1 U2562(.IN1(s_expo1[4:4]),.IN2(\sub_192_aco/carry[4] ),.Q(\sub_192_aco/carry[5] ));
  XNOR2X1 U2563(.IN1(\sub_192_aco/carry[4] ),.IN2(s_expo1[4:4]),.Q(s_expo2b[4:4]));
  OR2X1 U2564(.IN1(s_expo1[3:3]),.IN2(\sub_192_aco/carry[3] ),.Q(\sub_192_aco/carry[4] ));
  XNOR2X1 U2565(.IN1(\sub_192_aco/carry[3] ),.IN2(s_expo1[3:3]),.Q(s_expo2b[3:3]));
  OR2X1 U2566(.IN1(s_expo1[2:2]),.IN2(\sub_192_aco/carry[2] ),.Q(\sub_192_aco/carry[3] ));
  XNOR2X1 U2567(.IN1(\sub_192_aco/carry[2] ),.IN2(s_expo1[2:2]),.Q(s_expo2b[2:2]));
  OR2X1 U2568(.IN1(s_expo1[1:1]),.IN2(\sub_192_aco/carry[1] ),.Q(\sub_192_aco/carry[2] ));
  XNOR2X1 U2569(.IN1(\sub_192_aco/carry[1] ),.IN2(s_expo1[1:1]),.Q(s_expo2b[1:1]));
  OR2X1 U2570(.IN1(s_expo1[0:0]),.IN2(s_frac2a[46:46]),.Q(\sub_192_aco/carry[1] ));
  XNOR2X1 U2571(.IN1(s_frac2a[46:46]),.IN2(s_expo1[0:0]),.Q(s_expo2b[0:0]));
  XOR2X1 U2572(.IN1(n1280),.IN2(\add_197/carry[4] ),.Q(N3242));
  AND2X1 U2573(.IN1(\add_197/carry[3] ),.IN2(s_shr2[3:3]),.Q(\add_197/carry[4] ));
  XOR2X1 U2574(.IN1(s_shr2[3:3]),.IN2(\add_197/carry[3] ),.Q(N3241));
  AND2X1 U2575(.IN1(\add_197/carry[2] ),.IN2(s_shr2[2:2]),.Q(\add_197/carry[3] ));
  XOR2X1 U2576(.IN1(s_shr2[2:2]),.IN2(\add_197/carry[2] ),.Q(N3240));
  AND2X1 U2577(.IN1(\add_197/carry[1] ),.IN2(s_shr2[1:1]),.Q(\add_197/carry[2] ));
  XOR2X1 U2578(.IN1(s_shr2[1:1]),.IN2(\add_197/carry[1] ),.Q(N3239));
  AND2X1 U2579(.IN1(s_frac_rnd[24:24]),.IN2(s_shr2[0:0]),.Q(\add_197/carry[1] ));
  XOR2X1 U2580(.IN1(s_shr2[0:0]),.IN2(s_frac_rnd[24:24]),.Q(N3238));
  XOR2X1 U2581(.IN1(n1298),.IN2(\sub_0_root_add_0_root_add_148/carry[5] ),.Q(N3004));
  AND2X1 U2582(.IN1(\sub_0_root_add_0_root_add_148/carry[4] ),.IN2(n1297),.Q(\sub_0_root_add_0_root_add_148/carry[5] ));
  XOR2X1 U2583(.IN1(n1297),.IN2(\sub_0_root_add_0_root_add_148/carry[4] ),.Q(N3003));
  AND2X1 U2584(.IN1(\sub_0_root_add_0_root_add_148/carry[3] ),.IN2(n1296),.Q(\sub_0_root_add_0_root_add_148/carry[4] ));
  XOR2X1 U2585(.IN1(n1296),.IN2(\sub_0_root_add_0_root_add_148/carry[3] ),.Q(N3002));
  AND2X1 U2586(.IN1(\sub_0_root_add_0_root_add_148/carry[2] ),.IN2(n1295),.Q(\sub_0_root_add_0_root_add_148/carry[3] ));
  XOR2X1 U2587(.IN1(n1295),.IN2(\sub_0_root_add_0_root_add_148/carry[2] ),.Q(N3001));
  OR2X1 U2588(.IN1(n68),.IN2(n1293),.Q(\sub_0_root_add_0_root_add_148/carry[1] ));
  XNOR2X1 U2589(.IN1(n1293),.IN2(n68),.Q(N2999));
  XOR2X1 U2590(.IN1(s_exp_10_i[8:8]),.IN2(\add_140/carry[8] ),.Q(s_exp_10a[8:8]));
  AND2X1 U2591(.IN1(s_exp_10_i[7:7]),.IN2(\add_140/carry[7] ),.Q(\add_140/carry[8] ));
  XOR2X1 U2592(.IN1(s_exp_10_i[7:7]),.IN2(\add_140/carry[7] ),.Q(s_exp_10a[7:7]));
  AND2X1 U2593(.IN1(s_exp_10_i[6:6]),.IN2(\add_140/carry[6] ),.Q(\add_140/carry[7] ));
  XOR2X1 U2594(.IN1(s_exp_10_i[6:6]),.IN2(\add_140/carry[6] ),.Q(s_exp_10a[6:6]));
  AND2X1 U2595(.IN1(s_exp_10_i[5:5]),.IN2(\add_140/carry[5] ),.Q(\add_140/carry[6] ));
  XOR2X1 U2596(.IN1(s_exp_10_i[5:5]),.IN2(\add_140/carry[5] ),.Q(s_exp_10a[5:5]));
  AND2X1 U2597(.IN1(s_exp_10_i[4:4]),.IN2(\add_140/carry[4] ),.Q(\add_140/carry[5] ));
  XOR2X1 U2598(.IN1(s_exp_10_i[4:4]),.IN2(\add_140/carry[4] ),.Q(s_exp_10a[4:4]));
  AND2X1 U2599(.IN1(s_exp_10_i[3:3]),.IN2(\add_140/carry[3] ),.Q(\add_140/carry[4] ));
  XOR2X1 U2600(.IN1(s_exp_10_i[3:3]),.IN2(\add_140/carry[3] ),.Q(s_exp_10a[3:3]));
  AND2X1 U2601(.IN1(s_exp_10_i[2:2]),.IN2(\add_140/carry[2] ),.Q(\add_140/carry[3] ));
  XOR2X1 U2602(.IN1(s_exp_10_i[2:2]),.IN2(\add_140/carry[2] ),.Q(s_exp_10a[2:2]));
  AND2X1 U2603(.IN1(s_exp_10_i[1:1]),.IN2(\add_140/carry[1] ),.Q(\add_140/carry[2] ));
  XOR2X1 U2604(.IN1(s_exp_10_i[1:1]),.IN2(\add_140/carry[1] ),.Q(s_exp_10a[1:1]));
  AND2X1 U2605(.IN1(s_exp_10_i[0:0]),.IN2(N2993),.Q(\add_140/carry[1] ));
  XOR2X1 U2606(.IN1(s_exp_10_i[0:0]),.IN2(N2993),.Q(s_exp_10a[0:0]));
  XOR2X1 U2607(.IN1(\add_90_I9_L14036_C132/carry[5] ),.IN2(N401),.Q(N412));
  XOR2X1 U2608(.IN1(\add_90_I12_L14036_C132/carry[5] ),.IN2(N452),.Q(N463));
  XOR2X1 U2609(.IN1(\add_90_I13_L14036_C132/carry[5] ),.IN2(N469),.Q(N480));
  XOR2X1 U2610(.IN1(\add_90_I14_L14036_C132/carry[5] ),.IN2(N486),.Q(N497));
  XOR2X1 U2611(.IN1(\add_90_I16_L14036_C132/carry[5] ),.IN2(N520),.Q(N531));
  XOR2X1 U2612(.IN1(\add_90_I17_L14036_C132/carry[5] ),.IN2(N537),.Q(N548));
  XOR2X1 U2613(.IN1(\add_90_I19_L14036_C132/carry[5] ),.IN2(N571),.Q(N582));
  XOR2X1 U2614(.IN1(\add_90_I21_L14036_C132/carry[5] ),.IN2(n1015),.Q(N616));
  XOR2X1 U2615(.IN1(\add_90_I22_L14036_C132/carry[5] ),.IN2(N622),.Q(N633));
  XOR2X1 U2616(.IN1(\add_90_I25_L14036_C132/carry[5] ),.IN2(n979),.Q(N684));
  XOR2X1 U2617(.IN1(\add_90_I26_L14036_C132/carry[5] ),.IN2(N690),.Q(N701));
  XOR2X1 U2618(.IN1(\add_90_I27_L14036_C132/carry[5] ),.IN2(N707),.Q(N718));
  XOR2X1 U2619(.IN1(\add_90_I28_L14036_C132/carry[5] ),.IN2(n855),.Q(N735));
  XOR2X1 U2620(.IN1(\add_90_I31_L14036_C132/carry[5] ),.IN2(N775),.Q(N786));
  XOR2X1 U2621(.IN1(\add_105_I11_L14036_C136/carry[5] ),.IN2(N1761),.Q(N1771));
  XOR2X1 U2622(.IN1(\add_105_I15_L14036_C136/carry[5] ),.IN2(N1825),.Q(N1835));
  XOR2X1 U2623(.IN1(\add_105_I17_L14036_C136/carry[5] ),.IN2(N1857),.Q(N1867));
  XOR2X1 U2624(.IN1(\add_105_I18_L14036_C136/carry[5] ),.IN2(n897),.Q(N1883));
  XOR2X1 U2625(.IN1(\add_105_I22_L14036_C136/carry[5] ),.IN2(n975),.Q(N1947));
  XOR2X1 U2626(.IN1(\add_105_I24_L14036_C136/carry[5] ),.IN2(N1969),.Q(N1979));
  XOR2X1 U2627(.IN1(\add_105_I25_L14036_C136/carry[5] ),.IN2(n905),.Q(N1995));
  XOR2X1 U2628(.IN1(\add_105_I28_L14036_C136/carry[5] ),.IN2(n1038),.Q(N2043));
  XOR2X1 U2629(.IN1(\add_105_I35_L14036_C136/carry[5] ),.IN2(N2145),.Q(N2155));
  XOR2X1 U2630(.IN1(\add_105_I38_L14036_C136/carry[5] ),.IN2(N2193),.Q(N2203));
  AO22X1 U2631(.IN1(N3243),.IN2(n54),.IN3(N3242),.IN4(n78),.Q(n1309));
  OR2X1 U2632(.IN1(n54),.IN2(N3243),.Q(n1308));
  NOR2X0 U2633(.IN1(n74),.IN2(N3241),.QN(n1299));
  AOI21X1 U2634(.IN1(n1310),.IN2(s_r_zeros[2:2]),.IN3(n1299),.QN(n1305));
  NOR2X0 U2635(.IN1(s_r_zeros[2:2]),.IN2(n1299),.QN(n1300));
  AO22X1 U2636(.IN1(N3241),.IN2(n74),.IN3(n1300),.IN4(N3240),.Q(n1304));
  NOR2X0 U2637(.IN1(N3239),.IN2(n75),.QN(n1301));
  NOR2X0 U2638(.IN1(s_r_zeros[0:0]),.IN2(n1301),.QN(n1302));
  AO221X1 U2639(.IN1(N3239),.IN2(n75),.IN3(n1302),.IN4(N3238),.IN5(n1304),.Q(n1303));
  OA21X1 U2640(.IN1(n1305),.IN2(n1304),.IN3(n1303),.Q(n1307));
  OA21X1 U2641(.IN1(N3242),.IN2(n78),.IN3(n1308),.Q(n1306));
  AO22X1 U2642(.IN1(n1309),.IN2(n1308),.IN3(n1307),.IN4(n1306),.Q(N3244));
  AND2X1 U2643(.IN1(N1690),.IN2(n227),.Q(N1696));
  AND2X1 U2644(.IN1(N360),.IN2(n130),.Q(N366));
  MUX21X1 U2645(.IN1(s_fract_48_i[31:31]),.IN2(n1217),.S(n1242),.Q(n1527));
  MUX21X1 U2646(.IN1(s_fract_48_i[29:29]),.IN2(s_fract_48_i[28:28]),.S(n1242),.Q(n1526));
  MUX21X1 U2647(.IN1(n1527),.IN2(n1526),.S(n1239),.Q(n1546));
  MUX21X1 U2648(.IN1(s_fract_48_i[27:27]),.IN2(s_fract_48_i[26:26]),.S(n1242),.Q(n1525));
  MUX21X1 U2649(.IN1(s_fract_48_i[25:25]),.IN2(n1289),.S(n1242),.Q(n1532));
  MUX21X1 U2650(.IN1(n1525),.IN2(n1532),.S(n1239),.Q(n1549));
  MUX21X1 U2651(.IN1(n1546),.IN2(n1549),.S(n1236),.Q(n1650));
  MUX21X1 U2652(.IN1(s_fract_48_i[23:23]),.IN2(s_fract_48_i[22:22]),.S(n1242),.Q(n1531));
  MUX21X1 U2653(.IN1(s_fract_48_i[21:21]),.IN2(s_fract_48_i[20:20]),.S(n1242),.Q(n1530));
  MUX21X1 U2654(.IN1(n1531),.IN2(n1530),.S(n1239),.Q(n1548));
  MUX21X1 U2655(.IN1(s_fract_48_i[19:19]),.IN2(n1214),.S(n1242),.Q(n1529));
  MUX21X1 U2656(.IN1(s_fract_48_i[17:17]),.IN2(s_fract_48_i[16:16]),.S(n1242),.Q(n1536));
  MUX21X1 U2657(.IN1(n1529),.IN2(n1536),.S(n1239),.Q(n1551));
  MUX21X1 U2658(.IN1(n1548),.IN2(n1551),.S(n1236),.Q(n1744));
  MUX21X1 U2659(.IN1(n1650),.IN2(n1744),.S(n1234),.Q(n1597));
  MUX21X1 U2660(.IN1(s_fract_48_i[15:15]),.IN2(s_fract_48_i[14:14]),.S(n1242),.Q(n1535));
  MUX21X1 U2661(.IN1(s_fract_48_i[13:13]),.IN2(n1210),.S(n1242),.Q(n1534));
  MUX21X1 U2662(.IN1(n1535),.IN2(n1534),.S(n1239),.Q(n1550));
  MUX21X1 U2663(.IN1(s_fract_48_i[11:11]),.IN2(s_fract_48_i[10:10]),.S(n1242),.Q(n1533));
  MUX21X1 U2664(.IN1(s_fract_48_i[9:9]),.IN2(s_fract_48_i[8:8]),.S(n1241),.Q(n1671));
  MUX21X1 U2665(.IN1(n1533),.IN2(n1671),.S(n1239),.Q(n1713));
  MUX21X1 U2666(.IN1(n1550),.IN2(n1713),.S(n1236),.Q(n1745));
  MUX21X1 U2667(.IN1(s_fract_48_i[2:2]),.IN2(s_fract_48_i[3:3]),.S(s_shr2[0:0]),.Q(n1668));
  MUX21X1 U2668(.IN1(n1668),.IN2(n1516),.S(n1239),.Q(n1517));
  MUX21X1 U2669(.IN1(s_fract_48_i[7:7]),.IN2(n1227),.S(n1241),.Q(n1670));
  MUX21X1 U2670(.IN1(n1221),.IN2(s_fract_48_i[4:4]),.S(n1241),.Q(n1669));
  MUX21X1 U2671(.IN1(n1670),.IN2(n1669),.S(n1239),.Q(n1712));
  MUX21X1 U2672(.IN1(n1517),.IN2(n1712),.S(s_shr2[2:2]),.Q(n1518));
  MUX21X1 U2673(.IN1(n1745),.IN2(n1518),.S(n1234),.Q(n1519));
  MUX21X1 U2674(.IN1(n1597),.IN2(n1519),.S(n1281),.Q(n1520));
  MUX21X1 U2675(.IN1(N2993),.IN2(n1205),.S(n1241),.Q(n1540));
  MUX21X1 U2676(.IN1(s_fract_48_i[45:45]),.IN2(s_fract_48_i[44:44]),.S(n1241),.Q(n1539));
  MUX21X1 U2677(.IN1(n1540),.IN2(n1539),.S(n1239),.Q(n1553));
  MUX21X1 U2678(.IN1(s_fract_48_i[43:43]),.IN2(n1231),.S(n1241),.Q(n1538));
  MUX21X1 U2679(.IN1(s_fract_48_i[41:41]),.IN2(s_fract_48_i[40:40]),.S(n1241),.Q(n1524));
  MUX21X1 U2680(.IN1(n1538),.IN2(n1524),.S(n1239),.Q(n1545));
  MUX21X1 U2681(.IN1(n1553),.IN2(n1545),.S(n1236),.Q(n1648));
  MUX21X1 U2682(.IN1(s_fract_48_i[39:39]),.IN2(s_fract_48_i[38:38]),.S(n1241),.Q(n1523));
  MUX21X1 U2683(.IN1(s_fract_48_i[37:37]),.IN2(s_fract_48_i[36:36]),.S(n1241),.Q(n1522));
  MUX21X1 U2684(.IN1(n1523),.IN2(n1522),.S(n1239),.Q(n1544));
  MUX21X1 U2685(.IN1(s_fract_48_i[35:35]),.IN2(s_fract_48_i[34:34]),.S(n1241),.Q(n1521));
  MUX21X1 U2686(.IN1(s_fract_48_i[33:33]),.IN2(s_fract_48_i[32:32]),.S(n1241),.Q(n1528));
  MUX21X1 U2687(.IN1(n1521),.IN2(n1528),.S(n1239),.Q(n1547));
  MUX21X1 U2688(.IN1(n1544),.IN2(n1547),.S(n1236),.Q(n1649));
  MUX21X1 U2689(.IN1(n1648),.IN2(n1649),.S(n1233),.Q(n1598));
  MUX21X1 U2690(.IN1(n1520),.IN2(n1337),.S(n1285),.Q(N3093));
  MUX21X1 U2691(.IN1(n1522),.IN2(n1521),.S(n1238),.Q(n1578));
  MUX21X1 U2692(.IN1(n1524),.IN2(n1523),.S(n1238),.Q(n1575));
  MUX21X1 U2693(.IN1(n1578),.IN2(n1575),.S(s_shr2[2:2]),.Q(n1609));
  MUX21X1 U2694(.IN1(n1526),.IN2(n1525),.S(n1238),.Q(n1580));
  MUX21X1 U2695(.IN1(n1528),.IN2(n1527),.S(n1238),.Q(n1577));
  MUX21X1 U2696(.IN1(n1580),.IN2(n1577),.S(s_shr2[2:2]),.Q(n1612));
  MUX21X1 U2697(.IN1(n1609),.IN2(n1612),.S(n1233),.Q(n1656));
  MUX21X1 U2698(.IN1(n1530),.IN2(n1529),.S(n1238),.Q(n1582));
  MUX21X1 U2699(.IN1(n1532),.IN2(n1531),.S(n1238),.Q(n1579));
  MUX21X1 U2700(.IN1(n1582),.IN2(n1579),.S(s_shr2[2:2]),.Q(n1611));
  MUX21X1 U2701(.IN1(n1534),.IN2(n1533),.S(n1238),.Q(n1729));
  MUX21X1 U2702(.IN1(n1536),.IN2(n1535),.S(n1238),.Q(n1581));
  MUX21X1 U2703(.IN1(n1729),.IN2(n1581),.S(s_shr2[2:2]),.Q(n1674));
  MUX21X1 U2704(.IN1(n1611),.IN2(n1674),.S(n1233),.Q(n1537));
  MUX21X1 U2705(.IN1(n1656),.IN2(n1537),.S(n79),.Q(n1541));
  MUX21X1 U2706(.IN1(n1539),.IN2(n1538),.S(n1238),.Q(n1576));
  MUX21X1 U2707(.IN1(n1381),.IN2(n1584),.S(s_shr2[2:2]),.Q(n1610));
  OR2X1 U2708(.IN1(n1610),.IN2(s_shr2[3:3]),.Q(n1657));
  MUX21X1 U2709(.IN1(n1541),.IN2(n1706),.S(n1286),.Q(N3103));
  MUX21X1 U2710(.IN1(s_fract_48_i[38:38]),.IN2(s_fract_48_i[37:37]),.S(n1241),.Q(n1557));
  MUX21X1 U2711(.IN1(s_fract_48_i[36:36]),.IN2(s_fract_48_i[35:35]),.S(n1241),.Q(n1560));
  MUX21X1 U2712(.IN1(n1557),.IN2(n1560),.S(n1238),.Q(n1589));
  MUX21X1 U2713(.IN1(n1230),.IN2(s_fract_48_i[41:41]),.S(n1241),.Q(n1555));
  MUX21X1 U2714(.IN1(s_fract_48_i[40:40]),.IN2(s_fract_48_i[39:39]),.S(n1241),.Q(n1558));
  MUX21X1 U2715(.IN1(n1555),.IN2(n1558),.S(n1238),.Q(n1586));
  MUX21X1 U2716(.IN1(n1589),.IN2(n1586),.S(s_shr2[2:2]),.Q(n1614));
  MUX21X1 U2717(.IN1(n1216),.IN2(s_fract_48_i[29:29]),.S(n1241),.Q(n1561));
  MUX21X1 U2718(.IN1(s_fract_48_i[28:28]),.IN2(s_fract_48_i[27:27]),.S(n1241),.Q(n1564));
  MUX21X1 U2719(.IN1(n1561),.IN2(n1564),.S(n1238),.Q(n1591));
  MUX21X1 U2720(.IN1(s_fract_48_i[34:34]),.IN2(s_fract_48_i[33:33]),.S(n1240),.Q(n1559));
  MUX21X1 U2721(.IN1(s_fract_48_i[32:32]),.IN2(s_fract_48_i[31:31]),.S(n1240),.Q(n1562));
  MUX21X1 U2722(.IN1(n1559),.IN2(n1562),.S(n1238),.Q(n1588));
  MUX21X1 U2723(.IN1(n1591),.IN2(n1588),.S(s_shr2[2:2]),.Q(n1617));
  MUX21X1 U2724(.IN1(n1614),.IN2(n1617),.S(n1233),.Q(n1659));
  MUX21X1 U2725(.IN1(s_fract_48_i[22:22]),.IN2(s_fract_48_i[21:21]),.S(n1240),.Q(n1565));
  MUX21X1 U2726(.IN1(s_fract_48_i[20:20]),.IN2(s_fract_48_i[19:19]),.S(n1240),.Q(n1568));
  MUX21X1 U2727(.IN1(n1565),.IN2(n1568),.S(n1238),.Q(n1593));
  MUX21X1 U2728(.IN1(s_fract_48_i[26:26]),.IN2(s_fract_48_i[25:25]),.S(n1240),.Q(n1563));
  MUX21X1 U2729(.IN1(n1289),.IN2(s_fract_48_i[23:23]),.S(n1240),.Q(n1566));
  MUX21X1 U2730(.IN1(n1563),.IN2(n1566),.S(n1238),.Q(n1590));
  MUX21X1 U2731(.IN1(n1593),.IN2(n1590),.S(s_shr2[2:2]),.Q(n1616));
  MUX21X1 U2732(.IN1(s_fract_48_i[14:14]),.IN2(s_fract_48_i[13:13]),.S(n1240),.Q(n1569));
  MUX21X1 U2733(.IN1(n1211),.IN2(s_fract_48_i[11:11]),.S(n1240),.Q(n1619));
  MUX21X1 U2734(.IN1(n1569),.IN2(n1619),.S(n1238),.Q(n1737));
  MUX21X1 U2735(.IN1(n1213),.IN2(s_fract_48_i[17:17]),.S(n1240),.Q(n1567));
  MUX21X1 U2736(.IN1(s_fract_48_i[16:16]),.IN2(s_fract_48_i[15:15]),.S(n1240),.Q(n1570));
  MUX21X1 U2737(.IN1(n1567),.IN2(n1570),.S(n1238),.Q(n1592));
  MUX21X1 U2738(.IN1(n1737),.IN2(n1592),.S(s_shr2[2:2]),.Q(n1699));
  MUX21X1 U2739(.IN1(n1616),.IN2(n1699),.S(n1233),.Q(n1542));
  MUX21X1 U2740(.IN1(n1659),.IN2(n1542),.S(n79),.Q(n1543));
  MUX21X1 U2741(.IN1(n1205),.IN2(s_fract_48_i[45:45]),.S(n1240),.Q(n1572));
  MUX21X1 U2742(.IN1(s_fract_48_i[44:44]),.IN2(s_fract_48_i[43:43]),.S(n1240),.Q(n1556));
  MUX21X1 U2743(.IN1(n1572),.IN2(n1556),.S(n1238),.Q(n1587));
  OR2X1 U2744(.IN1(n1573),.IN2(s_shr2[1:1]),.Q(n1595));
  MUX21X1 U2745(.IN1(n1354),.IN2(n1595),.S(s_shr2[2:2]),.Q(n1615));
  OR2X1 U2746(.IN1(n1615),.IN2(s_shr2[3:3]),.Q(n1660));
  MUX21X1 U2747(.IN1(n1543),.IN2(n1707),.S(n1285),.Q(N3104));
  MUX21X1 U2748(.IN1(n1545),.IN2(n1544),.S(n1236),.Q(n1628));
  MUX21X1 U2749(.IN1(n1547),.IN2(n1546),.S(n1236),.Q(n1631));
  MUX21X1 U2750(.IN1(n1628),.IN2(n1631),.S(n1233),.Q(n1662));
  MUX21X1 U2751(.IN1(n1549),.IN2(n1548),.S(n1236),.Q(n1630));
  MUX21X1 U2752(.IN1(n1551),.IN2(n1550),.S(n1236),.Q(n1715));
  MUX21X1 U2753(.IN1(n1630),.IN2(n1715),.S(n1233),.Q(n1552));
  MUX21X1 U2754(.IN1(n1662),.IN2(n1552),.S(n79),.Q(n1554));
  OR2X1 U2755(.IN1(n1629),.IN2(s_shr2[3:3]),.Q(n1663));
  MUX21X1 U2756(.IN1(n1554),.IN2(n1708),.S(n1285),.Q(N3105));
  MUX21X1 U2757(.IN1(n1556),.IN2(n1555),.S(n1237),.Q(n1600));
  MUX21X1 U2758(.IN1(n1558),.IN2(n1557),.S(n1237),.Q(n1603));
  MUX21X1 U2759(.IN1(n1600),.IN2(n1603),.S(n1236),.Q(n1633));
  MUX21X1 U2760(.IN1(n1560),.IN2(n1559),.S(n1237),.Q(n1602));
  MUX21X1 U2761(.IN1(n1562),.IN2(n1561),.S(n1237),.Q(n1605));
  MUX21X1 U2762(.IN1(n1602),.IN2(n1605),.S(n1236),.Q(n1636));
  MUX21X1 U2763(.IN1(n1633),.IN2(n1636),.S(n1233),.Q(n1665));
  MUX21X1 U2764(.IN1(n1564),.IN2(n1563),.S(n1237),.Q(n1604));
  MUX21X1 U2765(.IN1(n1566),.IN2(n1565),.S(n1237),.Q(n1607));
  MUX21X1 U2766(.IN1(n1604),.IN2(n1607),.S(n1236),.Q(n1635));
  MUX21X1 U2767(.IN1(n1568),.IN2(n1567),.S(n1237),.Q(n1606));
  MUX21X1 U2768(.IN1(n1570),.IN2(n1569),.S(n1237),.Q(n1620));
  MUX21X1 U2769(.IN1(n1606),.IN2(n1620),.S(n1236),.Q(n1723));
  MUX21X1 U2770(.IN1(n1635),.IN2(n1723),.S(n1233),.Q(n1571));
  MUX21X1 U2771(.IN1(n1665),.IN2(n1571),.S(n1281),.Q(n1574));
  MUX21X1 U2772(.IN1(n1573),.IN2(n1357),.S(n1237),.Q(n1601));
  OR2X1 U2773(.IN1(n1601),.IN2(s_shr2[2:2]),.Q(n1634));
  OR2X1 U2774(.IN1(n1634),.IN2(s_shr2[3:3]),.Q(n1666));
  MUX21X1 U2775(.IN1(n1574),.IN2(n1709),.S(n1285),.Q(N3106));
  MUX21X1 U2776(.IN1(n1576),.IN2(n1575),.S(n1236),.Q(n1638));
  MUX21X1 U2777(.IN1(n1578),.IN2(n1577),.S(n1235),.Q(n1641));
  MUX21X1 U2778(.IN1(n1638),.IN2(n1641),.S(n1233),.Q(n1679));
  MUX21X1 U2779(.IN1(n1580),.IN2(n1579),.S(n1235),.Q(n1640));
  MUX21X1 U2780(.IN1(n1582),.IN2(n1581),.S(n1235),.Q(n1731));
  MUX21X1 U2781(.IN1(n1640),.IN2(n1731),.S(n1233),.Q(n1583));
  MUX21X1 U2782(.IN1(n1679),.IN2(n1583),.S(n79),.Q(n1585));
  OR2X1 U2783(.IN1(n1584),.IN2(s_shr2[2:2]),.Q(n1639));
  OR2X1 U2784(.IN1(n1639),.IN2(s_shr2[3:3]),.Q(n1680));
  MUX21X1 U2785(.IN1(n1585),.IN2(n1710),.S(n1286),.Q(N3107));
  MUX21X1 U2786(.IN1(n1587),.IN2(n1586),.S(n1235),.Q(n1643));
  MUX21X1 U2787(.IN1(n1589),.IN2(n1588),.S(n1235),.Q(n1646));
  MUX21X1 U2788(.IN1(n1643),.IN2(n1646),.S(n1233),.Q(n1682));
  MUX21X1 U2789(.IN1(n1591),.IN2(n1590),.S(n1235),.Q(n1645));
  MUX21X1 U2790(.IN1(n1593),.IN2(n1592),.S(n1235),.Q(n1739));
  MUX21X1 U2791(.IN1(n1645),.IN2(n1739),.S(n1233),.Q(n1594));
  MUX21X1 U2792(.IN1(n1682),.IN2(n1594),.S(n1281),.Q(n1596));
  OR2X1 U2793(.IN1(n1595),.IN2(s_shr2[2:2]),.Q(n1644));
  OR2X1 U2794(.IN1(n1644),.IN2(s_shr2[3:3]),.Q(n1683));
  MUX21X1 U2795(.IN1(n1596),.IN2(n1711),.S(n1285),.Q(N3108));
  MUX21X1 U2796(.IN1(n1598),.IN2(n1597),.S(n79),.Q(n1599));
  MUX21X1 U2797(.IN1(n1601),.IN2(n1386),.S(n1235),.Q(n1652));
  MUX21X1 U2798(.IN1(n1603),.IN2(n1602),.S(n1235),.Q(n1653));
  MUX21X1 U2799(.IN1(n1652),.IN2(n1405),.S(n1233),.Q(n1626));
  MUX21X1 U2800(.IN1(n1605),.IN2(n1604),.S(n1235),.Q(n1654));
  MUX21X1 U2801(.IN1(n1607),.IN2(n1606),.S(n1235),.Q(n1750));
  MUX21X1 U2802(.IN1(n1654),.IN2(n1750),.S(n1233),.Q(n1625));
  MUX21X1 U2803(.IN1(n1626),.IN2(n1444),.S(n79),.Q(n1608));
  MUX21X1 U2804(.IN1(n1610),.IN2(n1399),.S(n1233),.Q(n1677));
  MUX21X1 U2805(.IN1(n1612),.IN2(n1611),.S(n1233),.Q(n1676));
  MUX21X1 U2806(.IN1(n1677),.IN2(n1440),.S(n1281),.Q(n1613));
  MUX21X1 U2807(.IN1(n1615),.IN2(n1394),.S(n1233),.Q(n1688));
  MUX21X1 U2808(.IN1(n1617),.IN2(n1616),.S(n1232),.Q(n1700));
  MUX21X1 U2809(.IN1(n1688),.IN2(n1436),.S(n1281),.Q(n1618));
  MUX21X1 U2810(.IN1(s_fract_48_i[10:10]),.IN2(s_fract_48_i[9:9]),.S(n1240),.Q(n1696));
  MUX21X1 U2811(.IN1(n1619),.IN2(n1696),.S(n1237),.Q(n1721));
  MUX21X1 U2812(.IN1(n1620),.IN2(n1721),.S(n1235),.Q(n1751));
  MUX21X1 U2813(.IN1(s_fract_48_i[3:3]),.IN2(s_fract_48_i[4:4]),.S(s_shr2[0:0]),.Q(n1693));
  MUX21X1 U2814(.IN1(n1693),.IN2(n1621),.S(n1237),.Q(n1622));
  MUX21X1 U2815(.IN1(s_fract_48_i[8:8]),.IN2(s_fract_48_i[7:7]),.S(n1240),.Q(n1695));
  MUX21X1 U2816(.IN1(n1226),.IN2(n1223),.S(n1240),.Q(n1694));
  MUX21X1 U2817(.IN1(n1695),.IN2(n1694),.S(n1237),.Q(n1720));
  MUX21X1 U2818(.IN1(n1622),.IN2(n1720),.S(s_shr2[2:2]),.Q(n1623));
  MUX21X1 U2819(.IN1(n1751),.IN2(n1623),.S(n1232),.Q(n1624));
  MUX21X1 U2820(.IN1(n1625),.IN2(n1624),.S(n1281),.Q(n1627));
  MUX21X1 U2821(.IN1(n1627),.IN2(n1686),.S(n1286),.Q(N3094));
  MUX21X1 U2822(.IN1(n1629),.IN2(n1390),.S(n1232),.Q(n1689));
  MUX21X1 U2823(.IN1(n1631),.IN2(n1630),.S(n1232),.Q(n1716));
  MUX21X1 U2824(.IN1(n1689),.IN2(n1432),.S(n1281),.Q(n1632));
  MUX21X1 U2825(.IN1(n1634),.IN2(n1385),.S(n1232),.Q(n1690));
  MUX21X1 U2826(.IN1(n1636),.IN2(n1635),.S(n1232),.Q(n1724));
  MUX21X1 U2827(.IN1(n1690),.IN2(n1423),.S(n1281),.Q(n1637));
  MUX21X1 U2828(.IN1(n1639),.IN2(n1383),.S(n1232),.Q(n1691));
  MUX21X1 U2829(.IN1(n1641),.IN2(n1640),.S(n1232),.Q(n1732));
  MUX21X1 U2830(.IN1(n1691),.IN2(n1419),.S(n1281),.Q(n1642));
  MUX21X1 U2831(.IN1(n1644),.IN2(n1356),.S(n1232),.Q(n1692));
  MUX21X1 U2832(.IN1(n1646),.IN2(n1645),.S(n1232),.Q(n1740));
  MUX21X1 U2833(.IN1(n1692),.IN2(n1415),.S(n1281),.Q(n1647));
  MUX21X1 U2834(.IN1(n1650),.IN2(n1649),.S(s_shr2[3:3]),.Q(n1746));
  MUX21X1 U2835(.IN1(n1704),.IN2(n1411),.S(n79),.Q(n1651));
  OR2X1 U2836(.IN1(n1652),.IN2(s_shr2[3:3]),.Q(n1705));
  MUX21X1 U2837(.IN1(n1654),.IN2(n1653),.S(s_shr2[3:3]),.Q(n1752));
  MUX21X1 U2838(.IN1(n1705),.IN2(n1406),.S(n1281),.Q(n1655));
  MUX21X1 U2839(.IN1(n1657),.IN2(n1398),.S(n79),.Q(n1658));
  MUX21X1 U2840(.IN1(n1660),.IN2(n1393),.S(n79),.Q(n1661));
  MUX21X1 U2841(.IN1(n1663),.IN2(n1389),.S(n79),.Q(n1664));
  MUX21X1 U2842(.IN1(n1666),.IN2(n1384),.S(n79),.Q(n1667));
  MUX21X1 U2843(.IN1(n1669),.IN2(n1668),.S(n1237),.Q(n1672));
  MUX21X1 U2844(.IN1(n1671),.IN2(n1670),.S(n1237),.Q(n1728));
  MUX21X1 U2845(.IN1(n1672),.IN2(n1728),.S(s_shr2[2:2]),.Q(n1673));
  MUX21X1 U2846(.IN1(n1674),.IN2(n1673),.S(n1232),.Q(n1675));
  MUX21X1 U2847(.IN1(n1676),.IN2(n1675),.S(n79),.Q(n1678));
  MUX21X1 U2848(.IN1(n1678),.IN2(n1687),.S(n1286),.Q(N3095));
  MUX21X1 U2849(.IN1(n1680),.IN2(n1382),.S(n1282),.Q(n1681));
  MUX21X1 U2850(.IN1(n1683),.IN2(n1355),.S(n1282),.Q(n1684));
  MUX21X1 U2851(.IN1(n1694),.IN2(n1693),.S(n1237),.Q(n1697));
  MUX21X1 U2852(.IN1(n1696),.IN2(n1695),.S(n1237),.Q(n1736));
  MUX21X1 U2853(.IN1(n1697),.IN2(n1736),.S(s_shr2[2:2]),.Q(n1698));
  MUX21X1 U2854(.IN1(n1699),.IN2(n1698),.S(n1232),.Q(n1701));
  MUX21X1 U2855(.IN1(n1701),.IN2(n1700),.S(n1280),.Q(n1703));
  MUX21X1 U2856(.IN1(n1703),.IN2(n1702),.S(n1286),.Q(N3096));
  MUX21X1 U2857(.IN1(n1713),.IN2(n1712),.S(n1235),.Q(n1714));
  MUX21X1 U2858(.IN1(n1715),.IN2(n1714),.S(n1232),.Q(n1717));
  MUX21X1 U2859(.IN1(n1717),.IN2(n1716),.S(n1280),.Q(n1719));
  MUX21X1 U2860(.IN1(n1719),.IN2(n1718),.S(n1286),.Q(N3097));
  MUX21X1 U2861(.IN1(n1721),.IN2(n1720),.S(n1235),.Q(n1722));
  MUX21X1 U2862(.IN1(n1723),.IN2(n1722),.S(n1232),.Q(n1725));
  MUX21X1 U2863(.IN1(n1725),.IN2(n1724),.S(n1280),.Q(n1727));
  MUX21X1 U2864(.IN1(n1727),.IN2(n1726),.S(n1286),.Q(N3098));
  MUX21X1 U2865(.IN1(n1729),.IN2(n1728),.S(n1235),.Q(n1730));
  MUX21X1 U2866(.IN1(n1731),.IN2(n1730),.S(n1232),.Q(n1733));
  MUX21X1 U2867(.IN1(n1733),.IN2(n1732),.S(n1280),.Q(n1735));
  MUX21X1 U2868(.IN1(n1735),.IN2(n1734),.S(n1286),.Q(N3099));
  MUX21X1 U2869(.IN1(n1737),.IN2(n1736),.S(n1235),.Q(n1738));
  MUX21X1 U2870(.IN1(n1739),.IN2(n1738),.S(n1232),.Q(n1741));
  MUX21X1 U2871(.IN1(n1741),.IN2(n1740),.S(n1280),.Q(n1743));
  MUX21X1 U2872(.IN1(n1743),.IN2(n1742),.S(n1286),.Q(N3100));
  MUX21X1 U2873(.IN1(n1745),.IN2(n1744),.S(s_shr2[3:3]),.Q(n1747));
  MUX21X1 U2874(.IN1(n1747),.IN2(n1746),.S(n1280),.Q(n1749));
  MUX21X1 U2875(.IN1(n1749),.IN2(n1748),.S(n1286),.Q(N3101));
  MUX21X1 U2876(.IN1(n1751),.IN2(n1750),.S(s_shr2[3:3]),.Q(n1753));
  MUX21X1 U2877(.IN1(n1753),.IN2(n1752),.S(n1280),.Q(n1755));
  MUX21X1 U2878(.IN1(n1755),.IN2(n1754),.S(n1286),.Q(N3102));
  OR2X1 U2879(.IN1(n1761),.IN2(n1264),.Q(n1764));
  OR2X1 U2880(.IN1(n1764),.IN2(n1267),.Q(n1823));
  OR2X1 U2881(.IN1(n1823),.IN2(n1271),.Q(n1785));
  OR2X1 U2882(.IN1(n1785),.IN2(n1274),.Q(n1868));
  MUX21X1 U2883(.IN1(s_fract_48_i[10:10]),.IN2(s_fract_48_i[9:9]),.S(n1260),.Q(n1756));
  MUX21X1 U2884(.IN1(s_fract_48_i[8:8]),.IN2(s_fract_48_i[7:7]),.S(n1260),.Q(n1757));
  MUX21X1 U2885(.IN1(n1506),.IN2(n1508),.S(s_shl2[1:1]),.Q(n1773));
  MUX21X1 U2886(.IN1(n1227),.IN2(n1220),.S(n1260),.Q(n1758));
  MUX21X1 U2887(.IN1(s_fract_48_i[4:4]),.IN2(s_fract_48_i[3:3]),.S(n1260),.Q(n1759));
  MUX21X1 U2888(.IN1(n1510),.IN2(n1512),.S(s_shl2[1:1]),.Q(n1775));
  MUX21X1 U2889(.IN1(n1773),.IN2(n1775),.S(n1267),.Q(n1793));
  MUX21X1 U2890(.IN1(n1514),.IN2(n1761),.S(n1264),.Q(n1774));
  OR2X1 U2891(.IN1(n1774),.IN2(n1267),.Q(n1794));
  MUX21X1 U2892(.IN1(n1793),.IN2(n1794),.S(n1268),.Q(n1835));
  OR2X1 U2893(.IN1(n1835),.IN2(n1274),.Q(n1952));
  MUX21X1 U2894(.IN1(s_fract_48_i[11:11]),.IN2(s_fract_48_i[10:10]),.S(n1260),.Q(n1765));
  MUX21X1 U2895(.IN1(s_fract_48_i[9:9]),.IN2(s_fract_48_i[8:8]),.S(n1260),.Q(n1767));
  MUX21X1 U2896(.IN1(n1765),.IN2(n1767),.S(n1263),.Q(n1777));
  MUX21X1 U2897(.IN1(s_fract_48_i[7:7]),.IN2(n1225),.S(n1260),.Q(n1766));
  MUX21X1 U2898(.IN1(n1222),.IN2(s_fract_48_i[4:4]),.S(n1260),.Q(n1770));
  MUX21X1 U2899(.IN1(n1766),.IN2(n1770),.S(s_shl2[1:1]),.Q(n1779));
  MUX21X1 U2900(.IN1(n1777),.IN2(n1779),.S(n1267),.Q(n1762));
  MUX21X1 U2901(.IN1(s_fract_48_i[3:3]),.IN2(s_fract_48_i[2:2]),.S(n1260),.Q(n1769));
  MUX21X1 U2902(.IN1(n1769),.IN2(n1772),.S(s_shl2[1:1]),.Q(n1778));
  MUX21X1 U2903(.IN1(n1503),.IN2(n1798),.S(n1268),.Q(n1840));
  OR2X1 U2904(.IN1(n1840),.IN2(n1274),.Q(n1961));
  MUX21X1 U2905(.IN1(n1210),.IN2(s_fract_48_i[11:11]),.S(n1260),.Q(n1763));
  MUX21X1 U2906(.IN1(n1499),.IN2(n1506),.S(s_shl2[1:1]),.Q(n1782));
  MUX21X1 U2907(.IN1(n1508),.IN2(n1510),.S(s_shl2[1:1]),.Q(n1784));
  MUX21X1 U2908(.IN1(n1782),.IN2(n1784),.S(n1267),.Q(n1803));
  MUX21X1 U2909(.IN1(n1512),.IN2(n1514),.S(s_shl2[1:1]),.Q(n1783));
  MUX21X1 U2910(.IN1(n1783),.IN2(n1764),.S(n1267),.Q(n1804));
  MUX21X1 U2911(.IN1(n1803),.IN2(n1804),.S(n1268),.Q(n1845));
  MUX21X1 U2912(.IN1(n1496),.IN2(n1287),.S(n1261),.Q(n1776));
  MUX21X1 U2913(.IN1(n1776),.IN2(n1505),.S(s_shl2[1:1]),.Q(n1788));
  MUX21X1 U2914(.IN1(n1767),.IN2(n1766),.S(n1265),.Q(n1768));
  MUX21X1 U2915(.IN1(n1788),.IN2(n1507),.S(n1267),.Q(n1808));
  MUX21X1 U2916(.IN1(n1770),.IN2(n1769),.S(n1265),.Q(n1771));
  MUX21X1 U2917(.IN1(n1511),.IN2(n1789),.S(n1267),.Q(n1809));
  MUX21X1 U2918(.IN1(n1808),.IN2(n1809),.S(n1268),.Q(n1850));
  MUX21X1 U2919(.IN1(n1493),.IN2(n1496),.S(n1261),.Q(n1781));
  MUX21X1 U2920(.IN1(n1781),.IN2(n1499),.S(n1265),.Q(n1792));
  MUX21X1 U2921(.IN1(n1792),.IN2(n1773),.S(s_shl2[2:2]),.Q(n1813));
  MUX21X1 U2922(.IN1(n1775),.IN2(n1774),.S(n1267),.Q(n1814));
  MUX21X1 U2923(.IN1(n1813),.IN2(n1814),.S(n1268),.Q(n1856));
  MUX21X1 U2924(.IN1(n1490),.IN2(n1493),.S(n1261),.Q(n1787));
  MUX21X1 U2925(.IN1(n1787),.IN2(n1776),.S(n1265),.Q(n1797));
  MUX21X1 U2926(.IN1(n1797),.IN2(n1504),.S(n1267),.Q(n1818));
  MUX21X1 U2927(.IN1(n1779),.IN2(n1778),.S(s_shl2[2:2]),.Q(n1780));
  MUX21X1 U2928(.IN1(n1818),.IN2(n1509),.S(n1268),.Q(n1861));
  MUX21X1 U2929(.IN1(n1487),.IN2(n1490),.S(n1261),.Q(n1791));
  MUX21X1 U2930(.IN1(n1791),.IN2(n1781),.S(n1265),.Q(n1802));
  MUX21X1 U2931(.IN1(n1802),.IN2(n1782),.S(s_shl2[2:2]),.Q(n1822));
  MUX21X1 U2932(.IN1(n1784),.IN2(n1783),.S(s_shl2[2:2]),.Q(n1824));
  MUX21X1 U2933(.IN1(n1822),.IN2(n1824),.S(n1268),.Q(n1866));
  MUX21X1 U2934(.IN1(n1866),.IN2(n1785),.S(n1272),.Q(n1786));
  MUX21X1 U2935(.IN1(n1485),.IN2(n1487),.S(n1261),.Q(n1796));
  MUX21X1 U2936(.IN1(n1796),.IN2(n1787),.S(n1265),.Q(n1807));
  MUX21X1 U2937(.IN1(n1807),.IN2(n1788),.S(s_shl2[2:2]),.Q(n1828));
  MUX21X1 U2938(.IN1(n1507),.IN2(n1511),.S(s_shl2[2:2]),.Q(n1830));
  MUX21X1 U2939(.IN1(n1828),.IN2(n1830),.S(n1268),.Q(n1874));
  OR2X1 U2940(.IN1(n1789),.IN2(n1267),.Q(n1829));
  OR2X1 U2941(.IN1(n1829),.IN2(n1271),.Q(n1800));
  MUX21X1 U2942(.IN1(n1874),.IN2(n1800),.S(n1272),.Q(n1790));
  MUX21X1 U2943(.IN1(n1288),.IN2(n1485),.S(n1261),.Q(n1801));
  MUX21X1 U2944(.IN1(n1801),.IN2(n1791),.S(n1265),.Q(n1812));
  MUX21X1 U2945(.IN1(n1812),.IN2(n1792),.S(s_shl2[2:2]),.Q(n1834));
  MUX21X1 U2946(.IN1(n1834),.IN2(n1793),.S(n1268),.Q(n1882));
  OR2X1 U2947(.IN1(n1794),.IN2(n1271),.Q(n1852));
  MUX21X1 U2948(.IN1(n1882),.IN2(n1852),.S(n1272),.Q(n1795));
  MUX21X1 U2949(.IN1(n1479),.IN2(n1288),.S(n1261),.Q(n1806));
  MUX21X1 U2950(.IN1(n1806),.IN2(n1796),.S(n1265),.Q(n1817));
  MUX21X1 U2951(.IN1(n1817),.IN2(n1797),.S(s_shl2[2:2]),.Q(n1839));
  MUX21X1 U2952(.IN1(n1839),.IN2(n1503),.S(n1269),.Q(n1890));
  OR2X1 U2953(.IN1(n1798),.IN2(n1271),.Q(n1892));
  MUX21X1 U2954(.IN1(n1890),.IN2(n1892),.S(n1272),.Q(n1799));
  OR2X1 U2955(.IN1(n1800),.IN2(n1274),.Q(n1876));
  MUX21X1 U2956(.IN1(n1478),.IN2(n1479),.S(n1261),.Q(n1811));
  MUX21X1 U2957(.IN1(n1811),.IN2(n1801),.S(n1265),.Q(n1821));
  MUX21X1 U2958(.IN1(n1821),.IN2(n1802),.S(s_shl2[2:2]),.Q(n1844));
  MUX21X1 U2959(.IN1(n1844),.IN2(n1803),.S(n1268),.Q(n1898));
  OR2X1 U2960(.IN1(n1804),.IN2(n1271),.Q(n1900));
  MUX21X1 U2961(.IN1(n1898),.IN2(n1900),.S(n1272),.Q(n1805));
  MUX21X1 U2962(.IN1(n1477),.IN2(n1478),.S(n1261),.Q(n1816));
  MUX21X1 U2963(.IN1(n1816),.IN2(n1806),.S(n1265),.Q(n1827));
  MUX21X1 U2964(.IN1(n1827),.IN2(n1807),.S(n1266),.Q(n1849));
  MUX21X1 U2965(.IN1(n1849),.IN2(n1808),.S(n1268),.Q(n1906));
  OR2X1 U2966(.IN1(n1809),.IN2(n1271),.Q(n1908));
  MUX21X1 U2967(.IN1(n1906),.IN2(n1908),.S(n1272),.Q(n1810));
  MUX21X1 U2968(.IN1(n1473),.IN2(n1477),.S(n1261),.Q(n1820));
  MUX21X1 U2969(.IN1(n1820),.IN2(n1811),.S(n1265),.Q(n1833));
  MUX21X1 U2970(.IN1(n1833),.IN2(n1812),.S(n1267),.Q(n1855));
  MUX21X1 U2971(.IN1(n1855),.IN2(n1813),.S(n1269),.Q(n1914));
  OR2X1 U2972(.IN1(n1814),.IN2(n1271),.Q(n1916));
  MUX21X1 U2973(.IN1(n1914),.IN2(n1916),.S(n1272),.Q(n1815));
  MUX21X1 U2974(.IN1(n1468),.IN2(n1473),.S(n1261),.Q(n1826));
  MUX21X1 U2975(.IN1(n1826),.IN2(n1816),.S(n1265),.Q(n1838));
  MUX21X1 U2976(.IN1(n1838),.IN2(n1817),.S(s_shl2[2:2]),.Q(n1860));
  MUX21X1 U2977(.IN1(n1860),.IN2(n1818),.S(n1269),.Q(n1922));
  OR2X1 U2978(.IN1(n1509),.IN2(n1271),.Q(n1924));
  MUX21X1 U2979(.IN1(n1922),.IN2(n1924),.S(n1272),.Q(n1819));
  MUX21X1 U2980(.IN1(n1291),.IN2(n1468),.S(n1261),.Q(n1832));
  MUX21X1 U2981(.IN1(n1832),.IN2(n1820),.S(n1264),.Q(n1843));
  MUX21X1 U2982(.IN1(n1843),.IN2(n1821),.S(n1266),.Q(n1865));
  MUX21X1 U2983(.IN1(n1865),.IN2(n1822),.S(n1269),.Q(n1932));
  MUX21X1 U2984(.IN1(n1824),.IN2(n1823),.S(n1269),.Q(n1934));
  MUX21X1 U2985(.IN1(n1932),.IN2(n1934),.S(n1272),.Q(n1825));
  MUX21X1 U2986(.IN1(n1463),.IN2(n1291),.S(n1262),.Q(n1837));
  MUX21X1 U2987(.IN1(n1837),.IN2(n1826),.S(n1264),.Q(n1848));
  MUX21X1 U2988(.IN1(n1848),.IN2(n1827),.S(n1266),.Q(n1873));
  MUX21X1 U2989(.IN1(n1873),.IN2(n1828),.S(n1269),.Q(n1941));
  MUX21X1 U2990(.IN1(n1830),.IN2(n1829),.S(n1269),.Q(n1943));
  MUX21X1 U2991(.IN1(n1941),.IN2(n1943),.S(n1272),.Q(n1831));
  MUX21X1 U2992(.IN1(n1462),.IN2(n1463),.S(n1262),.Q(n1842));
  MUX21X1 U2993(.IN1(n1842),.IN2(n1832),.S(n1264),.Q(n1854));
  MUX21X1 U2994(.IN1(n1854),.IN2(n1833),.S(n1267),.Q(n1881));
  MUX21X1 U2995(.IN1(n1881),.IN2(n1834),.S(n1269),.Q(n1950));
  MUX21X1 U2996(.IN1(n1950),.IN2(n1835),.S(n1272),.Q(n1836));
  MUX21X1 U2997(.IN1(n1461),.IN2(n1462),.S(n1262),.Q(n1847));
  MUX21X1 U2998(.IN1(n1847),.IN2(n1837),.S(n1264),.Q(n1859));
  MUX21X1 U2999(.IN1(n1859),.IN2(n1838),.S(n1266),.Q(n1889));
  MUX21X1 U3000(.IN1(n1889),.IN2(n1839),.S(n1269),.Q(n1959));
  MUX21X1 U3001(.IN1(n1959),.IN2(n1840),.S(n1272),.Q(n1841));
  MUX21X1 U3002(.IN1(n1460),.IN2(n1461),.S(n1262),.Q(n1853));
  MUX21X1 U3003(.IN1(n1853),.IN2(n1842),.S(n1264),.Q(n1864));
  MUX21X1 U3004(.IN1(n1864),.IN2(n1843),.S(n1267),.Q(n1897));
  MUX21X1 U3005(.IN1(n1897),.IN2(n1844),.S(n1269),.Q(n1969));
  MUX21X1 U3006(.IN1(n1969),.IN2(n1845),.S(n1273),.Q(n1846));
  MUX21X1 U3007(.IN1(n1458),.IN2(n1460),.S(n1262),.Q(n1858));
  MUX21X1 U3008(.IN1(n1858),.IN2(n1847),.S(n1264),.Q(n1872));
  MUX21X1 U3009(.IN1(n1872),.IN2(n1848),.S(s_shl2[2:2]),.Q(n1905));
  MUX21X1 U3010(.IN1(n1905),.IN2(n1849),.S(n1269),.Q(n1978));
  MUX21X1 U3011(.IN1(n1978),.IN2(n1850),.S(n1273),.Q(n1851));
  OR2X1 U3012(.IN1(n1852),.IN2(n1274),.Q(n1884));
  MUX21X1 U3013(.IN1(n1292),.IN2(n1458),.S(n1262),.Q(n1863));
  MUX21X1 U3014(.IN1(n1863),.IN2(n1853),.S(n1264),.Q(n1880));
  MUX21X1 U3015(.IN1(n1880),.IN2(n1854),.S(s_shl2[2:2]),.Q(n1913));
  MUX21X1 U3016(.IN1(n1913),.IN2(n1855),.S(n1269),.Q(n1988));
  MUX21X1 U3017(.IN1(n1988),.IN2(n1856),.S(n1273),.Q(n1857));
  MUX21X1 U3018(.IN1(n1449),.IN2(n1292),.S(n1262),.Q(n1871));
  MUX21X1 U3019(.IN1(n1871),.IN2(n1858),.S(n1264),.Q(n1888));
  MUX21X1 U3020(.IN1(n1888),.IN2(n1859),.S(s_shl2[2:2]),.Q(n1921));
  MUX21X1 U3021(.IN1(n1921),.IN2(n1860),.S(n1270),.Q(n1998));
  MUX21X1 U3022(.IN1(n1998),.IN2(n1861),.S(n1273),.Q(n1862));
  MUX21X1 U3023(.IN1(n1446),.IN2(n1449),.S(n1262),.Q(n1879));
  MUX21X1 U3024(.IN1(n1879),.IN2(n1863),.S(n1264),.Q(n1896));
  MUX21X1 U3025(.IN1(n1896),.IN2(n1864),.S(s_shl2[2:2]),.Q(n1931));
  MUX21X1 U3026(.IN1(n1931),.IN2(n1865),.S(n1270),.Q(n1867));
  MUX21X1 U3027(.IN1(n1867),.IN2(n1866),.S(n1273),.Q(n1869));
  MUX21X1 U3028(.IN1(n1869),.IN2(n1868),.S(n1277),.Q(n1870));
  MUX21X1 U3029(.IN1(n1442),.IN2(n1446),.S(n1262),.Q(n1887));
  MUX21X1 U3030(.IN1(n1887),.IN2(n1871),.S(n1264),.Q(n1904));
  MUX21X1 U3031(.IN1(n1904),.IN2(n1872),.S(s_shl2[2:2]),.Q(n1940));
  MUX21X1 U3032(.IN1(n1940),.IN2(n1873),.S(n1270),.Q(n1875));
  MUX21X1 U3033(.IN1(n1875),.IN2(n1874),.S(n1273),.Q(n1877));
  MUX21X1 U3034(.IN1(n1877),.IN2(n1876),.S(n1277),.Q(n1878));
  MUX21X1 U3035(.IN1(s_fract_48_i[34:34]),.IN2(s_fract_48_i[33:33]),.S(n1262),.Q(n1895));
  MUX21X1 U3036(.IN1(n1438),.IN2(n1879),.S(n1264),.Q(n1912));
  MUX21X1 U3037(.IN1(n1912),.IN2(n1880),.S(s_shl2[2:2]),.Q(n1949));
  MUX21X1 U3038(.IN1(n1949),.IN2(n1881),.S(n1270),.Q(n1883));
  MUX21X1 U3039(.IN1(n1883),.IN2(n1882),.S(n1273),.Q(n1885));
  MUX21X1 U3040(.IN1(n1885),.IN2(n1884),.S(n1277),.Q(n1886));
  MUX21X1 U3041(.IN1(s_fract_48_i[35:35]),.IN2(s_fract_48_i[34:34]),.S(n1262),.Q(n1903));
  MUX21X1 U3042(.IN1(n1434),.IN2(n1887),.S(n1264),.Q(n1920));
  MUX21X1 U3043(.IN1(n1920),.IN2(n1888),.S(n1266),.Q(n1958));
  MUX21X1 U3044(.IN1(n1958),.IN2(n1889),.S(n1270),.Q(n1891));
  MUX21X1 U3045(.IN1(n1891),.IN2(n1890),.S(n1273),.Q(n1893));
  OR2X1 U3046(.IN1(n1892),.IN2(n1273),.Q(n1927));
  MUX21X1 U3047(.IN1(n1893),.IN2(n1927),.S(n1277),.Q(n1894));
  MUX21X1 U3048(.IN1(s_fract_48_i[36:36]),.IN2(s_fract_48_i[35:35]),.S(n1262),.Q(n1911));
  MUX21X1 U3049(.IN1(n1911),.IN2(n1895),.S(n1263),.Q(n1929));
  MUX21X1 U3050(.IN1(n1426),.IN2(n1896),.S(n1266),.Q(n1967));
  MUX21X1 U3051(.IN1(n1967),.IN2(n1897),.S(n1270),.Q(n1899));
  MUX21X1 U3052(.IN1(n1899),.IN2(n1898),.S(n1273),.Q(n1901));
  OR2X1 U3053(.IN1(n1900),.IN2(n1274),.Q(n2002));
  MUX21X1 U3054(.IN1(n1901),.IN2(n2002),.S(n1277),.Q(n1902));
  MUX21X1 U3055(.IN1(s_fract_48_i[37:37]),.IN2(s_fract_48_i[36:36]),.S(n55),.Q(n1919));
  MUX21X1 U3056(.IN1(n1919),.IN2(n1903),.S(n1263),.Q(n1938));
  MUX21X1 U3057(.IN1(n1422),.IN2(n1904),.S(n1266),.Q(n1976));
  MUX21X1 U3058(.IN1(n1976),.IN2(n1905),.S(n1270),.Q(n1907));
  MUX21X1 U3059(.IN1(n1907),.IN2(n1906),.S(n1273),.Q(n1909));
  OR2X1 U3060(.IN1(n1908),.IN2(n1274),.Q(n2003));
  MUX21X1 U3061(.IN1(n1909),.IN2(n2003),.S(n1277),.Q(n1910));
  MUX21X1 U3062(.IN1(s_fract_48_i[38:38]),.IN2(s_fract_48_i[37:37]),.S(n55),.Q(n1928));
  MUX21X1 U3063(.IN1(n1928),.IN2(n1911),.S(n1263),.Q(n1947));
  MUX21X1 U3064(.IN1(n1418),.IN2(n1912),.S(n1266),.Q(n1986));
  MUX21X1 U3065(.IN1(n1986),.IN2(n1913),.S(n1270),.Q(n1915));
  MUX21X1 U3066(.IN1(n1915),.IN2(n1914),.S(n1273),.Q(n1917));
  OR2X1 U3067(.IN1(n1916),.IN2(n1274),.Q(n2004));
  MUX21X1 U3068(.IN1(n1917),.IN2(n2004),.S(n1278),.Q(n1918));
  MUX21X1 U3069(.IN1(s_fract_48_i[39:39]),.IN2(s_fract_48_i[38:38]),.S(n55),.Q(n1937));
  MUX21X1 U3070(.IN1(n1937),.IN2(n1919),.S(n1263),.Q(n1956));
  MUX21X1 U3071(.IN1(n1414),.IN2(n1920),.S(n1266),.Q(n1996));
  MUX21X1 U3072(.IN1(n1996),.IN2(n1921),.S(n1270),.Q(n1923));
  MUX21X1 U3073(.IN1(n1923),.IN2(n1922),.S(n1273),.Q(n1925));
  OR2X1 U3074(.IN1(n1924),.IN2(n1274),.Q(n2005));
  MUX21X1 U3075(.IN1(n1925),.IN2(n2005),.S(n1278),.Q(n1926));
  MUX21X1 U3076(.IN1(s_fract_48_i[40:40]),.IN2(s_fract_48_i[39:39]),.S(n55),.Q(n1946));
  MUX21X1 U3077(.IN1(n1946),.IN2(n1928),.S(n1263),.Q(n1965));
  MUX21X1 U3078(.IN1(n1965),.IN2(n1929),.S(n1266),.Q(n1930));
  MUX21X1 U3079(.IN1(n1408),.IN2(n1931),.S(n1270),.Q(n1933));
  MUX21X1 U3080(.IN1(n1933),.IN2(n1932),.S(n1273),.Q(n1935));
  OR2X1 U3081(.IN1(n1934),.IN2(n1274),.Q(n2006));
  MUX21X1 U3082(.IN1(n1935),.IN2(n2006),.S(n1278),.Q(n1936));
  MUX21X1 U3083(.IN1(s_fract_48_i[41:41]),.IN2(s_fract_48_i[40:40]),.S(n55),.Q(n1955));
  MUX21X1 U3084(.IN1(n1955),.IN2(n1937),.S(n1263),.Q(n1974));
  MUX21X1 U3085(.IN1(n1974),.IN2(n1938),.S(n1266),.Q(n1939));
  MUX21X1 U3086(.IN1(n1401),.IN2(n1940),.S(n1270),.Q(n1942));
  MUX21X1 U3087(.IN1(n1942),.IN2(n1941),.S(n1273),.Q(n1944));
  OR2X1 U3088(.IN1(n1943),.IN2(n1274),.Q(n2007));
  MUX21X1 U3089(.IN1(n1944),.IN2(n2007),.S(n1278),.Q(n1945));
  MUX21X1 U3090(.IN1(n1230),.IN2(s_fract_48_i[41:41]),.S(n55),.Q(n1964));
  MUX21X1 U3091(.IN1(n1964),.IN2(n1946),.S(n1263),.Q(n1984));
  MUX21X1 U3092(.IN1(n1984),.IN2(n1947),.S(n1266),.Q(n1948));
  MUX21X1 U3093(.IN1(n1396),.IN2(n1949),.S(n1271),.Q(n1951));
  MUX21X1 U3094(.IN1(n1951),.IN2(n1950),.S(n1273),.Q(n1953));
  MUX21X1 U3095(.IN1(n1953),.IN2(n1952),.S(n1278),.Q(n1954));
  MUX21X1 U3096(.IN1(s_fract_48_i[43:43]),.IN2(n1228),.S(n55),.Q(n1973));
  MUX21X1 U3097(.IN1(n1973),.IN2(n1955),.S(n1263),.Q(n1994));
  MUX21X1 U3098(.IN1(n1994),.IN2(n1956),.S(n1266),.Q(n1957));
  MUX21X1 U3099(.IN1(n1392),.IN2(n1958),.S(n1271),.Q(n1960));
  MUX21X1 U3100(.IN1(n1960),.IN2(n1959),.S(n1273),.Q(n1962));
  MUX21X1 U3101(.IN1(n1962),.IN2(n1961),.S(n1278),.Q(n1963));
  MUX21X1 U3102(.IN1(s_fract_48_i[43:43]),.IN2(s_fract_48_i[44:44]),.S(n76),.Q(n1982));
  MUX21X1 U3103(.IN1(n1982),.IN2(n1964),.S(n1263),.Q(n1966));
  MUX21X1 U3104(.IN1(n1966),.IN2(n1965),.S(n1266),.Q(n1968));
  MUX21X1 U3105(.IN1(n1968),.IN2(n1425),.S(n1271),.Q(n1970));
  MUX21X1 U3106(.IN1(n1970),.IN2(n1459),.S(n1273),.Q(n1972));
  MUX21X1 U3107(.IN1(n1972),.IN2(n1971),.S(n1278),.Q(N3185));
  MUX21X1 U3108(.IN1(s_fract_48_i[44:44]),.IN2(s_fract_48_i[45:45]),.S(n76),.Q(n1992));
  MUX21X1 U3109(.IN1(n1992),.IN2(n1973),.S(n1263),.Q(n1975));
  MUX21X1 U3110(.IN1(n1975),.IN2(n1974),.S(n1266),.Q(n1977));
  MUX21X1 U3111(.IN1(n1977),.IN2(n1421),.S(n1271),.Q(n1979));
  MUX21X1 U3112(.IN1(n1979),.IN2(n1457),.S(n1273),.Q(n1981));
  MUX21X1 U3113(.IN1(n1981),.IN2(n1980),.S(n1278),.Q(N3186));
  MUX21X1 U3114(.IN1(n1205),.IN2(s_fract_48_i[45:45]),.S(n55),.Q(n1983));
  MUX21X1 U3115(.IN1(n1983),.IN2(n1982),.S(n1263),.Q(n1985));
  MUX21X1 U3116(.IN1(n1985),.IN2(n1984),.S(n1266),.Q(n1987));
  MUX21X1 U3117(.IN1(n1987),.IN2(n1417),.S(n1270),.Q(n1989));
  MUX21X1 U3118(.IN1(n1989),.IN2(n1452),.S(n1273),.Q(n1991));
  MUX21X1 U3119(.IN1(n1991),.IN2(n1990),.S(n1278),.Q(N3187));
  MUX21X1 U3120(.IN1(N2993),.IN2(n1205),.S(n55),.Q(n1993));
  MUX21X1 U3121(.IN1(n1993),.IN2(n1992),.S(n1263),.Q(n1995));
  MUX21X1 U3122(.IN1(n1995),.IN2(n1994),.S(s_shl2[2:2]),.Q(n1997));
  MUX21X1 U3123(.IN1(n1997),.IN2(n1413),.S(n1268),.Q(n1999));
  MUX21X1 U3124(.IN1(n1999),.IN2(n1448),.S(n1272),.Q(n2001));
  MUX21X1 U3125(.IN1(n2001),.IN2(n2000),.S(n1278),.Q(N3188));
endmodule
module pre_norm_div_DW01_add_3_inj (A,B,CI,SUM,CO);
input [9:0] A ;
input [9:0] B ;
output [9:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire [9:1] carry ;
// instances
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(carry[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  XOR2X1 U2(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
  XOR2X1 U3(.IN1(B[9:9]),.IN2(carry[9:9]),.Q(SUM[9:9]));
endmodule
module pre_norm_div_DW01_add_2_inj (A,B,CI,SUM,CO);
input [9:0] A ;
input [9:0] B ;
output [9:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire [9:1] carry ;
// instances
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  AND2X1 U2(.IN1(A[6:6]),.IN2(carry[6:6]),.Q(n2));
  AND2X1 U3(.IN1(A[7:7]),.IN2(n2),.Q(n3));
  AND2X1 U4(.IN1(A[8:8]),.IN2(n3),.Q(n4));
  XOR2X1 U5(.IN1(A[9:9]),.IN2(n4),.Q(SUM[9:9]));
  XOR2X1 U6(.IN1(A[8:8]),.IN2(n3),.Q(SUM[8:8]));
  XOR2X1 U7(.IN1(A[7:7]),.IN2(n2),.Q(SUM[7:7]));
  XOR2X1 U8(.IN1(A[6:6]),.IN2(carry[6:6]),.Q(SUM[6:6]));
  XOR2X1 U9(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module pre_norm_div_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [9:0] A ;
input [9:0] B ;
output [9:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire [10:0] carry ;
// instances
  FADDX1 U2_5(.A(A[5:5]),.B(n8),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n9),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n12),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n11),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n10),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  INVX0 U1(.INP(A[6:6]),.ZN(n3));
  INVX0 U2(.INP(A[7:7]),.ZN(n5));
  INVX0 U3(.INP(carry[6:6]),.ZN(n4));
  INVX0 U4(.INP(B[4:4]),.ZN(n9));
  INVX0 U5(.INP(B[3:3]),.ZN(n12));
  INVX0 U6(.INP(B[2:2]),.ZN(n11));
  NAND2X0 U7(.IN1(n7),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U8(.INP(B[1:1]),.ZN(n10));
  INVX0 U9(.INP(A[0:0]),.ZN(n7));
  INVX0 U10(.INP(B[5:5]),.ZN(n8));
  AND2X1 U11(.IN1(n3),.IN2(n4),.Q(n1));
  AND2X1 U12(.IN1(n5),.IN2(n1),.Q(n2));
  NAND2X0 U13(.IN1(n6),.IN2(n2),.QN(carry[9:9]));
  INVX0 U14(.INP(A[8:8]),.ZN(n6));
  XNOR2X1 U15(.IN1(carry[9:9]),.IN2(A[9:9]),.Q(DIFF[9:9]));
  XOR2X1 U16(.IN1(n4),.IN2(A[6:6]),.Q(DIFF[6:6]));
  XOR2X1 U17(.IN1(n1),.IN2(A[7:7]),.Q(DIFF[7:7]));
  XOR2X1 U18(.IN1(n2),.IN2(A[8:8]),.Q(DIFF[8:8]));
  XOR2X1 U19(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module pre_norm_div_inj (clk_i,opa_i,opb_i,exp_10_o,dvdnd_50_o,dvsor_27_o,p_desc1176_p_O_DFFX1,p_desc1177_p_O_DFFX1,p_desc1178_p_O_DFFX1,p_desc1179_p_O_DFFX1,p_desc1180_p_O_DFFX1,p_desc1181_p_O_DFFX1,p_desc1182_p_O_DFFX1,p_desc1183_p_O_DFFX1,p_desc1184_p_O_DFFX1,p_desc1185_p_O_DFFX1,p_desc1186_p_O_DFFX1,p_desc1187_p_O_DFFX1,p_desc1188_p_O_DFFX1,p_desc1189_p_O_DFFX1,p_desc1190_p_O_DFFX1,p_desc1191_p_O_DFFX1,p_desc1192_p_O_DFFX1,p_desc1193_p_O_DFFX1,p_desc1194_p_O_DFFX1,p_desc1195_p_O_DFFX1,p_desc1196_p_O_DFFX1,p_desc1197_p_O_DFFX1,p_desc1198_p_O_DFFX1,p_desc1199_p_O_DFFX1,p_desc1200_p_O_DFFX1,p_desc1201_p_O_DFFX1,p_desc1202_p_O_DFFX1,p_desc1203_p_O_DFFX1,p_desc1204_p_O_DFFX1,p_desc1205_p_O_DFFX1,p_desc1206_p_O_DFFX1,p_desc1207_p_O_DFFX1,p_desc1208_p_O_DFFX1,p_desc1209_p_O_DFFX1,p_desc1210_p_O_DFFX1,p_desc1211_p_O_DFFX1,p_desc1212_p_O_DFFX1,p_desc1213_p_O_DFFX1);
input [31:0] opa_i ;
input [31:0] opb_i ;
output [9:0] exp_10_o ;
output [49:0] dvdnd_50_o ;
output [26:0] dvsor_27_o ;
input clk_i ;
wire N192 ;
wire N199 ;
wire N229 ;
wire N230 ;
wire N231 ;
wire N238 ;
wire N239 ;
wire N240 ;
wire N241 ;
wire N243 ;
wire N244 ;
wire N245 ;
wire N246 ;
wire N253 ;
wire N254 ;
wire N255 ;
wire N256 ;
wire N257 ;
wire N259 ;
wire N260 ;
wire N261 ;
wire N262 ;
wire N263 ;
wire N270 ;
wire N271 ;
wire N272 ;
wire N273 ;
wire N274 ;
wire N275 ;
wire N276 ;
wire N277 ;
wire N278 ;
wire N279 ;
wire N280 ;
wire N287 ;
wire N288 ;
wire N289 ;
wire N290 ;
wire N291 ;
wire N292 ;
wire N293 ;
wire N294 ;
wire N295 ;
wire N296 ;
wire N297 ;
wire N298 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N308 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N313 ;
wire N314 ;
wire N315 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N324 ;
wire N325 ;
wire N326 ;
wire N327 ;
wire N328 ;
wire N329 ;
wire N330 ;
wire N331 ;
wire N332 ;
wire N338 ;
wire N339 ;
wire N340 ;
wire N341 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N345 ;
wire N346 ;
wire N347 ;
wire N348 ;
wire N349 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N361 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N365 ;
wire N366 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N377 ;
wire N378 ;
wire N379 ;
wire N380 ;
wire N381 ;
wire N382 ;
wire N383 ;
wire N389 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N394 ;
wire N395 ;
wire N396 ;
wire N397 ;
wire N398 ;
wire N399 ;
wire N400 ;
wire N406 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N411 ;
wire N412 ;
wire N413 ;
wire N414 ;
wire N415 ;
wire N416 ;
wire N417 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N433 ;
wire N434 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N450 ;
wire N451 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N462 ;
wire N463 ;
wire N464 ;
wire N465 ;
wire N466 ;
wire N467 ;
wire N468 ;
wire N474 ;
wire N475 ;
wire N476 ;
wire N477 ;
wire N478 ;
wire N479 ;
wire N480 ;
wire N481 ;
wire N482 ;
wire N483 ;
wire N484 ;
wire N485 ;
wire N491 ;
wire N492 ;
wire N493 ;
wire N494 ;
wire N495 ;
wire N496 ;
wire N497 ;
wire N498 ;
wire N499 ;
wire N500 ;
wire N501 ;
wire N502 ;
wire N508 ;
wire N509 ;
wire N510 ;
wire N511 ;
wire N512 ;
wire N513 ;
wire N514 ;
wire N515 ;
wire N516 ;
wire N517 ;
wire N518 ;
wire N519 ;
wire N525 ;
wire N526 ;
wire N527 ;
wire N528 ;
wire N529 ;
wire N530 ;
wire N531 ;
wire N532 ;
wire N533 ;
wire N534 ;
wire N535 ;
wire N536 ;
wire N542 ;
wire N543 ;
wire N544 ;
wire N545 ;
wire N546 ;
wire N547 ;
wire N548 ;
wire N549 ;
wire N550 ;
wire N551 ;
wire N552 ;
wire N553 ;
wire N559 ;
wire N560 ;
wire N561 ;
wire N562 ;
wire N563 ;
wire N564 ;
wire N892 ;
wire N893 ;
wire N894 ;
wire N901 ;
wire N902 ;
wire N903 ;
wire N904 ;
wire N906 ;
wire N907 ;
wire N908 ;
wire N909 ;
wire N916 ;
wire N917 ;
wire N918 ;
wire N919 ;
wire N920 ;
wire N922 ;
wire N923 ;
wire N924 ;
wire N925 ;
wire N926 ;
wire N933 ;
wire N934 ;
wire N935 ;
wire N936 ;
wire N937 ;
wire N938 ;
wire N939 ;
wire N940 ;
wire N941 ;
wire N942 ;
wire N943 ;
wire N950 ;
wire N951 ;
wire N952 ;
wire N953 ;
wire N954 ;
wire N955 ;
wire N956 ;
wire N957 ;
wire N958 ;
wire N959 ;
wire N960 ;
wire N961 ;
wire N967 ;
wire N968 ;
wire N969 ;
wire N970 ;
wire N971 ;
wire N972 ;
wire N973 ;
wire N974 ;
wire N975 ;
wire N976 ;
wire N977 ;
wire N978 ;
wire N984 ;
wire N985 ;
wire N986 ;
wire N987 ;
wire N988 ;
wire N989 ;
wire N990 ;
wire N991 ;
wire N992 ;
wire N993 ;
wire N994 ;
wire N995 ;
wire N1001 ;
wire N1002 ;
wire N1003 ;
wire N1004 ;
wire N1005 ;
wire N1006 ;
wire N1007 ;
wire N1008 ;
wire N1009 ;
wire N1010 ;
wire N1011 ;
wire N1012 ;
wire N1018 ;
wire N1019 ;
wire N1020 ;
wire N1021 ;
wire N1022 ;
wire N1023 ;
wire N1024 ;
wire N1025 ;
wire N1026 ;
wire N1027 ;
wire N1028 ;
wire N1029 ;
wire N1035 ;
wire N1036 ;
wire N1037 ;
wire N1038 ;
wire N1039 ;
wire N1040 ;
wire N1041 ;
wire N1042 ;
wire N1043 ;
wire N1044 ;
wire N1045 ;
wire N1046 ;
wire N1052 ;
wire N1053 ;
wire N1054 ;
wire N1055 ;
wire N1056 ;
wire N1057 ;
wire N1058 ;
wire N1059 ;
wire N1060 ;
wire N1061 ;
wire N1062 ;
wire N1063 ;
wire N1069 ;
wire N1070 ;
wire N1071 ;
wire N1072 ;
wire N1073 ;
wire N1074 ;
wire N1075 ;
wire N1076 ;
wire N1077 ;
wire N1078 ;
wire N1079 ;
wire N1080 ;
wire N1086 ;
wire N1087 ;
wire N1088 ;
wire N1089 ;
wire N1090 ;
wire N1091 ;
wire N1092 ;
wire N1093 ;
wire N1094 ;
wire N1095 ;
wire N1096 ;
wire N1097 ;
wire N1103 ;
wire N1104 ;
wire N1105 ;
wire N1106 ;
wire N1107 ;
wire N1108 ;
wire N1109 ;
wire N1110 ;
wire N1111 ;
wire N1112 ;
wire N1113 ;
wire N1114 ;
wire N1120 ;
wire N1121 ;
wire N1122 ;
wire N1123 ;
wire N1124 ;
wire N1125 ;
wire N1126 ;
wire N1127 ;
wire N1128 ;
wire N1129 ;
wire N1130 ;
wire N1131 ;
wire N1137 ;
wire N1138 ;
wire N1139 ;
wire N1140 ;
wire N1141 ;
wire N1142 ;
wire N1143 ;
wire N1144 ;
wire N1145 ;
wire N1146 ;
wire N1147 ;
wire N1148 ;
wire N1154 ;
wire N1155 ;
wire N1156 ;
wire N1157 ;
wire N1158 ;
wire N1159 ;
wire N1160 ;
wire N1161 ;
wire N1162 ;
wire N1163 ;
wire N1164 ;
wire N1165 ;
wire N1171 ;
wire N1172 ;
wire N1173 ;
wire N1174 ;
wire N1175 ;
wire N1176 ;
wire N1177 ;
wire N1178 ;
wire N1179 ;
wire N1180 ;
wire N1181 ;
wire N1182 ;
wire N1188 ;
wire N1189 ;
wire N1190 ;
wire N1191 ;
wire N1192 ;
wire N1193 ;
wire N1194 ;
wire N1195 ;
wire N1196 ;
wire N1197 ;
wire N1198 ;
wire N1199 ;
wire N1205 ;
wire N1206 ;
wire N1207 ;
wire N1208 ;
wire N1209 ;
wire N1210 ;
wire N1211 ;
wire N1212 ;
wire N1213 ;
wire N1214 ;
wire N1215 ;
wire N1216 ;
wire N1222 ;
wire N1223 ;
wire N1224 ;
wire N1225 ;
wire N1226 ;
wire N1227 ;
wire N1526 ;
wire N1527 ;
wire N1528 ;
wire N1529 ;
wire N1530 ;
wire N1531 ;
wire N1532 ;
wire N1533 ;
wire N1534 ;
wire N1535 ;
wire N1536 ;
wire N1537 ;
wire N1538 ;
wire N1539 ;
wire N1540 ;
wire N1541 ;
wire N1542 ;
wire N1543 ;
wire N1574 ;
wire N1575 ;
wire N1576 ;
wire N1577 ;
wire N1578 ;
wire N1579 ;
wire N1580 ;
wire N1581 ;
wire N1582 ;
wire N1583 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire N1573 ;
wire N1572 ;
wire N1571 ;
wire N1570 ;
wire N1569 ;
wire N1568 ;
wire N1567 ;
wire N1566 ;
wire N1565 ;
wire N1564 ;
wire N1562 ;
wire N1561 ;
wire N1553 ;
wire N1552 ;
wire N1551 ;
wire N1550 ;
wire N1549 ;
wire N1548 ;
wire N1547 ;
wire N1546 ;
wire N1545 ;
wire N1544 ;
wire \add_117/carry[7]  ;
wire \add_117/carry[6]  ;
wire \add_117/carry[5]  ;
wire \add_117/carry[4]  ;
wire \add_117/carry[3]  ;
wire \add_117/carry[2]  ;
wire \add_117/carry[1]  ;
wire \add_117/B[0]  ;
wire \add_116/carry[7]  ;
wire \add_116/carry[6]  ;
wire \add_116/carry[5]  ;
wire \add_116/carry[4]  ;
wire \add_116/carry[3]  ;
wire \add_116/carry[2]  ;
wire \add_116/carry[1]  ;
wire \add_116/B[0]  ;
wire \add_90_I24_L14036_C104/carry[5]  ;
wire \add_90_I24_L14036_C104/carry[4]  ;
wire \add_90_I24_L14036_C104/carry[3]  ;
wire \add_90_I24_L14036_C104/carry[2]  ;
wire \add_90_I23_L14036_C104/carry[5]  ;
wire \add_90_I23_L14036_C104/carry[4]  ;
wire \add_90_I23_L14036_C104/carry[3]  ;
wire \add_90_I23_L14036_C104/carry[2]  ;
wire \add_90_I22_L14036_C104/carry[5]  ;
wire \add_90_I22_L14036_C104/carry[4]  ;
wire \add_90_I22_L14036_C104/carry[3]  ;
wire \add_90_I22_L14036_C104/carry[2]  ;
wire \add_90_I21_L14036_C104/carry[5]  ;
wire \add_90_I21_L14036_C104/carry[4]  ;
wire \add_90_I21_L14036_C104/carry[3]  ;
wire \add_90_I21_L14036_C104/carry[2]  ;
wire \add_90_I20_L14036_C104/carry[5]  ;
wire \add_90_I20_L14036_C104/carry[4]  ;
wire \add_90_I20_L14036_C104/carry[3]  ;
wire \add_90_I20_L14036_C104/carry[2]  ;
wire \add_90_I19_L14036_C104/carry[5]  ;
wire \add_90_I19_L14036_C104/carry[4]  ;
wire \add_90_I19_L14036_C104/carry[3]  ;
wire \add_90_I19_L14036_C104/carry[2]  ;
wire \add_90_I18_L14036_C104/carry[5]  ;
wire \add_90_I18_L14036_C104/carry[4]  ;
wire \add_90_I18_L14036_C104/carry[3]  ;
wire \add_90_I18_L14036_C104/carry[2]  ;
wire \add_90_I17_L14036_C104/carry[5]  ;
wire \add_90_I17_L14036_C104/carry[4]  ;
wire \add_90_I17_L14036_C104/carry[3]  ;
wire \add_90_I17_L14036_C104/carry[2]  ;
wire \add_90_I16_L14036_C104/carry[5]  ;
wire \add_90_I16_L14036_C104/carry[4]  ;
wire \add_90_I16_L14036_C104/carry[3]  ;
wire \add_90_I16_L14036_C104/carry[2]  ;
wire \add_90_I15_L14036_C104/carry[5]  ;
wire \add_90_I15_L14036_C104/carry[4]  ;
wire \add_90_I15_L14036_C104/carry[3]  ;
wire \add_90_I15_L14036_C104/carry[2]  ;
wire \add_90_I14_L14036_C104/carry[5]  ;
wire \add_90_I14_L14036_C104/carry[4]  ;
wire \add_90_I14_L14036_C104/carry[3]  ;
wire \add_90_I14_L14036_C104/carry[2]  ;
wire \add_90_I13_L14036_C104/carry[5]  ;
wire \add_90_I13_L14036_C104/carry[4]  ;
wire \add_90_I13_L14036_C104/carry[3]  ;
wire \add_90_I13_L14036_C104/carry[2]  ;
wire \add_90_I12_L14036_C104/carry[5]  ;
wire \add_90_I12_L14036_C104/carry[4]  ;
wire \add_90_I12_L14036_C104/carry[3]  ;
wire \add_90_I12_L14036_C104/carry[2]  ;
wire \add_90_I11_L14036_C104/carry[5]  ;
wire \add_90_I11_L14036_C104/carry[4]  ;
wire \add_90_I11_L14036_C104/carry[3]  ;
wire \add_90_I11_L14036_C104/carry[2]  ;
wire \add_90_I10_L14036_C104/carry[5]  ;
wire \add_90_I10_L14036_C104/carry[4]  ;
wire \add_90_I10_L14036_C104/carry[3]  ;
wire \add_90_I10_L14036_C104/carry[2]  ;
wire \add_90_I9_L14036_C104/carry[5]  ;
wire \add_90_I9_L14036_C104/carry[4]  ;
wire \add_90_I9_L14036_C104/carry[3]  ;
wire \add_90_I9_L14036_C104/carry[2]  ;
wire \add_90_I8_L14036_C104/carry[5]  ;
wire \add_90_I8_L14036_C104/carry[4]  ;
wire \add_90_I8_L14036_C104/carry[3]  ;
wire \add_90_I8_L14036_C104/carry[2]  ;
wire \add_90_I7_L14036_C104/carry[4]  ;
wire \add_90_I7_L14036_C104/carry[3]  ;
wire \add_90_I7_L14036_C104/carry[2]  ;
wire \add_90_I6_L14036_C104/carry[2]  ;
wire \add_90_I6_L14036_C104/carry[3]  ;
wire \add_90_I5_L14036_C104/carry[2]  ;
wire \add_90_I24_L14036_C103/carry[5]  ;
wire \add_90_I24_L14036_C103/carry[4]  ;
wire \add_90_I24_L14036_C103/carry[3]  ;
wire \add_90_I24_L14036_C103/carry[2]  ;
wire \add_90_I23_L14036_C103/carry[5]  ;
wire \add_90_I23_L14036_C103/carry[4]  ;
wire \add_90_I23_L14036_C103/carry[3]  ;
wire \add_90_I23_L14036_C103/carry[2]  ;
wire \add_90_I22_L14036_C103/carry[5]  ;
wire \add_90_I22_L14036_C103/carry[4]  ;
wire \add_90_I22_L14036_C103/carry[3]  ;
wire \add_90_I22_L14036_C103/carry[2]  ;
wire \add_90_I21_L14036_C103/carry[5]  ;
wire \add_90_I21_L14036_C103/carry[4]  ;
wire \add_90_I21_L14036_C103/carry[3]  ;
wire \add_90_I21_L14036_C103/carry[2]  ;
wire \add_90_I20_L14036_C103/carry[5]  ;
wire \add_90_I20_L14036_C103/carry[4]  ;
wire \add_90_I20_L14036_C103/carry[3]  ;
wire \add_90_I20_L14036_C103/carry[2]  ;
wire \add_90_I19_L14036_C103/carry[5]  ;
wire \add_90_I19_L14036_C103/carry[4]  ;
wire \add_90_I19_L14036_C103/carry[3]  ;
wire \add_90_I19_L14036_C103/carry[2]  ;
wire \add_90_I18_L14036_C103/carry[5]  ;
wire \add_90_I18_L14036_C103/carry[4]  ;
wire \add_90_I18_L14036_C103/carry[3]  ;
wire \add_90_I18_L14036_C103/carry[2]  ;
wire \add_90_I17_L14036_C103/carry[5]  ;
wire \add_90_I17_L14036_C103/carry[4]  ;
wire \add_90_I17_L14036_C103/carry[3]  ;
wire \add_90_I17_L14036_C103/carry[2]  ;
wire \add_90_I16_L14036_C103/carry[5]  ;
wire \add_90_I16_L14036_C103/carry[4]  ;
wire \add_90_I16_L14036_C103/carry[3]  ;
wire \add_90_I16_L14036_C103/carry[2]  ;
wire \add_90_I15_L14036_C103/carry[5]  ;
wire \add_90_I15_L14036_C103/carry[4]  ;
wire \add_90_I15_L14036_C103/carry[3]  ;
wire \add_90_I15_L14036_C103/carry[2]  ;
wire \add_90_I14_L14036_C103/carry[5]  ;
wire \add_90_I14_L14036_C103/carry[4]  ;
wire \add_90_I14_L14036_C103/carry[3]  ;
wire \add_90_I14_L14036_C103/carry[2]  ;
wire \add_90_I13_L14036_C103/carry[5]  ;
wire \add_90_I13_L14036_C103/carry[4]  ;
wire \add_90_I13_L14036_C103/carry[3]  ;
wire \add_90_I13_L14036_C103/carry[2]  ;
wire \add_90_I12_L14036_C103/carry[5]  ;
wire \add_90_I12_L14036_C103/carry[4]  ;
wire \add_90_I12_L14036_C103/carry[3]  ;
wire \add_90_I12_L14036_C103/carry[2]  ;
wire \add_90_I11_L14036_C103/carry[5]  ;
wire \add_90_I11_L14036_C103/carry[4]  ;
wire \add_90_I11_L14036_C103/carry[3]  ;
wire \add_90_I11_L14036_C103/carry[2]  ;
wire \add_90_I10_L14036_C103/carry[5]  ;
wire \add_90_I10_L14036_C103/carry[4]  ;
wire \add_90_I10_L14036_C103/carry[3]  ;
wire \add_90_I10_L14036_C103/carry[2]  ;
wire \add_90_I9_L14036_C103/carry[5]  ;
wire \add_90_I9_L14036_C103/carry[4]  ;
wire \add_90_I9_L14036_C103/carry[3]  ;
wire \add_90_I9_L14036_C103/carry[2]  ;
wire \add_90_I8_L14036_C103/carry[5]  ;
wire \add_90_I8_L14036_C103/carry[4]  ;
wire \add_90_I8_L14036_C103/carry[3]  ;
wire \add_90_I8_L14036_C103/carry[2]  ;
wire \add_90_I7_L14036_C103/carry[4]  ;
wire \add_90_I7_L14036_C103/carry[3]  ;
wire \add_90_I7_L14036_C103/carry[2]  ;
wire \add_90_I6_L14036_C103/carry[2]  ;
wire \add_90_I6_L14036_C103/carry[3]  ;
wire \add_90_I5_L14036_C103/carry[2]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n381 ;
wire n382 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n416 ;
wire n417 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire n429 ;
wire n430 ;
wire n431 ;
wire n432 ;
wire n433 ;
wire n434 ;
wire n435 ;
wire n436 ;
wire n437 ;
wire n438 ;
wire n439 ;
wire n440 ;
wire n441 ;
wire n442 ;
wire n443 ;
wire n444 ;
wire n445 ;
wire n446 ;
wire n447 ;
wire n448 ;
wire n449 ;
wire n450 ;
wire n451 ;
wire n452 ;
wire n453 ;
wire n454 ;
wire n455 ;
wire n456 ;
wire n457 ;
wire n458 ;
wire n459 ;
wire n460 ;
wire n461 ;
wire n462 ;
wire n463 ;
wire n464 ;
wire n465 ;
wire n466 ;
wire n467 ;
wire n468 ;
wire n469 ;
wire n470 ;
wire n471 ;
wire n472 ;
wire n473 ;
wire n474 ;
wire n475 ;
wire n476 ;
wire n477 ;
wire n478 ;
wire n479 ;
wire n480 ;
wire n481 ;
wire n482 ;
wire n483 ;
wire n484 ;
wire n485 ;
wire n486 ;
wire n487 ;
wire n488 ;
wire n489 ;
wire n490 ;
wire n491 ;
wire n492 ;
wire n493 ;
wire n494 ;
wire n495 ;
wire n496 ;
wire n497 ;
wire n498 ;
wire n499 ;
wire n500 ;
wire n501 ;
wire n502 ;
wire n503 ;
wire n504 ;
wire n505 ;
wire n506 ;
wire n507 ;
wire n508 ;
wire n509 ;
wire n510 ;
wire n511 ;
wire n512 ;
wire n513 ;
wire n514 ;
wire n515 ;
wire n516 ;
wire n517 ;
wire n518 ;
wire n519 ;
wire n520 ;
wire n521 ;
wire n522 ;
wire n523 ;
wire n524 ;
wire n525 ;
wire n526 ;
wire n527 ;
wire n528 ;
wire n529 ;
wire n530 ;
wire n531 ;
wire n532 ;
wire n533 ;
wire n534 ;
wire n535 ;
wire n536 ;
wire n537 ;
wire n538 ;
wire n539 ;
wire n540 ;
wire n541 ;
wire n542 ;
wire n543 ;
wire n544 ;
wire n545 ;
wire n546 ;
wire n547 ;
wire n548 ;
wire n549 ;
wire n550 ;
wire n551 ;
wire n552 ;
wire n553 ;
wire n554 ;
wire n555 ;
wire n556 ;
wire n557 ;
wire n558 ;
wire n559 ;
wire n560 ;
wire n561 ;
wire n562 ;
wire n563 ;
wire n564 ;
wire n565 ;
wire n566 ;
wire n567 ;
wire n568 ;
wire n569 ;
wire n570 ;
wire n571 ;
wire n572 ;
wire n573 ;
wire n574 ;
wire n575 ;
wire n576 ;
wire n577 ;
wire n578 ;
wire n579 ;
wire n580 ;
wire n581 ;
wire n582 ;
wire n583 ;
wire n584 ;
wire n585 ;
wire n586 ;
wire n587 ;
wire n588 ;
wire n589 ;
wire n590 ;
wire n591 ;
wire n592 ;
wire n593 ;
wire n594 ;
wire n595 ;
wire n596 ;
wire n597 ;
wire n598 ;
wire n599 ;
wire n600 ;
wire n601 ;
wire n602 ;
wire n603 ;
wire n604 ;
wire n605 ;
wire n606 ;
wire n607 ;
wire n608 ;
wire n609 ;
wire n610 ;
wire n611 ;
wire n612 ;
wire n613 ;
wire n614 ;
wire n615 ;
wire [9:0] s_exp_10_o ;
wire [5:0] s_dvd_zeros ;
wire [5:0] s_div_zeros ;
wire [9:0] s_expa_in ;
input p_desc1176_p_O_DFFX1 ;
input p_desc1177_p_O_DFFX1 ;
input p_desc1178_p_O_DFFX1 ;
input p_desc1179_p_O_DFFX1 ;
input p_desc1180_p_O_DFFX1 ;
input p_desc1181_p_O_DFFX1 ;
input p_desc1182_p_O_DFFX1 ;
input p_desc1183_p_O_DFFX1 ;
input p_desc1184_p_O_DFFX1 ;
input p_desc1185_p_O_DFFX1 ;
input p_desc1186_p_O_DFFX1 ;
input p_desc1187_p_O_DFFX1 ;
input p_desc1188_p_O_DFFX1 ;
input p_desc1189_p_O_DFFX1 ;
input p_desc1190_p_O_DFFX1 ;
input p_desc1191_p_O_DFFX1 ;
input p_desc1192_p_O_DFFX1 ;
input p_desc1193_p_O_DFFX1 ;
input p_desc1194_p_O_DFFX1 ;
input p_desc1195_p_O_DFFX1 ;
input p_desc1196_p_O_DFFX1 ;
input p_desc1197_p_O_DFFX1 ;
input p_desc1198_p_O_DFFX1 ;
input p_desc1199_p_O_DFFX1 ;
input p_desc1200_p_O_DFFX1 ;
input p_desc1201_p_O_DFFX1 ;
input p_desc1202_p_O_DFFX1 ;
input p_desc1203_p_O_DFFX1 ;
input p_desc1204_p_O_DFFX1 ;
input p_desc1205_p_O_DFFX1 ;
input p_desc1206_p_O_DFFX1 ;
input p_desc1207_p_O_DFFX1 ;
input p_desc1208_p_O_DFFX1 ;
input p_desc1209_p_O_DFFX1 ;
input p_desc1210_p_O_DFFX1 ;
input p_desc1211_p_O_DFFX1 ;
input p_desc1212_p_O_DFFX1 ;
input p_desc1213_p_O_DFFX1 ;
// instances
  p_O_DFFX1 desc1176(.D(N1534),.CLK(clk_i),.Q(s_expa_in[8:8]),.E(p_desc1176_p_O_DFFX1));
  p_O_DFFX1 desc1177(.D(N1533),.CLK(clk_i),.Q(s_expa_in[7:7]),.E(p_desc1177_p_O_DFFX1));
  p_O_DFFX1 desc1178(.D(N1532),.CLK(clk_i),.Q(s_expa_in[6:6]),.E(p_desc1178_p_O_DFFX1));
  p_O_DFFX1 desc1179(.D(N1531),.CLK(clk_i),.Q(s_expa_in[5:5]),.E(p_desc1179_p_O_DFFX1));
  p_O_DFFX1 desc1180(.D(N1530),.CLK(clk_i),.Q(s_expa_in[4:4]),.E(p_desc1180_p_O_DFFX1));
  p_O_DFFX1 desc1181(.D(N1529),.CLK(clk_i),.Q(s_expa_in[3:3]),.E(p_desc1181_p_O_DFFX1));
  p_O_DFFX1 desc1182(.D(N1528),.CLK(clk_i),.Q(s_expa_in[2:2]),.E(p_desc1182_p_O_DFFX1));
  p_O_DFFX1 desc1183(.D(N1527),.CLK(clk_i),.Q(s_expa_in[1:1]),.E(p_desc1183_p_O_DFFX1));
  p_O_DFFX1 desc1184(.D(N1526),.CLK(clk_i),.Q(s_expa_in[0:0]),.E(p_desc1184_p_O_DFFX1));
  p_O_DFFX1 desc1185(.D(N1543),.CLK(clk_i),.QN(n9),.E(p_desc1185_p_O_DFFX1));
  p_O_DFFX1 desc1186(.D(N1542),.CLK(clk_i),.Q(N1561),.QN(n1),.E(p_desc1186_p_O_DFFX1));
  p_O_DFFX1 desc1187(.D(N1541),.CLK(clk_i),.QN(n8),.E(p_desc1187_p_O_DFFX1));
  p_O_DFFX1 desc1188(.D(N1540),.CLK(clk_i),.QN(n7),.E(p_desc1188_p_O_DFFX1));
  p_O_DFFX1 desc1189(.D(N1539),.CLK(clk_i),.QN(n6),.E(p_desc1189_p_O_DFFX1));
  p_O_DFFX1 desc1190(.D(N1538),.CLK(clk_i),.QN(n5),.E(p_desc1190_p_O_DFFX1));
  p_O_DFFX1 desc1191(.D(N1537),.CLK(clk_i),.QN(n4),.E(p_desc1191_p_O_DFFX1));
  p_O_DFFX1 desc1192(.D(N1536),.CLK(clk_i),.QN(n2),.E(p_desc1192_p_O_DFFX1));
  p_O_DFFX1 desc1193(.D(N1535),.CLK(clk_i),.QN(n3),.E(p_desc1193_p_O_DFFX1));
  p_O_DFFX1 desc1194(.D(N1583),.CLK(clk_i),.Q(s_exp_10_o[9:9]),.E(p_desc1194_p_O_DFFX1));
  p_O_DFFX1 desc1195(.D(s_exp_10_o[9:9]),.CLK(clk_i),.Q(exp_10_o[9:9]),.E(p_desc1195_p_O_DFFX1));
  p_O_DFFX1 desc1196(.D(N1582),.CLK(clk_i),.Q(s_exp_10_o[8:8]),.E(p_desc1196_p_O_DFFX1));
  p_O_DFFX1 desc1197(.D(s_exp_10_o[8:8]),.CLK(clk_i),.Q(exp_10_o[8:8]),.E(p_desc1197_p_O_DFFX1));
  p_O_DFFX1 desc1198(.D(N1581),.CLK(clk_i),.Q(s_exp_10_o[7:7]),.E(p_desc1198_p_O_DFFX1));
  p_O_DFFX1 desc1199(.D(s_exp_10_o[7:7]),.CLK(clk_i),.Q(exp_10_o[7:7]),.E(p_desc1199_p_O_DFFX1));
  p_O_DFFX1 desc1200(.D(N1580),.CLK(clk_i),.Q(s_exp_10_o[6:6]),.E(p_desc1200_p_O_DFFX1));
  p_O_DFFX1 desc1201(.D(s_exp_10_o[6:6]),.CLK(clk_i),.Q(exp_10_o[6:6]),.E(p_desc1201_p_O_DFFX1));
  p_O_DFFX1 desc1202(.D(N1579),.CLK(clk_i),.Q(s_exp_10_o[5:5]),.E(p_desc1202_p_O_DFFX1));
  p_O_DFFX1 desc1203(.D(s_exp_10_o[5:5]),.CLK(clk_i),.Q(exp_10_o[5:5]),.E(p_desc1203_p_O_DFFX1));
  p_O_DFFX1 desc1204(.D(N1578),.CLK(clk_i),.Q(s_exp_10_o[4:4]),.E(p_desc1204_p_O_DFFX1));
  p_O_DFFX1 desc1205(.D(s_exp_10_o[4:4]),.CLK(clk_i),.Q(exp_10_o[4:4]),.E(p_desc1205_p_O_DFFX1));
  p_O_DFFX1 desc1206(.D(N1577),.CLK(clk_i),.Q(s_exp_10_o[3:3]),.E(p_desc1206_p_O_DFFX1));
  p_O_DFFX1 desc1207(.D(s_exp_10_o[3:3]),.CLK(clk_i),.Q(exp_10_o[3:3]),.E(p_desc1207_p_O_DFFX1));
  p_O_DFFX1 desc1208(.D(N1576),.CLK(clk_i),.Q(s_exp_10_o[2:2]),.E(p_desc1208_p_O_DFFX1));
  p_O_DFFX1 desc1209(.D(s_exp_10_o[2:2]),.CLK(clk_i),.Q(exp_10_o[2:2]),.E(p_desc1209_p_O_DFFX1));
  p_O_DFFX1 desc1210(.D(N1575),.CLK(clk_i),.Q(s_exp_10_o[1:1]),.E(p_desc1210_p_O_DFFX1));
  p_O_DFFX1 desc1211(.D(s_exp_10_o[1:1]),.CLK(clk_i),.Q(exp_10_o[1:1]),.E(p_desc1211_p_O_DFFX1));
  p_O_DFFX1 desc1212(.D(N1574),.CLK(clk_i),.Q(s_exp_10_o[0:0]),.E(p_desc1212_p_O_DFFX1));
  p_O_DFFX1 desc1213(.D(s_exp_10_o[0:0]),.CLK(clk_i),.Q(exp_10_o[0:0]),.E(p_desc1213_p_O_DFFX1));
  AO222X1 U207(.IN1(n157),.IN2(N298),.IN3(n158),.IN4(n10),.IN5(n159),.IN6(N315),.Q(n156));
  AO221X1 U208(.IN1(n160),.IN2(N366),.IN3(n111),.IN4(n161),.IN5(n162),.Q(n155));
  AO22X1 U209(.IN1(n163),.IN2(N349),.IN3(n164),.IN4(N332),.Q(n162));
  NAND3X0 U210(.IN1(n165),.IN2(n166),.IN3(n167),.QN(n161));
  OA222X1 U211(.IN1(n53),.IN2(n168),.IN3(n50),.IN4(n169),.IN5(n170),.IN6(n171),.Q(n167));
  AO222X1 U212(.IN1(n174),.IN2(N502),.IN3(n31),.IN4(N485),.IN5(n175),.IN6(N519),.Q(n173));
  AO222X1 U213(.IN1(N564),.IN2(n176),.IN3(n177),.IN4(N536),.IN5(n178),.IN6(N553),.Q(n172));
  AOI22X1 U214(.IN1(N383),.IN2(n40),.IN3(N400),.IN4(n179),.QN(n166));
  OA22X1 U215(.IN1(n52),.IN2(n180),.IN3(n51),.IN4(n181),.Q(n165));
  AO221X1 U216(.IN1(n159),.IN2(N314),.IN3(n47),.IN4(N263),.IN5(n184),.Q(n183));
  AO22X1 U217(.IN1(n157),.IN2(N297),.IN3(n158),.IN4(N280),.Q(n184));
  AO221X1 U218(.IN1(n160),.IN2(N365),.IN3(n111),.IN4(n185),.IN5(n186),.Q(n182));
  AO22X1 U219(.IN1(n163),.IN2(N348),.IN3(n164),.IN4(N331),.Q(n186));
  NAND3X0 U220(.IN1(n187),.IN2(n188),.IN3(n189),.QN(n185));
  OA222X1 U221(.IN1(n58),.IN2(n168),.IN3(n55),.IN4(n169),.IN5(n190),.IN6(n171),.Q(n189));
  AO222X1 U222(.IN1(n174),.IN2(N501),.IN3(n31),.IN4(N484),.IN5(n175),.IN6(N518),.Q(n192));
  AO222X1 U223(.IN1(N563),.IN2(n176),.IN3(n177),.IN4(N535),.IN5(n178),.IN6(N552),.Q(n191));
  AOI22X1 U224(.IN1(N382),.IN2(n40),.IN3(N399),.IN4(n179),.QN(n188));
  OA22X1 U225(.IN1(n57),.IN2(n180),.IN3(n56),.IN4(n181),.Q(n187));
  AO221X1 U226(.IN1(n159),.IN2(N313),.IN3(n47),.IN4(N262),.IN5(n195),.Q(n194));
  AO22X1 U227(.IN1(n157),.IN2(N296),.IN3(n158),.IN4(N279),.Q(n195));
  AO221X1 U228(.IN1(n160),.IN2(N364),.IN3(n111),.IN4(n196),.IN5(n197),.Q(n193));
  AO22X1 U229(.IN1(n163),.IN2(N347),.IN3(n164),.IN4(N330),.Q(n197));
  NAND3X0 U230(.IN1(n198),.IN2(n199),.IN3(n200),.QN(n196));
  OA222X1 U231(.IN1(n99),.IN2(n168),.IN3(n96),.IN4(n169),.IN5(n201),.IN6(n171),.Q(n200));
  AO222X1 U232(.IN1(n174),.IN2(N500),.IN3(n31),.IN4(N483),.IN5(n175),.IN6(N517),.Q(n203));
  AO222X1 U233(.IN1(N562),.IN2(n176),.IN3(n177),.IN4(N534),.IN5(n178),.IN6(N551),.Q(n202));
  AOI22X1 U234(.IN1(N381),.IN2(n40),.IN3(N398),.IN4(n179),.QN(n199));
  OA22X1 U235(.IN1(n98),.IN2(n180),.IN3(n97),.IN4(n181),.Q(n198));
  AO22X1 U236(.IN1(n95),.IN2(n204),.IN3(n205),.IN4(n206),.Q(s_dvd_zeros[2:2]));
  NAND4X0 U237(.IN1(n207),.IN2(n208),.IN3(n209),.IN4(n210),.QN(n204));
  AOI221X1 U238(.IN1(N261),.IN2(n47),.IN3(N312),.IN4(n159),.IN5(n211),.QN(n210));
  AO22X1 U239(.IN1(N278),.IN2(n158),.IN3(N295),.IN4(n157),.Q(n211));
  AOI22X1 U240(.IN1(N329),.IN2(n164),.IN3(N346),.IN4(n163),.QN(n209));
  AO21X1 U241(.IN1(n212),.IN2(n213),.IN3(n214),.Q(n207));
  OA221X1 U242(.IN1(n101),.IN2(n181),.IN3(n102),.IN4(n180),.IN5(n215),.Q(n213));
  AOI22X1 U243(.IN1(N380),.IN2(n40),.IN3(N397),.IN4(n179),.QN(n215));
  OA222X1 U244(.IN1(n103),.IN2(n168),.IN3(n100),.IN4(n169),.IN5(n216),.IN6(n171),.Q(n212));
  AO222X1 U245(.IN1(n174),.IN2(N499),.IN3(n31),.IN4(N482),.IN5(n175),.IN6(N516),.Q(n218));
  AO222X1 U246(.IN1(N561),.IN2(n176),.IN3(n177),.IN4(N533),.IN5(n178),.IN6(N550),.Q(n217));
  AO22X1 U247(.IN1(n95),.IN2(n219),.IN3(n220),.IN4(N230),.Q(s_dvd_zeros[1:1]));
  NAND4X0 U248(.IN1(n221),.IN2(n222),.IN3(n223),.IN4(n224),.QN(n219));
  AOI221X1 U249(.IN1(N260),.IN2(n47),.IN3(N311),.IN4(n159),.IN5(n225),.QN(n224));
  AO22X1 U250(.IN1(N277),.IN2(n158),.IN3(N294),.IN4(n157),.Q(n225));
  AOI22X1 U251(.IN1(N328),.IN2(n164),.IN3(N345),.IN4(n163),.QN(n223));
  AO21X1 U252(.IN1(n226),.IN2(n227),.IN3(n214),.Q(n221));
  OA221X1 U253(.IN1(n105),.IN2(n181),.IN3(n106),.IN4(n180),.IN5(n228),.Q(n227));
  AOI22X1 U254(.IN1(N379),.IN2(n40),.IN3(N396),.IN4(n179),.QN(n228));
  OA222X1 U255(.IN1(n107),.IN2(n168),.IN3(n104),.IN4(n169),.IN5(n229),.IN6(n171),.Q(n226));
  AO222X1 U256(.IN1(n174),.IN2(N498),.IN3(n31),.IN4(N481),.IN5(n175),.IN6(N515),.Q(n231));
  AO222X1 U257(.IN1(N560),.IN2(n176),.IN3(n177),.IN4(N532),.IN5(n178),.IN6(N549),.Q(n230));
  AO22X1 U258(.IN1(n232),.IN2(\add_116/B[0] ),.IN3(n95),.IN4(n233),.Q(s_dvd_zeros[0:0]));
  NAND4X0 U259(.IN1(n234),.IN2(n235),.IN3(n236),.IN4(n237),.QN(n233));
  AOI221X1 U260(.IN1(N259),.IN2(n47),.IN3(N310),.IN4(n159),.IN5(n238),.QN(n237));
  AO22X1 U261(.IN1(N276),.IN2(n158),.IN3(N293),.IN4(n157),.Q(n238));
  AOI22X1 U262(.IN1(N327),.IN2(n164),.IN3(N344),.IN4(n163),.QN(n236));
  AO21X1 U263(.IN1(n244),.IN2(n245),.IN3(n214),.Q(n234));
  OA221X1 U264(.IN1(N457),.IN2(n181),.IN3(N440),.IN4(n180),.IN5(n246),.Q(n245));
  AOI22X1 U265(.IN1(N378),.IN2(n40),.IN3(N395),.IN4(n179),.QN(n246));
  OR2X1 U266(.IN1(n248),.IN2(n249),.Q(n180));
  OA222X1 U267(.IN1(N423),.IN2(n168),.IN3(N474),.IN4(n169),.IN5(n251),.IN6(n171),.Q(n244));
  AO222X1 U268(.IN1(n174),.IN2(N497),.IN3(n31),.IN4(N480),.IN5(n175),.IN6(N514),.Q(n253));
  AND2X1 U269(.IN1(n254),.IN2(n32),.Q(n174));
  AO222X1 U270(.IN1(N559),.IN2(n176),.IN3(n177),.IN4(N531),.IN5(n178),.IN6(N548),.Q(n252));
  AND2X1 U271(.IN1(n255),.IN2(n256),.Q(n177));
  NOR3X0 U272(.IN1(n25),.IN2(opa_i[0:0]),.IN3(n256),.QN(n176));
  OAI21X1 U273(.IN1(n257),.IN2(n205),.IN3(n108),.QN(n232));
  AO222X1 U274(.IN1(n261),.IN2(N961),.IN3(n262),.IN4(n11),.IN5(n263),.IN6(N978),.Q(n260));
  AO221X1 U275(.IN1(n264),.IN2(N1029),.IN3(n379),.IN4(n265),.IN5(n266),.Q(n259));
  AO22X1 U276(.IN1(n267),.IN2(N1012),.IN3(n268),.IN4(N995),.Q(n266));
  NAND3X0 U277(.IN1(n269),.IN2(n270),.IN3(n271),.QN(n265));
  OA222X1 U278(.IN1(n63),.IN2(n272),.IN3(n60),.IN4(n273),.IN5(n274),.IN6(n275),.Q(n271));
  AO222X1 U279(.IN1(n278),.IN2(N1165),.IN3(n13),.IN4(N1148),.IN5(n279),.IN6(N1182),.Q(n277));
  AO222X1 U280(.IN1(N1227),.IN2(n280),.IN3(n281),.IN4(N1199),.IN5(n282),.IN6(N1216),.Q(n276));
  AOI22X1 U281(.IN1(N1046),.IN2(n14),.IN3(N1063),.IN4(n283),.QN(n270));
  OA22X1 U282(.IN1(n62),.IN2(n284),.IN3(n61),.IN4(n285),.Q(n269));
  AO221X1 U283(.IN1(n263),.IN2(N977),.IN3(n16),.IN4(N926),.IN5(n288),.Q(n287));
  AO22X1 U284(.IN1(n261),.IN2(N960),.IN3(n262),.IN4(N943),.Q(n288));
  AO221X1 U285(.IN1(n264),.IN2(N1028),.IN3(n379),.IN4(n289),.IN5(n290),.Q(n286));
  AO22X1 U286(.IN1(n267),.IN2(N1011),.IN3(n268),.IN4(N994),.Q(n290));
  NAND3X0 U287(.IN1(n291),.IN2(n292),.IN3(n293),.QN(n289));
  OA222X1 U288(.IN1(n68),.IN2(n272),.IN3(n65),.IN4(n273),.IN5(n294),.IN6(n275),.Q(n293));
  AO222X1 U289(.IN1(n278),.IN2(N1164),.IN3(n13),.IN4(N1147),.IN5(n279),.IN6(N1181),.Q(n296));
  AO222X1 U290(.IN1(N1226),.IN2(n280),.IN3(n281),.IN4(N1198),.IN5(n282),.IN6(N1215),.Q(n295));
  AOI22X1 U291(.IN1(N1045),.IN2(n14),.IN3(N1062),.IN4(n283),.QN(n292));
  OA22X1 U292(.IN1(n67),.IN2(n284),.IN3(n66),.IN4(n285),.Q(n291));
  AO221X1 U293(.IN1(n263),.IN2(N976),.IN3(n16),.IN4(N925),.IN5(n299),.Q(n298));
  AO22X1 U294(.IN1(n261),.IN2(N959),.IN3(n262),.IN4(N942),.Q(n299));
  AO221X1 U295(.IN1(n264),.IN2(N1027),.IN3(n379),.IN4(n300),.IN5(n301),.Q(n297));
  AO22X1 U296(.IN1(n267),.IN2(N1010),.IN3(n268),.IN4(N993),.Q(n301));
  NAND3X0 U297(.IN1(n302),.IN2(n303),.IN3(n304),.QN(n300));
  OA222X1 U298(.IN1(n149),.IN2(n272),.IN3(n146),.IN4(n273),.IN5(n305),.IN6(n275),.Q(n304));
  AO222X1 U299(.IN1(n278),.IN2(N1163),.IN3(n13),.IN4(N1146),.IN5(n279),.IN6(N1180),.Q(n307));
  AO222X1 U300(.IN1(N1225),.IN2(n280),.IN3(n281),.IN4(N1197),.IN5(n282),.IN6(N1214),.Q(n306));
  AOI22X1 U301(.IN1(N1044),.IN2(n14),.IN3(N1061),.IN4(n283),.QN(n303));
  OA22X1 U302(.IN1(n148),.IN2(n284),.IN3(n147),.IN4(n285),.Q(n302));
  AO22X1 U303(.IN1(n145),.IN2(n308),.IN3(n309),.IN4(n310),.Q(s_div_zeros[2:2]));
  NAND4X0 U304(.IN1(n311),.IN2(n312),.IN3(n313),.IN4(n314),.QN(n308));
  AOI221X1 U305(.IN1(N924),.IN2(n16),.IN3(N975),.IN4(n263),.IN5(n315),.QN(n314));
  AO22X1 U306(.IN1(N941),.IN2(n262),.IN3(N958),.IN4(n261),.Q(n315));
  AOI22X1 U307(.IN1(N992),.IN2(n268),.IN3(N1009),.IN4(n267),.QN(n313));
  AO21X1 U308(.IN1(n316),.IN2(n317),.IN3(n318),.Q(n311));
  OA221X1 U309(.IN1(n151),.IN2(n285),.IN3(n152),.IN4(n284),.IN5(n319),.Q(n317));
  AOI22X1 U310(.IN1(N1043),.IN2(n14),.IN3(N1060),.IN4(n283),.QN(n319));
  OA222X1 U311(.IN1(n153),.IN2(n272),.IN3(n150),.IN4(n273),.IN5(n320),.IN6(n275),.Q(n316));
  AO222X1 U312(.IN1(n278),.IN2(N1162),.IN3(n13),.IN4(N1145),.IN5(n279),.IN6(N1179),.Q(n322));
  AO222X1 U313(.IN1(N1224),.IN2(n280),.IN3(n281),.IN4(N1196),.IN5(n282),.IN6(N1213),.Q(n321));
  AO22X1 U314(.IN1(n145),.IN2(n323),.IN3(n324),.IN4(N893),.Q(s_div_zeros[1:1]));
  NAND4X0 U315(.IN1(n325),.IN2(n326),.IN3(n327),.IN4(n328),.QN(n323));
  AOI221X1 U316(.IN1(N923),.IN2(n16),.IN3(N974),.IN4(n263),.IN5(n329),.QN(n328));
  AO22X1 U317(.IN1(N940),.IN2(n262),.IN3(N957),.IN4(n261),.Q(n329));
  AOI22X1 U318(.IN1(N991),.IN2(n268),.IN3(N1008),.IN4(n267),.QN(n327));
  AO21X1 U319(.IN1(n330),.IN2(n331),.IN3(n318),.Q(n325));
  OA221X1 U320(.IN1(n373),.IN2(n285),.IN3(n374),.IN4(n284),.IN5(n332),.Q(n331));
  AOI22X1 U321(.IN1(N1042),.IN2(n14),.IN3(N1059),.IN4(n283),.QN(n332));
  OA222X1 U322(.IN1(n375),.IN2(n272),.IN3(n154),.IN4(n273),.IN5(n333),.IN6(n275),.Q(n330));
  AO222X1 U323(.IN1(n278),.IN2(N1161),.IN3(n13),.IN4(N1144),.IN5(n279),.IN6(N1178),.Q(n335));
  AO222X1 U324(.IN1(N1223),.IN2(n280),.IN3(n281),.IN4(N1195),.IN5(n282),.IN6(N1212),.Q(n334));
  AO22X1 U325(.IN1(n336),.IN2(\add_117/B[0] ),.IN3(n145),.IN4(n337),.Q(s_div_zeros[0:0]));
  NAND4X0 U326(.IN1(n338),.IN2(n339),.IN3(n340),.IN4(n341),.QN(n337));
  AOI221X1 U327(.IN1(N922),.IN2(n16),.IN3(N973),.IN4(n263),.IN5(n342),.QN(n341));
  AO22X1 U328(.IN1(N939),.IN2(n262),.IN3(N956),.IN4(n261),.Q(n342));
  AOI22X1 U329(.IN1(N990),.IN2(n268),.IN3(N1007),.IN4(n267),.QN(n340));
  AO21X1 U330(.IN1(n348),.IN2(n349),.IN3(n318),.Q(n338));
  OA221X1 U331(.IN1(N1120),.IN2(n285),.IN3(N1103),.IN4(n284),.IN5(n350),.Q(n349));
  AOI22X1 U332(.IN1(N1041),.IN2(n14),.IN3(N1058),.IN4(n283),.QN(n350));
  OR2X1 U333(.IN1(n352),.IN2(n353),.Q(n284));
  OA222X1 U334(.IN1(N1086),.IN2(n272),.IN3(N1137),.IN4(n273),.IN5(n355),.IN6(n275),.Q(n348));
  AO222X1 U335(.IN1(n278),.IN2(N1160),.IN3(n13),.IN4(N1143),.IN5(n279),.IN6(N1177),.Q(n357));
  AND2X1 U336(.IN1(n358),.IN2(n399),.Q(n278));
  AO222X1 U337(.IN1(N1222),.IN2(n280),.IN3(n281),.IN4(N1194),.IN5(n282),.IN6(N1211),.Q(n356));
  AND2X1 U338(.IN1(n359),.IN2(n360),.Q(n281));
  NOR3X0 U339(.IN1(opb_i[1:1]),.IN2(opb_i[0:0]),.IN3(n360),.QN(n280));
  OAI21X1 U340(.IN1(n361),.IN2(n309),.IN3(n376),.QN(n336));
  AO22X1 U341(.IN1(N547),.IN2(n26),.IN3(n25),.IN4(N536),.Q(N553));
  AO22X1 U342(.IN1(N546),.IN2(n26),.IN3(n25),.IN4(N535),.Q(N552));
  AO22X1 U343(.IN1(N545),.IN2(n26),.IN3(n25),.IN4(N534),.Q(N551));
  AO22X1 U344(.IN1(N544),.IN2(n26),.IN3(n25),.IN4(N533),.Q(N550));
  AO22X1 U345(.IN1(N543),.IN2(n26),.IN3(n25),.IN4(N532),.Q(N549));
  AO22X1 U346(.IN1(N542),.IN2(n26),.IN3(n25),.IN4(N531),.Q(N548));
  AO22X1 U347(.IN1(N530),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N519),.Q(N536));
  AO22X1 U348(.IN1(N529),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N518),.Q(N535));
  AO22X1 U349(.IN1(N528),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N517),.Q(N534));
  AO22X1 U350(.IN1(N527),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N516),.Q(N533));
  AO22X1 U351(.IN1(N526),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N515),.Q(N532));
  AO22X1 U352(.IN1(N525),.IN2(n27),.IN3(opa_i[2:2]),.IN4(N514),.Q(N531));
  AO22X1 U353(.IN1(N513),.IN2(n29),.IN3(n28),.IN4(N502),.Q(N519));
  AO22X1 U354(.IN1(N512),.IN2(n29),.IN3(n28),.IN4(N501),.Q(N518));
  AO22X1 U355(.IN1(N511),.IN2(n29),.IN3(n28),.IN4(N500),.Q(N517));
  AO22X1 U356(.IN1(N510),.IN2(n29),.IN3(n28),.IN4(N499),.Q(N516));
  AO22X1 U357(.IN1(N509),.IN2(n29),.IN3(n28),.IN4(N498),.Q(N515));
  AO22X1 U358(.IN1(N508),.IN2(n29),.IN3(n28),.IN4(N497),.Q(N514));
  AO22X1 U359(.IN1(N496),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N485),.Q(N502));
  AO22X1 U360(.IN1(N495),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N484),.Q(N501));
  AO22X1 U361(.IN1(N494),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N483),.Q(N500));
  AO22X1 U362(.IN1(N493),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N482),.Q(N499));
  AO22X1 U363(.IN1(N492),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N481),.Q(N498));
  AO22X1 U364(.IN1(N491),.IN2(n30),.IN3(opa_i[4:4]),.IN4(N480),.Q(N497));
  AO22X1 U365(.IN1(N479),.IN2(n32),.IN3(n31),.IN4(N468),.Q(N485));
  AO22X1 U366(.IN1(N478),.IN2(n32),.IN3(n31),.IN4(N467),.Q(N484));
  AO22X1 U367(.IN1(N477),.IN2(n32),.IN3(n31),.IN4(N466),.Q(N483));
  AO22X1 U368(.IN1(N476),.IN2(n32),.IN3(n31),.IN4(N465),.Q(N482));
  AO22X1 U369(.IN1(N475),.IN2(n32),.IN3(n31),.IN4(N464),.Q(N481));
  AO22X1 U370(.IN1(N474),.IN2(n32),.IN3(n31),.IN4(N463),.Q(N480));
  AO22X1 U371(.IN1(N462),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N451),.Q(N468));
  AO22X1 U372(.IN1(N461),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N450),.Q(N467));
  AO22X1 U373(.IN1(N460),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N449),.Q(N466));
  AO22X1 U374(.IN1(N459),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N448),.Q(N465));
  AO22X1 U375(.IN1(N458),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N447),.Q(N464));
  AO22X1 U376(.IN1(N457),.IN2(n33),.IN3(opa_i[6:6]),.IN4(N446),.Q(N463));
  AO22X1 U377(.IN1(N445),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N434),.Q(N451));
  AO22X1 U378(.IN1(N444),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N433),.Q(N450));
  AO22X1 U379(.IN1(N443),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N432),.Q(N449));
  AO22X1 U380(.IN1(N442),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N431),.Q(N448));
  AO22X1 U381(.IN1(N441),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N430),.Q(N447));
  AO22X1 U382(.IN1(N440),.IN2(n34),.IN3(opa_i[7:7]),.IN4(N429),.Q(N446));
  AO22X1 U383(.IN1(N428),.IN2(n36),.IN3(n35),.IN4(N417),.Q(N434));
  AO22X1 U384(.IN1(N427),.IN2(n36),.IN3(n35),.IN4(N416),.Q(N433));
  AO22X1 U385(.IN1(N426),.IN2(n36),.IN3(n35),.IN4(N415),.Q(N432));
  AO22X1 U386(.IN1(N425),.IN2(n36),.IN3(n35),.IN4(N414),.Q(N431));
  AO22X1 U387(.IN1(N424),.IN2(n36),.IN3(n35),.IN4(N413),.Q(N430));
  AO22X1 U388(.IN1(N423),.IN2(n36),.IN3(n35),.IN4(N412),.Q(N429));
  AO22X1 U389(.IN1(N411),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N400),.Q(N417));
  AO22X1 U390(.IN1(N410),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N399),.Q(N416));
  AO22X1 U391(.IN1(N409),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N398),.Q(N415));
  AO22X1 U392(.IN1(N408),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N397),.Q(N414));
  AO22X1 U393(.IN1(N407),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N396),.Q(N413));
  AO22X1 U394(.IN1(N406),.IN2(n37),.IN3(opa_i[9:9]),.IN4(N395),.Q(N412));
  AO22X1 U395(.IN1(N394),.IN2(n39),.IN3(n38),.IN4(N383),.Q(N400));
  AO22X1 U396(.IN1(N393),.IN2(n39),.IN3(n38),.IN4(N382),.Q(N399));
  AO22X1 U397(.IN1(N392),.IN2(n39),.IN3(n38),.IN4(N381),.Q(N398));
  AO22X1 U398(.IN1(N391),.IN2(n39),.IN3(n38),.IN4(N380),.Q(N397));
  AO22X1 U399(.IN1(N390),.IN2(n39),.IN3(n38),.IN4(N379),.Q(N396));
  AO22X1 U400(.IN1(N389),.IN2(n39),.IN3(n38),.IN4(N378),.Q(N395));
  AO22X1 U401(.IN1(N377),.IN2(n41),.IN3(n40),.IN4(N366),.Q(N383));
  AO22X1 U402(.IN1(N376),.IN2(n41),.IN3(n40),.IN4(N365),.Q(N382));
  AO22X1 U403(.IN1(N375),.IN2(n41),.IN3(n40),.IN4(N364),.Q(N381));
  AO22X1 U404(.IN1(N374),.IN2(n41),.IN3(n40),.IN4(N363),.Q(N380));
  AO22X1 U405(.IN1(N373),.IN2(n41),.IN3(n40),.IN4(N362),.Q(N379));
  AO22X1 U406(.IN1(N372),.IN2(n41),.IN3(n40),.IN4(N361),.Q(N378));
  AO22X1 U407(.IN1(N360),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N349),.Q(N366));
  AO22X1 U408(.IN1(N359),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N348),.Q(N365));
  AO22X1 U409(.IN1(N358),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N347),.Q(N364));
  AO22X1 U410(.IN1(N357),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N346),.Q(N363));
  AO22X1 U411(.IN1(N356),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N345),.Q(N362));
  AO22X1 U412(.IN1(N355),.IN2(n117),.IN3(opa_i[12:12]),.IN4(N344),.Q(N361));
  AO22X1 U413(.IN1(N343),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N332),.Q(N349));
  AO22X1 U414(.IN1(N342),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N331),.Q(N348));
  AO22X1 U415(.IN1(N341),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N330),.Q(N347));
  AO22X1 U416(.IN1(N340),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N329),.Q(N346));
  AO22X1 U417(.IN1(N339),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N328),.Q(N345));
  AO22X1 U418(.IN1(N338),.IN2(n42),.IN3(opa_i[13:13]),.IN4(N327),.Q(N344));
  AO22X1 U419(.IN1(N326),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N315),.Q(N332));
  AO22X1 U420(.IN1(N325),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N314),.Q(N331));
  AO22X1 U421(.IN1(N324),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N313),.Q(N330));
  AO22X1 U422(.IN1(N323),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N312),.Q(N329));
  AO22X1 U423(.IN1(N322),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N311),.Q(N328));
  AO22X1 U424(.IN1(N321),.IN2(n43),.IN3(opa_i[14:14]),.IN4(N310),.Q(N327));
  AO22X1 U425(.IN1(N309),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N298),.Q(N315));
  AO22X1 U426(.IN1(N308),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N297),.Q(N314));
  AO22X1 U427(.IN1(N307),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N296),.Q(N313));
  AO22X1 U428(.IN1(N306),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N295),.Q(N312));
  AO22X1 U429(.IN1(N305),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N294),.Q(N311));
  AO22X1 U430(.IN1(N304),.IN2(n44),.IN3(opa_i[15:15]),.IN4(N293),.Q(N310));
  AO22X1 U431(.IN1(N292),.IN2(n45),.IN3(opa_i[16:16]),.IN4(n10),.Q(N298));
  AO22X1 U432(.IN1(N291),.IN2(n45),.IN3(opa_i[16:16]),.IN4(N280),.Q(N297));
  AO22X1 U433(.IN1(N290),.IN2(n45),.IN3(opa_i[16:16]),.IN4(N279),.Q(N296));
  AO22X1 U434(.IN1(N289),.IN2(n45),.IN3(opa_i[16:16]),.IN4(N278),.Q(N295));
  AO22X1 U435(.IN1(N288),.IN2(n45),.IN3(opa_i[16:16]),.IN4(N277),.Q(N294));
  AO22X1 U436(.IN1(N287),.IN2(n45),.IN3(opa_i[16:16]),.IN4(N276),.Q(N293));
  AO22X1 U438(.IN1(N274),.IN2(n46),.IN3(opa_i[17:17]),.IN4(N263),.Q(N280));
  AO22X1 U439(.IN1(N273),.IN2(n46),.IN3(opa_i[17:17]),.IN4(N262),.Q(N279));
  AO22X1 U440(.IN1(N272),.IN2(n46),.IN3(opa_i[17:17]),.IN4(N261),.Q(N278));
  AO22X1 U441(.IN1(N271),.IN2(n46),.IN3(opa_i[17:17]),.IN4(N260),.Q(N277));
  AO22X1 U442(.IN1(N270),.IN2(n46),.IN3(opa_i[17:17]),.IN4(N259),.Q(N276));
  AO22X1 U445(.IN1(N256),.IN2(n48),.IN3(N246),.IN4(n47),.Q(N262));
  AO22X1 U446(.IN1(N255),.IN2(n48),.IN3(n47),.IN4(N245),.Q(N261));
  AO22X1 U447(.IN1(N254),.IN2(n48),.IN3(n47),.IN4(N244),.Q(N260));
  AO22X1 U448(.IN1(N253),.IN2(n48),.IN3(n47),.IN4(N243),.Q(N259));
  AND2X1 U450(.IN1(N241),.IN2(n110),.Q(N246));
  AO22X1 U451(.IN1(N240),.IN2(n110),.IN3(opa_i[19:19]),.IN4(N231),.Q(N245));
  AO22X1 U452(.IN1(N239),.IN2(n110),.IN3(opa_i[19:19]),.IN4(N230),.Q(N244));
  AO22X1 U453(.IN1(N238),.IN2(n110),.IN3(N229),.IN4(opa_i[19:19]),.Q(N243));
  AND2X1 U455(.IN1(n363),.IN2(n364),.Q(N231));
  XOR2X1 U456(.IN1(n364),.IN2(n363),.Q(N230));
  AO21X1 U457(.IN1(n258),.IN2(n109),.IN3(n220),.Q(n364));
  XOR2X1 U458(.IN1(n365),.IN2(opa_i[20:20]),.Q(N229));
  XOR2X1 U459(.IN1(n258),.IN2(opa_i[21:21]),.Q(n365));
  XOR2X1 U460(.IN1(N192),.IN2(opa_i[22:22]),.Q(n258));
  NOR4X0 U461(.IN1(opa_i[30:30]),.IN2(opa_i[29:29]),.IN3(opa_i[28:28]),.IN4(opa_i[27:27]),.QN(n367));
  NOR4X0 U462(.IN1(opa_i[26:26]),.IN2(opa_i[25:25]),.IN3(opa_i[24:24]),.IN4(opa_i[23:23]),.QN(n366));
  AO22X1 U463(.IN1(N1210),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1199),.Q(N1216));
  AO22X1 U464(.IN1(N1209),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1198),.Q(N1215));
  AO22X1 U465(.IN1(N1208),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1197),.Q(N1214));
  AO22X1 U466(.IN1(N1207),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1196),.Q(N1213));
  AO22X1 U467(.IN1(N1206),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1195),.Q(N1212));
  AO22X1 U468(.IN1(N1205),.IN2(n403),.IN3(opb_i[1:1]),.IN4(N1194),.Q(N1211));
  AO22X1 U469(.IN1(N1193),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1182),.Q(N1199));
  AO22X1 U470(.IN1(N1192),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1181),.Q(N1198));
  AO22X1 U471(.IN1(N1191),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1180),.Q(N1197));
  AO22X1 U472(.IN1(N1190),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1179),.Q(N1196));
  AO22X1 U473(.IN1(N1189),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1178),.Q(N1195));
  AO22X1 U474(.IN1(N1188),.IN2(n402),.IN3(opb_i[2:2]),.IN4(N1177),.Q(N1194));
  AO22X1 U475(.IN1(N1176),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1165),.Q(N1182));
  AO22X1 U476(.IN1(N1175),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1164),.Q(N1181));
  AO22X1 U477(.IN1(N1174),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1163),.Q(N1180));
  AO22X1 U478(.IN1(N1173),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1162),.Q(N1179));
  AO22X1 U479(.IN1(N1172),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1161),.Q(N1178));
  AO22X1 U480(.IN1(N1171),.IN2(n401),.IN3(opb_i[3:3]),.IN4(N1160),.Q(N1177));
  AO22X1 U481(.IN1(N1159),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1148),.Q(N1165));
  AO22X1 U482(.IN1(N1158),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1147),.Q(N1164));
  AO22X1 U483(.IN1(N1157),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1146),.Q(N1163));
  AO22X1 U484(.IN1(N1156),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1145),.Q(N1162));
  AO22X1 U485(.IN1(N1155),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1144),.Q(N1161));
  AO22X1 U486(.IN1(N1154),.IN2(n400),.IN3(opb_i[4:4]),.IN4(N1143),.Q(N1160));
  AO22X1 U487(.IN1(N1142),.IN2(n399),.IN3(n13),.IN4(N1131),.Q(N1148));
  AO22X1 U488(.IN1(N1141),.IN2(n399),.IN3(n13),.IN4(N1130),.Q(N1147));
  AO22X1 U489(.IN1(N1140),.IN2(n399),.IN3(n13),.IN4(N1129),.Q(N1146));
  AO22X1 U490(.IN1(N1139),.IN2(n399),.IN3(n13),.IN4(N1128),.Q(N1145));
  AO22X1 U491(.IN1(N1138),.IN2(n399),.IN3(n13),.IN4(N1127),.Q(N1144));
  AO22X1 U492(.IN1(N1137),.IN2(n399),.IN3(n13),.IN4(N1126),.Q(N1143));
  AO22X1 U493(.IN1(N1125),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1114),.Q(N1131));
  AO22X1 U494(.IN1(N1124),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1113),.Q(N1130));
  AO22X1 U495(.IN1(N1123),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1112),.Q(N1129));
  AO22X1 U496(.IN1(N1122),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1111),.Q(N1128));
  AO22X1 U497(.IN1(N1121),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1110),.Q(N1127));
  AO22X1 U498(.IN1(N1120),.IN2(n398),.IN3(opb_i[6:6]),.IN4(N1109),.Q(N1126));
  AO22X1 U499(.IN1(N1108),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1097),.Q(N1114));
  AO22X1 U500(.IN1(N1107),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1096),.Q(N1113));
  AO22X1 U501(.IN1(N1106),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1095),.Q(N1112));
  AO22X1 U502(.IN1(N1105),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1094),.Q(N1111));
  AO22X1 U503(.IN1(N1104),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1093),.Q(N1110));
  AO22X1 U504(.IN1(N1103),.IN2(n397),.IN3(opb_i[7:7]),.IN4(N1092),.Q(N1109));
  AO22X1 U505(.IN1(N1091),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1080),.Q(N1097));
  AO22X1 U506(.IN1(N1090),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1079),.Q(N1096));
  AO22X1 U507(.IN1(N1089),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1078),.Q(N1095));
  AO22X1 U508(.IN1(N1088),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1077),.Q(N1094));
  AO22X1 U509(.IN1(N1087),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1076),.Q(N1093));
  AO22X1 U510(.IN1(N1086),.IN2(n396),.IN3(opb_i[8:8]),.IN4(N1075),.Q(N1092));
  AO22X1 U511(.IN1(N1074),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1063),.Q(N1080));
  AO22X1 U512(.IN1(N1073),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1062),.Q(N1079));
  AO22X1 U513(.IN1(N1072),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1061),.Q(N1078));
  AO22X1 U514(.IN1(N1071),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1060),.Q(N1077));
  AO22X1 U515(.IN1(N1070),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1059),.Q(N1076));
  AO22X1 U516(.IN1(N1069),.IN2(n395),.IN3(opb_i[9:9]),.IN4(N1058),.Q(N1075));
  AO22X1 U517(.IN1(N1057),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1046),.Q(N1063));
  AO22X1 U518(.IN1(N1056),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1045),.Q(N1062));
  AO22X1 U519(.IN1(N1055),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1044),.Q(N1061));
  AO22X1 U520(.IN1(N1054),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1043),.Q(N1060));
  AO22X1 U521(.IN1(N1053),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1042),.Q(N1059));
  AO22X1 U522(.IN1(N1052),.IN2(n394),.IN3(opb_i[10:10]),.IN4(N1041),.Q(N1058));
  AO22X1 U523(.IN1(N1040),.IN2(n392),.IN3(n14),.IN4(N1029),.Q(N1046));
  AO22X1 U524(.IN1(N1039),.IN2(n392),.IN3(n14),.IN4(N1028),.Q(N1045));
  AO22X1 U525(.IN1(N1038),.IN2(n392),.IN3(n14),.IN4(N1027),.Q(N1044));
  AO22X1 U526(.IN1(N1037),.IN2(n392),.IN3(n14),.IN4(N1026),.Q(N1043));
  AO22X1 U527(.IN1(N1036),.IN2(n392),.IN3(n14),.IN4(N1025),.Q(N1042));
  AO22X1 U528(.IN1(N1035),.IN2(n392),.IN3(n14),.IN4(N1024),.Q(N1041));
  AO22X1 U529(.IN1(N1023),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1012),.Q(N1029));
  AO22X1 U530(.IN1(N1022),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1011),.Q(N1028));
  AO22X1 U531(.IN1(N1021),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1010),.Q(N1027));
  AO22X1 U532(.IN1(N1020),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1009),.Q(N1026));
  AO22X1 U533(.IN1(N1019),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1008),.Q(N1025));
  AO22X1 U534(.IN1(N1018),.IN2(n391),.IN3(opb_i[12:12]),.IN4(N1007),.Q(N1024));
  AO22X1 U535(.IN1(N1006),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N995),.Q(N1012));
  AO22X1 U536(.IN1(N989),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N978),.Q(N995));
  AO22X1 U537(.IN1(N972),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N961),.Q(N978));
  AO22X1 U538(.IN1(N955),.IN2(n387),.IN3(opb_i[16:16]),.IN4(n11),.Q(N961));
  AO22X1 U541(.IN1(N1005),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N994),.Q(N1011));
  AO22X1 U542(.IN1(N988),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N977),.Q(N994));
  AO22X1 U543(.IN1(N971),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N960),.Q(N977));
  AO22X1 U544(.IN1(N954),.IN2(n387),.IN3(opb_i[16:16]),.IN4(N943),.Q(N960));
  AO22X1 U545(.IN1(N937),.IN2(n386),.IN3(opb_i[17:17]),.IN4(N926),.Q(N943));
  AO22X1 U548(.IN1(N1004),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N993),.Q(N1010));
  AO22X1 U549(.IN1(N987),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N976),.Q(N993));
  AO22X1 U550(.IN1(N970),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N959),.Q(N976));
  AO22X1 U551(.IN1(N953),.IN2(n387),.IN3(opb_i[16:16]),.IN4(N942),.Q(N959));
  AO22X1 U552(.IN1(N936),.IN2(n386),.IN3(opb_i[17:17]),.IN4(N925),.Q(N942));
  AO22X1 U553(.IN1(N919),.IN2(n385),.IN3(N909),.IN4(n16),.Q(N925));
  AND2X1 U554(.IN1(N904),.IN2(n378),.Q(N909));
  AO22X1 U555(.IN1(N1003),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N992),.Q(N1009));
  AO22X1 U556(.IN1(N986),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N975),.Q(N992));
  AO22X1 U557(.IN1(N969),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N958),.Q(N975));
  AO22X1 U558(.IN1(N952),.IN2(n387),.IN3(opb_i[16:16]),.IN4(N941),.Q(N958));
  AO22X1 U559(.IN1(N935),.IN2(n386),.IN3(opb_i[17:17]),.IN4(N924),.Q(N941));
  AO22X1 U560(.IN1(N918),.IN2(n385),.IN3(n16),.IN4(N908),.Q(N924));
  AO22X1 U561(.IN1(N903),.IN2(n378),.IN3(opb_i[19:19]),.IN4(N894),.Q(N908));
  AND2X1 U562(.IN1(n368),.IN2(n369),.Q(N894));
  AO22X1 U563(.IN1(N1002),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N991),.Q(N1008));
  AO22X1 U564(.IN1(N985),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N974),.Q(N991));
  AO22X1 U565(.IN1(N968),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N957),.Q(N974));
  AO22X1 U566(.IN1(N951),.IN2(n387),.IN3(opb_i[16:16]),.IN4(N940),.Q(N957));
  AO22X1 U567(.IN1(N934),.IN2(n386),.IN3(opb_i[17:17]),.IN4(N923),.Q(N940));
  AO22X1 U568(.IN1(N917),.IN2(n385),.IN3(n16),.IN4(N907),.Q(N923));
  AO22X1 U569(.IN1(N902),.IN2(n378),.IN3(opb_i[19:19]),.IN4(N893),.Q(N907));
  XOR2X1 U570(.IN1(n369),.IN2(n368),.Q(N893));
  AO21X1 U571(.IN1(n362),.IN2(n377),.IN3(n324),.Q(n369));
  AO22X1 U572(.IN1(N1001),.IN2(n390),.IN3(opb_i[13:13]),.IN4(N990),.Q(N1007));
  AO22X1 U573(.IN1(N984),.IN2(n389),.IN3(opb_i[14:14]),.IN4(N973),.Q(N990));
  AO22X1 U574(.IN1(N967),.IN2(n388),.IN3(opb_i[15:15]),.IN4(N956),.Q(N973));
  AO22X1 U575(.IN1(N950),.IN2(n387),.IN3(opb_i[16:16]),.IN4(N939),.Q(N956));
  AO22X1 U576(.IN1(N933),.IN2(n386),.IN3(opb_i[17:17]),.IN4(N922),.Q(N939));
  AO22X1 U577(.IN1(N916),.IN2(n385),.IN3(n16),.IN4(N906),.Q(N922));
  AO22X1 U578(.IN1(N901),.IN2(n378),.IN3(N892),.IN4(opb_i[19:19]),.Q(N906));
  XOR2X1 U579(.IN1(n370),.IN2(opb_i[20:20]),.Q(N892));
  XOR2X1 U580(.IN1(n362),.IN2(opb_i[21:21]),.Q(n370));
  XOR2X1 U581(.IN1(N199),.IN2(opb_i[22:22]),.Q(n362));
  NOR4X0 U582(.IN1(opb_i[30:30]),.IN2(opb_i[29:29]),.IN3(opb_i[28:28]),.IN4(opb_i[27:27]),.QN(n372));
  NOR4X0 U583(.IN1(opb_i[26:26]),.IN2(opb_i[25:25]),.IN3(opb_i[24:24]),.IN4(opb_i[23:23]),.QN(n371));
  pre_norm_div_DW01_add_3_inj add_2_root_sub_0_root_add_118_2(.A({1'b0,s_expa_in[8:0]}),.B({n12,N1562,N1561,n8,n7,n6,n5,n4,n2,n3}),.CI(1'b0),.SUM({N1553,N1552,N1551,N1550,N1549,N1548,N1547,N1546,N1545,N1544}));
  pre_norm_div_DW01_add_2_inj add_1_root_sub_0_root_add_118_2(.A({N1553,N1552,N1551,N1550,N1549,N1548,N1547,N1546,N1545,N1544}),.B({1'b0,1'b0,1'b0,1'b0,n18,s_div_zeros[4:0]}),.CI(1'b0),.SUM({N1573,N1572,N1571,N1570,N1569,N1568,N1567,N1566,N1565,N1564}));
  pre_norm_div_DW01_sub_0_inj sub_0_root_sub_0_root_add_118_2(.A({N1573,N1572,N1571,N1570,N1569,N1568,N1567,N1566,N1565,N1564}),.B({1'b0,1'b0,1'b0,1'b0,n20,s_dvd_zeros[4:0]}),.CI(1'b0),.DIFF({N1583,N1582,N1581,N1580,N1579,N1578,N1577,N1576,N1575,N1574}));
  HADDX1 desc1214(.A0(N1212),.B0(N1211),.C1(\add_90_I24_L14036_C104/carry[2] ),.SO(N1223));
  HADDX1 desc1215(.A0(N1213),.B0(\add_90_I24_L14036_C104/carry[2] ),.C1(\add_90_I24_L14036_C104/carry[3] ),.SO(N1224));
  HADDX1 desc1216(.A0(N1214),.B0(\add_90_I24_L14036_C104/carry[3] ),.C1(\add_90_I24_L14036_C104/carry[4] ),.SO(N1225));
  HADDX1 desc1217(.A0(N1215),.B0(\add_90_I24_L14036_C104/carry[4] ),.C1(\add_90_I24_L14036_C104/carry[5] ),.SO(N1226));
  HADDX1 desc1218(.A0(N1195),.B0(N1194),.C1(\add_90_I23_L14036_C104/carry[2] ),.SO(N1206));
  HADDX1 desc1219(.A0(N1196),.B0(\add_90_I23_L14036_C104/carry[2] ),.C1(\add_90_I23_L14036_C104/carry[3] ),.SO(N1207));
  HADDX1 desc1220(.A0(N1197),.B0(\add_90_I23_L14036_C104/carry[3] ),.C1(\add_90_I23_L14036_C104/carry[4] ),.SO(N1208));
  HADDX1 desc1221(.A0(N1198),.B0(\add_90_I23_L14036_C104/carry[4] ),.C1(\add_90_I23_L14036_C104/carry[5] ),.SO(N1209));
  HADDX1 desc1222(.A0(N1178),.B0(N1177),.C1(\add_90_I22_L14036_C104/carry[2] ),.SO(N1189));
  HADDX1 desc1223(.A0(N1179),.B0(\add_90_I22_L14036_C104/carry[2] ),.C1(\add_90_I22_L14036_C104/carry[3] ),.SO(N1190));
  HADDX1 desc1224(.A0(N1180),.B0(\add_90_I22_L14036_C104/carry[3] ),.C1(\add_90_I22_L14036_C104/carry[4] ),.SO(N1191));
  HADDX1 desc1225(.A0(N1181),.B0(\add_90_I22_L14036_C104/carry[4] ),.C1(\add_90_I22_L14036_C104/carry[5] ),.SO(N1192));
  HADDX1 desc1226(.A0(N1161),.B0(N1160),.C1(\add_90_I21_L14036_C104/carry[2] ),.SO(N1172));
  HADDX1 desc1227(.A0(N1162),.B0(\add_90_I21_L14036_C104/carry[2] ),.C1(\add_90_I21_L14036_C104/carry[3] ),.SO(N1173));
  HADDX1 desc1228(.A0(N1163),.B0(\add_90_I21_L14036_C104/carry[3] ),.C1(\add_90_I21_L14036_C104/carry[4] ),.SO(N1174));
  HADDX1 desc1229(.A0(N1164),.B0(\add_90_I21_L14036_C104/carry[4] ),.C1(\add_90_I21_L14036_C104/carry[5] ),.SO(N1175));
  HADDX1 desc1230(.A0(N1144),.B0(N1143),.C1(\add_90_I20_L14036_C104/carry[2] ),.SO(N1155));
  HADDX1 desc1231(.A0(N1145),.B0(\add_90_I20_L14036_C104/carry[2] ),.C1(\add_90_I20_L14036_C104/carry[3] ),.SO(N1156));
  HADDX1 desc1232(.A0(N1146),.B0(\add_90_I20_L14036_C104/carry[3] ),.C1(\add_90_I20_L14036_C104/carry[4] ),.SO(N1157));
  HADDX1 desc1233(.A0(N1147),.B0(\add_90_I20_L14036_C104/carry[4] ),.C1(\add_90_I20_L14036_C104/carry[5] ),.SO(N1158));
  HADDX1 desc1234(.A0(N1127),.B0(N1126),.C1(\add_90_I19_L14036_C104/carry[2] ),.SO(N1138));
  HADDX1 desc1235(.A0(N1128),.B0(\add_90_I19_L14036_C104/carry[2] ),.C1(\add_90_I19_L14036_C104/carry[3] ),.SO(N1139));
  HADDX1 desc1236(.A0(N1129),.B0(\add_90_I19_L14036_C104/carry[3] ),.C1(\add_90_I19_L14036_C104/carry[4] ),.SO(N1140));
  HADDX1 desc1237(.A0(N1130),.B0(\add_90_I19_L14036_C104/carry[4] ),.C1(\add_90_I19_L14036_C104/carry[5] ),.SO(N1141));
  HADDX1 desc1238(.A0(N1110),.B0(N1109),.C1(\add_90_I18_L14036_C104/carry[2] ),.SO(N1121));
  HADDX1 desc1239(.A0(N1111),.B0(\add_90_I18_L14036_C104/carry[2] ),.C1(\add_90_I18_L14036_C104/carry[3] ),.SO(N1122));
  HADDX1 desc1240(.A0(N1112),.B0(\add_90_I18_L14036_C104/carry[3] ),.C1(\add_90_I18_L14036_C104/carry[4] ),.SO(N1123));
  HADDX1 desc1241(.A0(N1113),.B0(\add_90_I18_L14036_C104/carry[4] ),.C1(\add_90_I18_L14036_C104/carry[5] ),.SO(N1124));
  HADDX1 desc1242(.A0(N1093),.B0(N1092),.C1(\add_90_I17_L14036_C104/carry[2] ),.SO(N1104));
  HADDX1 desc1243(.A0(N1094),.B0(\add_90_I17_L14036_C104/carry[2] ),.C1(\add_90_I17_L14036_C104/carry[3] ),.SO(N1105));
  HADDX1 desc1244(.A0(N1095),.B0(\add_90_I17_L14036_C104/carry[3] ),.C1(\add_90_I17_L14036_C104/carry[4] ),.SO(N1106));
  HADDX1 desc1245(.A0(N1096),.B0(\add_90_I17_L14036_C104/carry[4] ),.C1(\add_90_I17_L14036_C104/carry[5] ),.SO(N1107));
  HADDX1 desc1246(.A0(N1076),.B0(N1075),.C1(\add_90_I16_L14036_C104/carry[2] ),.SO(N1087));
  HADDX1 desc1247(.A0(N1077),.B0(\add_90_I16_L14036_C104/carry[2] ),.C1(\add_90_I16_L14036_C104/carry[3] ),.SO(N1088));
  HADDX1 desc1248(.A0(N1078),.B0(\add_90_I16_L14036_C104/carry[3] ),.C1(\add_90_I16_L14036_C104/carry[4] ),.SO(N1089));
  HADDX1 desc1249(.A0(N1079),.B0(\add_90_I16_L14036_C104/carry[4] ),.C1(\add_90_I16_L14036_C104/carry[5] ),.SO(N1090));
  HADDX1 desc1250(.A0(N1059),.B0(N1058),.C1(\add_90_I15_L14036_C104/carry[2] ),.SO(N1070));
  HADDX1 desc1251(.A0(N1060),.B0(\add_90_I15_L14036_C104/carry[2] ),.C1(\add_90_I15_L14036_C104/carry[3] ),.SO(N1071));
  HADDX1 desc1252(.A0(N1061),.B0(\add_90_I15_L14036_C104/carry[3] ),.C1(\add_90_I15_L14036_C104/carry[4] ),.SO(N1072));
  HADDX1 desc1253(.A0(N1062),.B0(\add_90_I15_L14036_C104/carry[4] ),.C1(\add_90_I15_L14036_C104/carry[5] ),.SO(N1073));
  HADDX1 desc1254(.A0(N1042),.B0(N1041),.C1(\add_90_I14_L14036_C104/carry[2] ),.SO(N1053));
  HADDX1 desc1255(.A0(N1043),.B0(\add_90_I14_L14036_C104/carry[2] ),.C1(\add_90_I14_L14036_C104/carry[3] ),.SO(N1054));
  HADDX1 desc1256(.A0(N1044),.B0(\add_90_I14_L14036_C104/carry[3] ),.C1(\add_90_I14_L14036_C104/carry[4] ),.SO(N1055));
  HADDX1 desc1257(.A0(N1045),.B0(\add_90_I14_L14036_C104/carry[4] ),.C1(\add_90_I14_L14036_C104/carry[5] ),.SO(N1056));
  HADDX1 desc1258(.A0(N1025),.B0(N1024),.C1(\add_90_I13_L14036_C104/carry[2] ),.SO(N1036));
  HADDX1 desc1259(.A0(N1026),.B0(\add_90_I13_L14036_C104/carry[2] ),.C1(\add_90_I13_L14036_C104/carry[3] ),.SO(N1037));
  HADDX1 desc1260(.A0(N1027),.B0(\add_90_I13_L14036_C104/carry[3] ),.C1(\add_90_I13_L14036_C104/carry[4] ),.SO(N1038));
  HADDX1 desc1261(.A0(N1028),.B0(\add_90_I13_L14036_C104/carry[4] ),.C1(\add_90_I13_L14036_C104/carry[5] ),.SO(N1039));
  HADDX1 desc1262(.A0(N1008),.B0(N1007),.C1(\add_90_I12_L14036_C104/carry[2] ),.SO(N1019));
  HADDX1 desc1263(.A0(N1009),.B0(\add_90_I12_L14036_C104/carry[2] ),.C1(\add_90_I12_L14036_C104/carry[3] ),.SO(N1020));
  HADDX1 desc1264(.A0(N1010),.B0(\add_90_I12_L14036_C104/carry[3] ),.C1(\add_90_I12_L14036_C104/carry[4] ),.SO(N1021));
  HADDX1 desc1265(.A0(N1011),.B0(\add_90_I12_L14036_C104/carry[4] ),.C1(\add_90_I12_L14036_C104/carry[5] ),.SO(N1022));
  HADDX1 desc1266(.A0(N991),.B0(N990),.C1(\add_90_I11_L14036_C104/carry[2] ),.SO(N1002));
  HADDX1 desc1267(.A0(N992),.B0(\add_90_I11_L14036_C104/carry[2] ),.C1(\add_90_I11_L14036_C104/carry[3] ),.SO(N1003));
  HADDX1 desc1268(.A0(N993),.B0(\add_90_I11_L14036_C104/carry[3] ),.C1(\add_90_I11_L14036_C104/carry[4] ),.SO(N1004));
  HADDX1 desc1269(.A0(N994),.B0(\add_90_I11_L14036_C104/carry[4] ),.C1(\add_90_I11_L14036_C104/carry[5] ),.SO(N1005));
  HADDX1 desc1270(.A0(N974),.B0(N973),.C1(\add_90_I10_L14036_C104/carry[2] ),.SO(N985));
  HADDX1 desc1271(.A0(N975),.B0(\add_90_I10_L14036_C104/carry[2] ),.C1(\add_90_I10_L14036_C104/carry[3] ),.SO(N986));
  HADDX1 desc1272(.A0(N976),.B0(\add_90_I10_L14036_C104/carry[3] ),.C1(\add_90_I10_L14036_C104/carry[4] ),.SO(N987));
  HADDX1 desc1273(.A0(N977),.B0(\add_90_I10_L14036_C104/carry[4] ),.C1(\add_90_I10_L14036_C104/carry[5] ),.SO(N988));
  HADDX1 desc1274(.A0(N957),.B0(N956),.C1(\add_90_I9_L14036_C104/carry[2] ),.SO(N968));
  HADDX1 desc1275(.A0(N958),.B0(\add_90_I9_L14036_C104/carry[2] ),.C1(\add_90_I9_L14036_C104/carry[3] ),.SO(N969));
  HADDX1 desc1276(.A0(N959),.B0(\add_90_I9_L14036_C104/carry[3] ),.C1(\add_90_I9_L14036_C104/carry[4] ),.SO(N970));
  HADDX1 desc1277(.A0(N960),.B0(\add_90_I9_L14036_C104/carry[4] ),.C1(\add_90_I9_L14036_C104/carry[5] ),.SO(N971));
  HADDX1 desc1278(.A0(N940),.B0(N939),.C1(\add_90_I8_L14036_C104/carry[2] ),.SO(N951));
  HADDX1 desc1279(.A0(N941),.B0(\add_90_I8_L14036_C104/carry[2] ),.C1(\add_90_I8_L14036_C104/carry[3] ),.SO(N952));
  HADDX1 desc1280(.A0(N942),.B0(\add_90_I8_L14036_C104/carry[3] ),.C1(\add_90_I8_L14036_C104/carry[4] ),.SO(N953));
  HADDX1 desc1281(.A0(N943),.B0(\add_90_I8_L14036_C104/carry[4] ),.C1(\add_90_I8_L14036_C104/carry[5] ),.SO(N954));
  HADDX1 desc1282(.A0(N923),.B0(N922),.C1(\add_90_I7_L14036_C104/carry[2] ),.SO(N934));
  HADDX1 desc1283(.A0(N924),.B0(\add_90_I7_L14036_C104/carry[2] ),.C1(\add_90_I7_L14036_C104/carry[3] ),.SO(N935));
  HADDX1 desc1284(.A0(N925),.B0(\add_90_I7_L14036_C104/carry[3] ),.C1(\add_90_I7_L14036_C104/carry[4] ),.SO(N936));
  HADDX1 desc1285(.A0(N926),.B0(\add_90_I7_L14036_C104/carry[4] ),.C1(N938),.SO(N937));
  HADDX1 desc1286(.A0(N907),.B0(N906),.C1(\add_90_I6_L14036_C104/carry[2] ),.SO(N917));
  HADDX1 desc1287(.A0(N908),.B0(\add_90_I6_L14036_C104/carry[2] ),.C1(\add_90_I6_L14036_C104/carry[3] ),.SO(N918));
  HADDX1 desc1288(.A0(N909),.B0(\add_90_I6_L14036_C104/carry[3] ),.C1(N920),.SO(N919));
  HADDX1 desc1289(.A0(N893),.B0(N892),.C1(\add_90_I5_L14036_C104/carry[2] ),.SO(N902));
  HADDX1 desc1290(.A0(N894),.B0(\add_90_I5_L14036_C104/carry[2] ),.C1(N904),.SO(N903));
  HADDX1 desc1291(.A0(N549),.B0(N548),.C1(\add_90_I24_L14036_C103/carry[2] ),.SO(N560));
  HADDX1 desc1292(.A0(N550),.B0(\add_90_I24_L14036_C103/carry[2] ),.C1(\add_90_I24_L14036_C103/carry[3] ),.SO(N561));
  HADDX1 desc1293(.A0(N551),.B0(\add_90_I24_L14036_C103/carry[3] ),.C1(\add_90_I24_L14036_C103/carry[4] ),.SO(N562));
  HADDX1 desc1294(.A0(N552),.B0(\add_90_I24_L14036_C103/carry[4] ),.C1(\add_90_I24_L14036_C103/carry[5] ),.SO(N563));
  HADDX1 desc1295(.A0(N532),.B0(N531),.C1(\add_90_I23_L14036_C103/carry[2] ),.SO(N543));
  HADDX1 desc1296(.A0(N533),.B0(\add_90_I23_L14036_C103/carry[2] ),.C1(\add_90_I23_L14036_C103/carry[3] ),.SO(N544));
  HADDX1 desc1297(.A0(N534),.B0(\add_90_I23_L14036_C103/carry[3] ),.C1(\add_90_I23_L14036_C103/carry[4] ),.SO(N545));
  HADDX1 desc1298(.A0(N535),.B0(\add_90_I23_L14036_C103/carry[4] ),.C1(\add_90_I23_L14036_C103/carry[5] ),.SO(N546));
  HADDX1 desc1299(.A0(N515),.B0(N514),.C1(\add_90_I22_L14036_C103/carry[2] ),.SO(N526));
  HADDX1 desc1300(.A0(N516),.B0(\add_90_I22_L14036_C103/carry[2] ),.C1(\add_90_I22_L14036_C103/carry[3] ),.SO(N527));
  HADDX1 desc1301(.A0(N517),.B0(\add_90_I22_L14036_C103/carry[3] ),.C1(\add_90_I22_L14036_C103/carry[4] ),.SO(N528));
  HADDX1 desc1302(.A0(N518),.B0(\add_90_I22_L14036_C103/carry[4] ),.C1(\add_90_I22_L14036_C103/carry[5] ),.SO(N529));
  HADDX1 desc1303(.A0(N498),.B0(N497),.C1(\add_90_I21_L14036_C103/carry[2] ),.SO(N509));
  HADDX1 desc1304(.A0(N499),.B0(\add_90_I21_L14036_C103/carry[2] ),.C1(\add_90_I21_L14036_C103/carry[3] ),.SO(N510));
  HADDX1 desc1305(.A0(N500),.B0(\add_90_I21_L14036_C103/carry[3] ),.C1(\add_90_I21_L14036_C103/carry[4] ),.SO(N511));
  HADDX1 desc1306(.A0(N501),.B0(\add_90_I21_L14036_C103/carry[4] ),.C1(\add_90_I21_L14036_C103/carry[5] ),.SO(N512));
  HADDX1 desc1307(.A0(N481),.B0(N480),.C1(\add_90_I20_L14036_C103/carry[2] ),.SO(N492));
  HADDX1 desc1308(.A0(N482),.B0(\add_90_I20_L14036_C103/carry[2] ),.C1(\add_90_I20_L14036_C103/carry[3] ),.SO(N493));
  HADDX1 desc1309(.A0(N483),.B0(\add_90_I20_L14036_C103/carry[3] ),.C1(\add_90_I20_L14036_C103/carry[4] ),.SO(N494));
  HADDX1 desc1310(.A0(N484),.B0(\add_90_I20_L14036_C103/carry[4] ),.C1(\add_90_I20_L14036_C103/carry[5] ),.SO(N495));
  HADDX1 desc1311(.A0(N464),.B0(N463),.C1(\add_90_I19_L14036_C103/carry[2] ),.SO(N475));
  HADDX1 desc1312(.A0(N465),.B0(\add_90_I19_L14036_C103/carry[2] ),.C1(\add_90_I19_L14036_C103/carry[3] ),.SO(N476));
  HADDX1 desc1313(.A0(N466),.B0(\add_90_I19_L14036_C103/carry[3] ),.C1(\add_90_I19_L14036_C103/carry[4] ),.SO(N477));
  HADDX1 desc1314(.A0(N467),.B0(\add_90_I19_L14036_C103/carry[4] ),.C1(\add_90_I19_L14036_C103/carry[5] ),.SO(N478));
  HADDX1 desc1315(.A0(N447),.B0(N446),.C1(\add_90_I18_L14036_C103/carry[2] ),.SO(N458));
  HADDX1 desc1316(.A0(N448),.B0(\add_90_I18_L14036_C103/carry[2] ),.C1(\add_90_I18_L14036_C103/carry[3] ),.SO(N459));
  HADDX1 desc1317(.A0(N449),.B0(\add_90_I18_L14036_C103/carry[3] ),.C1(\add_90_I18_L14036_C103/carry[4] ),.SO(N460));
  HADDX1 desc1318(.A0(N450),.B0(\add_90_I18_L14036_C103/carry[4] ),.C1(\add_90_I18_L14036_C103/carry[5] ),.SO(N461));
  HADDX1 desc1319(.A0(N430),.B0(N429),.C1(\add_90_I17_L14036_C103/carry[2] ),.SO(N441));
  HADDX1 desc1320(.A0(N431),.B0(\add_90_I17_L14036_C103/carry[2] ),.C1(\add_90_I17_L14036_C103/carry[3] ),.SO(N442));
  HADDX1 desc1321(.A0(N432),.B0(\add_90_I17_L14036_C103/carry[3] ),.C1(\add_90_I17_L14036_C103/carry[4] ),.SO(N443));
  HADDX1 desc1322(.A0(N433),.B0(\add_90_I17_L14036_C103/carry[4] ),.C1(\add_90_I17_L14036_C103/carry[5] ),.SO(N444));
  HADDX1 desc1323(.A0(N413),.B0(N412),.C1(\add_90_I16_L14036_C103/carry[2] ),.SO(N424));
  HADDX1 desc1324(.A0(N414),.B0(\add_90_I16_L14036_C103/carry[2] ),.C1(\add_90_I16_L14036_C103/carry[3] ),.SO(N425));
  HADDX1 desc1325(.A0(N415),.B0(\add_90_I16_L14036_C103/carry[3] ),.C1(\add_90_I16_L14036_C103/carry[4] ),.SO(N426));
  HADDX1 desc1326(.A0(N416),.B0(\add_90_I16_L14036_C103/carry[4] ),.C1(\add_90_I16_L14036_C103/carry[5] ),.SO(N427));
  HADDX1 desc1327(.A0(N396),.B0(N395),.C1(\add_90_I15_L14036_C103/carry[2] ),.SO(N407));
  HADDX1 desc1328(.A0(N397),.B0(\add_90_I15_L14036_C103/carry[2] ),.C1(\add_90_I15_L14036_C103/carry[3] ),.SO(N408));
  HADDX1 desc1329(.A0(N398),.B0(\add_90_I15_L14036_C103/carry[3] ),.C1(\add_90_I15_L14036_C103/carry[4] ),.SO(N409));
  HADDX1 desc1330(.A0(N399),.B0(\add_90_I15_L14036_C103/carry[4] ),.C1(\add_90_I15_L14036_C103/carry[5] ),.SO(N410));
  HADDX1 desc1331(.A0(N379),.B0(N378),.C1(\add_90_I14_L14036_C103/carry[2] ),.SO(N390));
  HADDX1 desc1332(.A0(N380),.B0(\add_90_I14_L14036_C103/carry[2] ),.C1(\add_90_I14_L14036_C103/carry[3] ),.SO(N391));
  HADDX1 desc1333(.A0(N381),.B0(\add_90_I14_L14036_C103/carry[3] ),.C1(\add_90_I14_L14036_C103/carry[4] ),.SO(N392));
  HADDX1 desc1334(.A0(N382),.B0(\add_90_I14_L14036_C103/carry[4] ),.C1(\add_90_I14_L14036_C103/carry[5] ),.SO(N393));
  HADDX1 desc1335(.A0(N362),.B0(N361),.C1(\add_90_I13_L14036_C103/carry[2] ),.SO(N373));
  HADDX1 desc1336(.A0(N363),.B0(\add_90_I13_L14036_C103/carry[2] ),.C1(\add_90_I13_L14036_C103/carry[3] ),.SO(N374));
  HADDX1 desc1337(.A0(N364),.B0(\add_90_I13_L14036_C103/carry[3] ),.C1(\add_90_I13_L14036_C103/carry[4] ),.SO(N375));
  HADDX1 desc1338(.A0(N365),.B0(\add_90_I13_L14036_C103/carry[4] ),.C1(\add_90_I13_L14036_C103/carry[5] ),.SO(N376));
  HADDX1 desc1339(.A0(N345),.B0(N344),.C1(\add_90_I12_L14036_C103/carry[2] ),.SO(N356));
  HADDX1 desc1340(.A0(N346),.B0(\add_90_I12_L14036_C103/carry[2] ),.C1(\add_90_I12_L14036_C103/carry[3] ),.SO(N357));
  HADDX1 desc1341(.A0(N347),.B0(\add_90_I12_L14036_C103/carry[3] ),.C1(\add_90_I12_L14036_C103/carry[4] ),.SO(N358));
  HADDX1 desc1342(.A0(N348),.B0(\add_90_I12_L14036_C103/carry[4] ),.C1(\add_90_I12_L14036_C103/carry[5] ),.SO(N359));
  HADDX1 desc1343(.A0(N328),.B0(N327),.C1(\add_90_I11_L14036_C103/carry[2] ),.SO(N339));
  HADDX1 desc1344(.A0(N329),.B0(\add_90_I11_L14036_C103/carry[2] ),.C1(\add_90_I11_L14036_C103/carry[3] ),.SO(N340));
  HADDX1 desc1345(.A0(N330),.B0(\add_90_I11_L14036_C103/carry[3] ),.C1(\add_90_I11_L14036_C103/carry[4] ),.SO(N341));
  HADDX1 desc1346(.A0(N331),.B0(\add_90_I11_L14036_C103/carry[4] ),.C1(\add_90_I11_L14036_C103/carry[5] ),.SO(N342));
  HADDX1 desc1347(.A0(N311),.B0(N310),.C1(\add_90_I10_L14036_C103/carry[2] ),.SO(N322));
  HADDX1 desc1348(.A0(N312),.B0(\add_90_I10_L14036_C103/carry[2] ),.C1(\add_90_I10_L14036_C103/carry[3] ),.SO(N323));
  HADDX1 desc1349(.A0(N313),.B0(\add_90_I10_L14036_C103/carry[3] ),.C1(\add_90_I10_L14036_C103/carry[4] ),.SO(N324));
  HADDX1 desc1350(.A0(N314),.B0(\add_90_I10_L14036_C103/carry[4] ),.C1(\add_90_I10_L14036_C103/carry[5] ),.SO(N325));
  HADDX1 desc1351(.A0(N294),.B0(N293),.C1(\add_90_I9_L14036_C103/carry[2] ),.SO(N305));
  HADDX1 desc1352(.A0(N295),.B0(\add_90_I9_L14036_C103/carry[2] ),.C1(\add_90_I9_L14036_C103/carry[3] ),.SO(N306));
  HADDX1 desc1353(.A0(N296),.B0(\add_90_I9_L14036_C103/carry[3] ),.C1(\add_90_I9_L14036_C103/carry[4] ),.SO(N307));
  HADDX1 desc1354(.A0(N297),.B0(\add_90_I9_L14036_C103/carry[4] ),.C1(\add_90_I9_L14036_C103/carry[5] ),.SO(N308));
  HADDX1 desc1355(.A0(N277),.B0(N276),.C1(\add_90_I8_L14036_C103/carry[2] ),.SO(N288));
  HADDX1 desc1356(.A0(N278),.B0(\add_90_I8_L14036_C103/carry[2] ),.C1(\add_90_I8_L14036_C103/carry[3] ),.SO(N289));
  HADDX1 desc1357(.A0(N279),.B0(\add_90_I8_L14036_C103/carry[3] ),.C1(\add_90_I8_L14036_C103/carry[4] ),.SO(N290));
  HADDX1 desc1358(.A0(N280),.B0(\add_90_I8_L14036_C103/carry[4] ),.C1(\add_90_I8_L14036_C103/carry[5] ),.SO(N291));
  HADDX1 desc1359(.A0(N260),.B0(N259),.C1(\add_90_I7_L14036_C103/carry[2] ),.SO(N271));
  HADDX1 desc1360(.A0(N261),.B0(\add_90_I7_L14036_C103/carry[2] ),.C1(\add_90_I7_L14036_C103/carry[3] ),.SO(N272));
  HADDX1 desc1361(.A0(N262),.B0(\add_90_I7_L14036_C103/carry[3] ),.C1(\add_90_I7_L14036_C103/carry[4] ),.SO(N273));
  HADDX1 desc1362(.A0(N263),.B0(\add_90_I7_L14036_C103/carry[4] ),.C1(N275),.SO(N274));
  HADDX1 desc1363(.A0(N244),.B0(N243),.C1(\add_90_I6_L14036_C103/carry[2] ),.SO(N254));
  HADDX1 desc1364(.A0(N245),.B0(\add_90_I6_L14036_C103/carry[2] ),.C1(\add_90_I6_L14036_C103/carry[3] ),.SO(N255));
  HADDX1 desc1365(.A0(N246),.B0(\add_90_I6_L14036_C103/carry[3] ),.C1(N257),.SO(N256));
  HADDX1 desc1366(.A0(N230),.B0(N229),.C1(\add_90_I5_L14036_C103/carry[2] ),.SO(N239));
  HADDX1 desc1367(.A0(N231),.B0(\add_90_I5_L14036_C103/carry[2] ),.C1(N241),.SO(N240));
  NAND2X0 U3(.IN1(n611),.IN2(n144),.QN(n548));
  NAND2X0 U5(.IN1(n613),.IN2(n144),.QN(n570));
  NAND2X0 U6(.IN1(n324),.IN2(n377),.QN(n361));
  NAND2X0 U7(.IN1(n309),.IN2(n378),.QN(n310));
  NBUFFX2 U8(.INP(opb_i[18:18]),.Z(n16));
  NAND2X0 U9(.IN1(n220),.IN2(n109),.QN(n257));
  NOR2X0 U10(.IN1(s_dvd_zeros[5:5]),.IN2(n451),.QN(dvdnd_50_o[43:43]));
  INVX0 U11(.INP(s_dvd_zeros[5:5]),.ZN(n49));
  INVX0 U12(.INP(n492),.ZN(n80));
  OA21X1 U13(.IN1(n155),.IN2(n156),.IN3(n95),.Q(n20));
  INVX0 U14(.INP(s_dvd_zeros[2:2]),.ZN(n93));
  INVX0 U15(.INP(s_dvd_zeros[3:3]),.ZN(n94));
  INVX0 U16(.INP(s_dvd_zeros[4:4]),.ZN(n54));
  INVX0 U17(.INP(n509),.ZN(n76));
  OA21X1 U18(.IN1(n155),.IN2(n156),.IN3(n95),.Q(n19));
  OA21X1 U19(.IN1(n155),.IN2(n156),.IN3(n95),.Q(s_dvd_zeros[5:5]));
  NAND2X0 U20(.IN1(n509),.IN2(n94),.QN(n466));
  NAND2X0 U21(.IN1(n507),.IN2(n94),.QN(n444));
  INVX0 U22(.INP(n432),.ZN(n78));
  NOR2X0 U23(.IN1(n75),.IN2(s_dvd_zeros[3:3]),.QN(n505));
  NOR2X0 U24(.IN1(n19),.IN2(n445),.QN(dvdnd_50_o[42:42]));
  NOR2X0 U25(.IN1(n19),.IN2(n465),.QN(dvdnd_50_o[45:45]));
  NOR2X0 U26(.IN1(n20),.IN2(n458),.QN(dvdnd_50_o[44:44]));
  INVX0 U27(.INP(n506),.ZN(n69));
  INVX0 U28(.INP(n470),.ZN(n83));
  INVX0 U29(.INP(n487),.ZN(n88));
  INVX0 U30(.INP(n478),.ZN(n86));
  NBUFFX2 U31(.INP(n91),.Z(n21));
  NBUFFX2 U32(.INP(n91),.Z(n22));
  NOR2X0 U33(.IN1(s_div_zeros[5:5]),.IN2(n555),.QN(dvsor_27_o[17:17]));
  INVX0 U34(.INP(n610),.ZN(n119));
  INVX0 U35(.INP(s_div_zeros[5:5]),.ZN(n59));
  INVX0 U36(.INP(N430),.ZN(n106));
  INVX0 U37(.INP(N431),.ZN(n102));
  INVX0 U38(.INP(n596),.ZN(n130));
  NBUFFX2 U39(.INP(n141),.Z(n23));
  NBUFFX2 U40(.INP(n141),.Z(n24));
  INVX0 U41(.INP(N432),.ZN(n98));
  INVX0 U42(.INP(N433),.ZN(n57));
  NOR2X0 U43(.IN1(n38),.IN2(n40),.QN(n247));
  NOR2X0 U44(.IN1(n248),.IN2(n35),.QN(n249));
  NAND2X0 U45(.IN1(n249),.IN2(n250),.QN(n181));
  INVX0 U46(.INP(n250),.ZN(n118));
  NAND2X0 U47(.IN1(n118),.IN2(n171),.QN(n169));
  NOR2X0 U48(.IN1(n247),.IN2(n40),.QN(n179));
  NAND2X0 U49(.IN1(n247),.IN2(n248),.QN(n168));
  NOR2X0 U50(.IN1(n243),.IN2(n111),.QN(n160));
  NOR2X0 U51(.IN1(n254),.IN2(n28),.QN(n255));
  INVX0 U52(.INP(n239),.ZN(n116));
  INVX0 U53(.INP(n243),.ZN(n112));
  INVX0 U54(.INP(n240),.ZN(n115));
  INVX0 U55(.INP(n241),.ZN(n113));
  INVX0 U56(.INP(n242),.ZN(n114));
  INVX0 U57(.INP(n214),.ZN(n111));
  NOR2X0 U58(.IN1(n254),.IN2(n255),.QN(n175));
  NOR2X0 U59(.IN1(n239),.IN2(n115),.QN(n157));
  NOR2X0 U60(.IN1(n240),.IN2(n114),.QN(n159));
  NOR2X0 U61(.IN1(n241),.IN2(n112),.QN(n163));
  NOR2X0 U62(.IN1(n242),.IN2(n113),.QN(n164));
  NOR2X0 U63(.IN1(n116),.IN2(n47),.QN(n158));
  OA21X1 U64(.IN1(n182),.IN2(n183),.IN3(n95),.Q(s_dvd_zeros[4:4]));
  OA21X1 U65(.IN1(n193),.IN2(n194),.IN3(n95),.Q(s_dvd_zeros[3:3]));
  INVX0 U66(.INP(N417),.ZN(n53));
  INVX0 U67(.INP(N468),.ZN(n50));
  NOR2X0 U68(.IN1(n172),.IN2(n173),.QN(n170));
  INVX0 U69(.INP(s_dvd_zeros[1:1]),.ZN(n92));
  OA21X1 U70(.IN1(n259),.IN2(n260),.IN3(n145),.Q(n18));
  NAND2X0 U71(.IN1(n433),.IN2(n93),.QN(n459));
  INVX0 U72(.INP(N412),.ZN(N423));
  NOR2X0 U73(.IN1(n446),.IN2(s_dvd_zeros[2:2]),.QN(n509));
  INVX0 U74(.INP(N361),.ZN(N372));
  NOR2X0 U75(.IN1(n416),.IN2(s_dvd_zeros[2:2]),.QN(n507));
  AND2X1 U76(.IN1(N275),.IN2(n46),.Q(n10));
  INVX0 U77(.INP(n447),.ZN(n85));
  INVX0 U78(.INP(n422),.ZN(n81));
  INVX0 U79(.INP(n440),.ZN(n82));
  INVX0 U80(.INP(n434),.ZN(n75));
  NOR2X0 U81(.IN1(n20),.IN2(n482),.QN(dvdnd_50_o[47:47]));
  INVX0 U82(.INP(n479),.ZN(n87));
  NOR2X0 U83(.IN1(s_dvd_zeros[5:5]),.IN2(n474),.QN(dvdnd_50_o[46:46]));
  INVX0 U84(.INP(n471),.ZN(n84));
  INVX0 U85(.INP(n424),.ZN(n79));
  INVX0 U86(.INP(n421),.ZN(n77));
  INVX0 U87(.INP(N463),.ZN(N474));
  INVX0 U88(.INP(N531),.ZN(N542));
  INVX0 U89(.INP(N497),.ZN(N508));
  INVX0 U90(.INP(N378),.ZN(N389));
  INVX0 U91(.INP(n496),.ZN(n90));
  INVX0 U92(.INP(s_div_zeros[1:1]),.ZN(n142));
  INVX0 U93(.INP(s_div_zeros[2:2]),.ZN(n143));
  INVX0 U94(.INP(s_div_zeros[3:3]),.ZN(n144));
  INVX0 U95(.INP(s_div_zeros[4:4]),.ZN(n64));
  INVX0 U96(.INP(n613),.ZN(n126));
  OA21X1 U97(.IN1(n259),.IN2(n260),.IN3(n145),.Q(n17));
  NAND2X0 U98(.IN1(n537),.IN2(n143),.QN(n563));
  OA21X1 U99(.IN1(n259),.IN2(n260),.IN3(n145),.Q(s_div_zeros[5:5]));
  NOR2X0 U100(.IN1(n550),.IN2(s_div_zeros[2:2]),.QN(n613));
  NOR2X0 U101(.IN1(n520),.IN2(s_div_zeros[2:2]),.QN(n611));
  NOR2X0 U102(.IN1(n125),.IN2(s_div_zeros[3:3]),.QN(n609));
  INVX0 U103(.INP(n536),.ZN(n128));
  NOR2X0 U104(.IN1(n18),.IN2(n586),.QN(dvsor_27_o[21:21]));
  INVX0 U105(.INP(n583),.ZN(n137));
  NOR2X0 U106(.IN1(n18),.IN2(n562),.QN(dvsor_27_o[18:18]));
  INVX0 U107(.INP(n538),.ZN(n125));
  NOR2X0 U108(.IN1(n17),.IN2(n569),.QN(dvsor_27_o[19:19]));
  NOR2X0 U109(.IN1(n17),.IN2(n549),.QN(dvsor_27_o[16:16]));
  NOR2X0 U110(.IN1(s_div_zeros[5:5]),.IN2(n578),.QN(dvsor_27_o[20:20]));
  INVX0 U111(.INP(n575),.ZN(n134));
  INVX0 U112(.INP(s_dvd_zeros[0:0]),.ZN(n91));
  INVX0 U113(.INP(N434),.ZN(n52));
  INVX0 U114(.INP(N451),.ZN(n51));
  INVX0 U115(.INP(N447),.ZN(n105));
  INVX0 U116(.INP(N448),.ZN(n101));
  INVX0 U117(.INP(N449),.ZN(n97));
  INVX0 U118(.INP(N450),.ZN(n56));
  INVX0 U119(.INP(n591),.ZN(n138));
  INVX0 U120(.INP(n574),.ZN(n133));
  INVX0 U121(.INP(n600),.ZN(n140));
  INVX0 U122(.INP(n582),.ZN(n136));
  INVX0 U123(.INP(N464),.ZN(n104));
  INVX0 U124(.INP(N465),.ZN(n100));
  INVX0 U125(.INP(N466),.ZN(n96));
  INVX0 U126(.INP(N467),.ZN(n55));
  INVX0 U127(.INP(s_div_zeros[0:0]),.ZN(n141));
  INVX0 U128(.INP(N413),.ZN(n107));
  INVX0 U129(.INP(N414),.ZN(n103));
  INVX0 U130(.INP(N415),.ZN(n99));
  INVX0 U131(.INP(N416),.ZN(n58));
  NOR2X0 U132(.IN1(n347),.IN2(n379),.QN(n264));
  NOR2X0 U133(.IN1(n345),.IN2(n380),.QN(n267));
  INVX0 U134(.INP(n343),.ZN(n384));
  INVX0 U135(.INP(n318),.ZN(n379));
  INVX0 U136(.INP(n347),.ZN(n380));
  INVX0 U137(.INP(n346),.ZN(n382));
  INVX0 U138(.INP(n345),.ZN(n381));
  INVX0 U139(.INP(n344),.ZN(n383));
  NAND2X0 U140(.IN1(n160),.IN2(N361),.QN(n235));
  NAND2X0 U141(.IN1(n160),.IN2(N363),.QN(n208));
  NAND2X0 U142(.IN1(n160),.IN2(N362),.QN(n222));
  NAND2X1 U143(.IN1(n118),.IN2(n33),.QN(n171));
  NAND2X1 U144(.IN1(n247),.IN2(n37),.QN(n248));
  NOR2X0 U145(.IN1(n344),.IN2(n382),.QN(n263));
  NOR2X0 U146(.IN1(n343),.IN2(n383),.QN(n261));
  NAND2X0 U147(.IN1(n249),.IN2(n34),.QN(n250));
  NOR2X0 U148(.IN1(n346),.IN2(n381),.QN(n268));
  INVX0 U149(.INP(n354),.ZN(n393));
  NAND2X0 U150(.IN1(n393),.IN2(n275),.QN(n273));
  INVX0 U151(.INP(n206),.ZN(n95));
  NAND2X1 U152(.IN1(n113),.IN2(n42),.QN(n243));
  NAND2X1 U153(.IN1(n255),.IN2(n27),.QN(n256));
  NAND2X0 U154(.IN1(n114),.IN2(n43),.QN(n241));
  NAND2X0 U155(.IN1(n116),.IN2(n45),.QN(n240));
  NAND2X0 U156(.IN1(n115),.IN2(n44),.QN(n242));
  NAND2X0 U157(.IN1(n46),.IN2(n48),.QN(n239));
  NAND2X1 U158(.IN1(n112),.IN2(n117),.QN(n214));
  INVX0 U159(.INP(n310),.ZN(n145));
  NAND2X1 U160(.IN1(n30),.IN2(n32),.QN(n254));
  INVX0 U161(.INP(N276),.ZN(N287));
  INVX0 U162(.INP(N259),.ZN(N270));
  INVX0 U163(.INP(N293),.ZN(N304));
  INVX0 U164(.INP(N310),.ZN(N321));
  NOR2X0 U165(.IN1(n230),.IN2(n231),.QN(n229));
  NOR2X0 U166(.IN1(n217),.IN2(n218),.QN(n216));
  NOR2X0 U167(.IN1(n202),.IN2(n203),.QN(n201));
  NOR2X0 U168(.IN1(n191),.IN2(n192),.QN(n190));
  NOR2X0 U169(.IN1(n365),.IN2(opa_i[20:20]),.QN(n363));
  INVX0 U170(.INP(N243),.ZN(N253));
  NAND2X0 U171(.IN1(n418),.IN2(n92),.QN(n446));
  OA21X1 U172(.IN1(n297),.IN2(n298),.IN3(n145),.Q(s_div_zeros[3:3]));
  INVX0 U173(.INP(N344),.ZN(N355));
  INVX0 U174(.INP(N446),.ZN(N457));
  INVX0 U175(.INP(n362),.ZN(n376));
  INVX0 U176(.INP(N395),.ZN(N406));
  INVX0 U177(.INP(n258),.ZN(n108));
  INVX0 U178(.INP(n15),.ZN(n385));
  INVX0 U179(.INP(N514),.ZN(N525));
  INVX0 U180(.INP(N327),.ZN(N338));
  INVX0 U181(.INP(N1126),.ZN(N1137));
  INVX0 U182(.INP(N906),.ZN(N916));
  INVX0 U183(.INP(N1024),.ZN(N1035));
  NOR2X0 U184(.IN1(n252),.IN2(n253),.QN(n251));
  INVX0 U185(.INP(N548),.ZN(N559));
  OA21X1 U186(.IN1(n286),.IN2(n287),.IN3(n145),.Q(s_div_zeros[4:4]));
  INVX0 U187(.INP(N1080),.ZN(n63));
  INVX0 U188(.INP(N1131),.ZN(n60));
  NOR2X0 U189(.IN1(n276),.IN2(n277),.QN(n274));
  AND2X1 U190(.IN1(N938),.IN2(n386),.Q(n11));
  NOR2X0 U191(.IN1(n19),.IN2(n491),.QN(dvdnd_50_o[48:48]));
  INVX0 U192(.INP(n488),.ZN(n89));
  NOR2X0 U193(.IN1(n295),.IN2(n296),.QN(n294));
  NOR2X0 U194(.IN1(n334),.IN2(n335),.QN(n333));
  NOR2X0 U195(.IN1(n321),.IN2(n322),.QN(n320));
  NOR2X0 U196(.IN1(n306),.IN2(n307),.QN(n305));
  NOR2X0 U197(.IN1(n356),.IN2(n357),.QN(n355));
  INVX0 U198(.INP(N1211),.ZN(N1222));
  INVX0 U199(.INP(N429),.ZN(N440));
  INVX0 U200(.INP(N480),.ZN(N491));
  NAND2X0 U201(.IN1(n522),.IN2(n142),.QN(n550));
  INVX0 U202(.INP(n14),.ZN(n392));
  INVX0 U203(.INP(n551),.ZN(n135));
  INVX0 U204(.INP(n526),.ZN(n131));
  INVX0 U205(.INP(n544),.ZN(n132));
  NOR2X0 U206(.IN1(n17),.IN2(n595),.QN(dvsor_27_o[22:22]));
  INVX0 U437(.INP(n592),.ZN(n139));
  INVX0 U443(.INP(n411),.ZN(n72));
  INVX0 U444(.INP(n412),.ZN(n73));
  INVX0 U449(.INP(n413),.ZN(n74));
  INVX0 U454(.INP(n410),.ZN(n71));
  INVX0 U539(.INP(n408),.ZN(n70));
  INVX0 U540(.INP(n528),.ZN(n129));
  INVX0 U546(.INP(n525),.ZN(n127));
  INVX0 U547(.INP(N1130),.ZN(n65));
  INVX0 U584(.INP(N1127),.ZN(n154));
  INVX0 U585(.INP(N1128),.ZN(n150));
  INVX0 U586(.INP(N1129),.ZN(n146));
  INVX0 U587(.INP(opa_i[10:10]),.ZN(n39));
  INVX0 U588(.INP(N1096),.ZN(n67));
  INVX0 U589(.INP(N1095),.ZN(n148));
  INVX0 U590(.INP(N1110),.ZN(n373));
  INVX0 U591(.INP(N1111),.ZN(n151));
  INVX0 U592(.INP(N1113),.ZN(n66));
  INVX0 U593(.INP(N1112),.ZN(n147));
  INVX0 U594(.INP(N1097),.ZN(n62));
  INVX0 U595(.INP(N1114),.ZN(n61));
  INVX0 U596(.INP(N1093),.ZN(n374));
  INVX0 U597(.INP(N1094),.ZN(n152));
  INVX0 U598(.INP(N1079),.ZN(n68));
  INVX0 U599(.INP(N1076),.ZN(n375));
  INVX0 U600(.INP(N1077),.ZN(n153));
  INVX0 U601(.INP(N1078),.ZN(n149));
  INVX0 U602(.INP(opa_i[12:12]),.ZN(n117));
  INVX0 U603(.INP(n13),.ZN(n399));
  NAND2X0 U604(.IN1(n380),.IN2(n391),.QN(n318));
  NAND2X0 U605(.IN1(n381),.IN2(n390),.QN(n347));
  NAND2X0 U606(.IN1(n382),.IN2(n389),.QN(n345));
  NAND2X0 U607(.IN1(n384),.IN2(n387),.QN(n344));
  NAND2X0 U608(.IN1(n383),.IN2(n388),.QN(n346));
  NAND2X0 U609(.IN1(n386),.IN2(n385),.QN(n343));
  NAND2X0 U610(.IN1(n264),.IN2(N1024),.QN(n339));
  NAND2X0 U611(.IN1(n264),.IN2(N1026),.QN(n312));
  NAND2X0 U612(.IN1(n264),.IN2(N1025),.QN(n326));
  NOR2X0 U613(.IN1(n360),.IN2(n280),.QN(n282));
  INVX0 U614(.INP(opa_i[18:18]),.ZN(n48));
  NOR2X0 U615(.IN1(n358),.IN2(n359),.QN(n279));
  NAND2X1 U616(.IN1(n393),.IN2(n398),.QN(n275));
  NOR2X0 U617(.IN1(n351),.IN2(n14),.QN(n283));
  NOR2X0 U618(.IN1(n384),.IN2(n15),.QN(n262));
  NAND2X1 U619(.IN1(n351),.IN2(n395),.QN(n352));
  NAND2X0 U620(.IN1(n400),.IN2(n399),.QN(n358));
  NAND2X1 U621(.IN1(n359),.IN2(n402),.QN(n360));
  NAND2X1 U622(.IN1(n351),.IN2(n352),.QN(n272));
  NAND2X1 U623(.IN1(n353),.IN2(n354),.QN(n285));
  NAND2X1 U624(.IN1(n353),.IN2(n397),.QN(n354));
  NOR2X0 U625(.IN1(n257),.IN2(opa_i[20:20]),.QN(n205));
  INVX0 U626(.INP(opa_i[11:11]),.ZN(n41));
  NAND2X0 U627(.IN1(n205),.IN2(n110),.QN(n206));
  NOR2X0 U628(.IN1(n256),.IN2(n176),.QN(n178));
  INVX0 U629(.INP(opa_i[8:8]),.ZN(n36));
  INVX0 U630(.INP(opa_i[3:3]),.ZN(n29));
  INVX0 U631(.INP(N192),.ZN(\add_116/B[0] ));
  INVX0 U632(.INP(opa_i[1:1]),.ZN(n26));
  INVX0 U633(.INP(N199),.ZN(\add_117/B[0] ));
  NAND2X1 U634(.IN1(n1),.IN2(n9),.QN(n12));
  NAND2X0 U635(.IN1(n366),.IN2(n367),.QN(N192));
  NOR2X0 U636(.IN1(N192),.IN2(opa_i[22:22]),.QN(n220));
  INVX0 U637(.INP(N229),.ZN(N238));
  NBUFFX2 U638(.INP(opb_i[18:18]),.Z(n15));
  INVX0 U639(.INP(N1092),.ZN(N1103));
  INVX0 U640(.INP(N1177),.ZN(N1188));
  INVX0 U641(.INP(N1160),.ZN(N1171));
  INVX0 U642(.INP(N939),.ZN(N950));
  INVX0 U643(.INP(N990),.ZN(N1001));
  INVX0 U644(.INP(N922),.ZN(N933));
  INVX0 U645(.INP(N973),.ZN(N984));
  INVX0 U646(.INP(N1194),.ZN(N1205));
  INVX0 U647(.INP(N1075),.ZN(N1086));
  INVX0 U648(.INP(N1109),.ZN(N1120));
  INVX0 U649(.INP(N1143),.ZN(N1154));
  INVX0 U650(.INP(N956),.ZN(N967));
  INVX0 U651(.INP(N1007),.ZN(N1018));
  INVX0 U652(.INP(N1058),.ZN(N1069));
  INVX0 U653(.INP(N1041),.ZN(N1052));
  NBUFFX2 U654(.INP(opb_i[11:11]),.Z(n14));
  NAND2X0 U655(.IN1(opa_i[0:0]),.IN2(n21),.QN(n409));
  NAND2X0 U656(.IN1(opb_i[0:0]),.IN2(n23),.QN(n513));
  INVX0 U657(.INP(n516),.ZN(n123));
  INVX0 U658(.INP(n517),.ZN(n124));
  INVX0 U659(.INP(n515),.ZN(n122));
  INVX0 U660(.INP(n514),.ZN(n121));
  INVX0 U661(.INP(n512),.ZN(n120));
  NAND2X0 U662(.IN1(n371),.IN2(n372),.QN(N199));
  NBUFFX2 U663(.INP(opb_i[5:5]),.Z(n13));
  INVX0 U664(.INP(opa_i[19:19]),.ZN(n110));
  NOR2X0 U665(.IN1(N199),.IN2(opb_i[22:22]),.QN(n324));
  NOR2X0 U666(.IN1(n370),.IN2(opb_i[20:20]),.QN(n368));
  INVX0 U667(.INP(N892),.ZN(N901));
  NOR2X0 U668(.IN1(opb_i[10:10]),.IN2(n14),.QN(n351));
  NOR2X0 U669(.IN1(n352),.IN2(opb_i[8:8]),.QN(n353));
  NOR2X0 U670(.IN1(n358),.IN2(opb_i[3:3]),.QN(n359));
  INVX0 U671(.INP(opb_i[16:16]),.ZN(n387));
  INVX0 U672(.INP(opa_i[21:21]),.ZN(n109));
  INVX0 U673(.INP(opb_i[21:21]),.ZN(n377));
  INVX0 U674(.INP(opb_i[17:17]),.ZN(n386));
  INVX0 U675(.INP(opb_i[15:15]),.ZN(n388));
  INVX0 U676(.INP(opb_i[14:14]),.ZN(n389));
  INVX0 U677(.INP(opb_i[19:19]),.ZN(n378));
  INVX0 U678(.INP(opb_i[12:12]),.ZN(n391));
  INVX0 U679(.INP(opb_i[13:13]),.ZN(n390));
  INVX0 U680(.INP(opb_i[6:6]),.ZN(n398));
  INVX0 U681(.INP(opb_i[7:7]),.ZN(n397));
  INVX0 U682(.INP(opb_i[9:9]),.ZN(n395));
  INVX0 U683(.INP(opb_i[10:10]),.ZN(n394));
  INVX0 U684(.INP(opb_i[8:8]),.ZN(n396));
  INVX0 U685(.INP(opb_i[4:4]),.ZN(n400));
  NOR2X0 U686(.IN1(n361),.IN2(opb_i[20:20]),.QN(n309));
  INVX0 U687(.INP(opb_i[3:3]),.ZN(n401));
  INVX0 U688(.INP(opb_i[1:1]),.ZN(n403));
  INVX0 U689(.INP(opb_i[2:2]),.ZN(n402));
  INVX0 U690(.INP(n26),.ZN(n25));
  INVX0 U691(.INP(opa_i[2:2]),.ZN(n27));
  INVX0 U692(.INP(n29),.ZN(n28));
  INVX0 U693(.INP(opa_i[4:4]),.ZN(n30));
  INVX0 U694(.INP(n32),.ZN(n31));
  INVX0 U695(.INP(opa_i[5:5]),.ZN(n32));
  INVX0 U696(.INP(opa_i[6:6]),.ZN(n33));
  INVX0 U697(.INP(opa_i[7:7]),.ZN(n34));
  INVX0 U698(.INP(n36),.ZN(n35));
  INVX0 U699(.INP(opa_i[9:9]),.ZN(n37));
  INVX0 U700(.INP(n39),.ZN(n38));
  INVX0 U701(.INP(n41),.ZN(n40));
  INVX0 U702(.INP(opa_i[13:13]),.ZN(n42));
  INVX0 U703(.INP(opa_i[14:14]),.ZN(n43));
  INVX0 U704(.INP(opa_i[15:15]),.ZN(n44));
  INVX0 U705(.INP(opa_i[16:16]),.ZN(n45));
  INVX0 U706(.INP(opa_i[17:17]),.ZN(n46));
  INVX0 U707(.INP(n48),.ZN(n47));
  XOR2X1 U708(.IN1(n9),.IN2(n1),.Q(N1562));
  AND2X1 U709(.IN1(\add_117/carry[7] ),.IN2(opb_i[30:30]),.Q(N1543));
  XOR2X1 U710(.IN1(opb_i[30:30]),.IN2(\add_117/carry[7] ),.Q(N1542));
  AND2X1 U711(.IN1(\add_117/carry[6] ),.IN2(opb_i[29:29]),.Q(\add_117/carry[7] ));
  XOR2X1 U712(.IN1(opb_i[29:29]),.IN2(\add_117/carry[6] ),.Q(N1541));
  AND2X1 U713(.IN1(\add_117/carry[5] ),.IN2(opb_i[28:28]),.Q(\add_117/carry[6] ));
  XOR2X1 U714(.IN1(opb_i[28:28]),.IN2(\add_117/carry[5] ),.Q(N1540));
  AND2X1 U715(.IN1(\add_117/carry[4] ),.IN2(opb_i[27:27]),.Q(\add_117/carry[5] ));
  XOR2X1 U716(.IN1(opb_i[27:27]),.IN2(\add_117/carry[4] ),.Q(N1539));
  AND2X1 U717(.IN1(\add_117/carry[3] ),.IN2(opb_i[26:26]),.Q(\add_117/carry[4] ));
  XOR2X1 U718(.IN1(opb_i[26:26]),.IN2(\add_117/carry[3] ),.Q(N1538));
  AND2X1 U719(.IN1(\add_117/carry[2] ),.IN2(opb_i[25:25]),.Q(\add_117/carry[3] ));
  XOR2X1 U720(.IN1(opb_i[25:25]),.IN2(\add_117/carry[2] ),.Q(N1537));
  AND2X1 U721(.IN1(\add_117/carry[1] ),.IN2(opb_i[24:24]),.Q(\add_117/carry[2] ));
  XOR2X1 U722(.IN1(opb_i[24:24]),.IN2(\add_117/carry[1] ),.Q(N1536));
  AND2X1 U723(.IN1(\add_117/B[0] ),.IN2(opb_i[23:23]),.Q(\add_117/carry[1] ));
  XOR2X1 U724(.IN1(opb_i[23:23]),.IN2(\add_117/B[0] ),.Q(N1535));
  AND2X1 U725(.IN1(\add_116/carry[7] ),.IN2(opa_i[30:30]),.Q(N1534));
  XOR2X1 U726(.IN1(opa_i[30:30]),.IN2(\add_116/carry[7] ),.Q(N1533));
  AND2X1 U727(.IN1(\add_116/carry[6] ),.IN2(opa_i[29:29]),.Q(\add_116/carry[7] ));
  XOR2X1 U728(.IN1(opa_i[29:29]),.IN2(\add_116/carry[6] ),.Q(N1532));
  AND2X1 U729(.IN1(\add_116/carry[5] ),.IN2(opa_i[28:28]),.Q(\add_116/carry[6] ));
  XOR2X1 U730(.IN1(opa_i[28:28]),.IN2(\add_116/carry[5] ),.Q(N1531));
  AND2X1 U731(.IN1(\add_116/carry[4] ),.IN2(opa_i[27:27]),.Q(\add_116/carry[5] ));
  XOR2X1 U732(.IN1(opa_i[27:27]),.IN2(\add_116/carry[4] ),.Q(N1530));
  AND2X1 U733(.IN1(\add_116/carry[3] ),.IN2(opa_i[26:26]),.Q(\add_116/carry[4] ));
  XOR2X1 U734(.IN1(opa_i[26:26]),.IN2(\add_116/carry[3] ),.Q(N1529));
  AND2X1 U735(.IN1(\add_116/carry[2] ),.IN2(opa_i[25:25]),.Q(\add_116/carry[3] ));
  XOR2X1 U736(.IN1(opa_i[25:25]),.IN2(\add_116/carry[2] ),.Q(N1528));
  AND2X1 U737(.IN1(\add_116/carry[1] ),.IN2(opa_i[24:24]),.Q(\add_116/carry[2] ));
  XOR2X1 U738(.IN1(opa_i[24:24]),.IN2(\add_116/carry[1] ),.Q(N1527));
  AND2X1 U739(.IN1(\add_116/B[0] ),.IN2(opa_i[23:23]),.Q(\add_116/carry[1] ));
  XOR2X1 U740(.IN1(opa_i[23:23]),.IN2(\add_116/B[0] ),.Q(N1526));
  XOR2X1 U741(.IN1(\add_90_I8_L14036_C103/carry[5] ),.IN2(n10),.Q(N292));
  XOR2X1 U742(.IN1(\add_90_I9_L14036_C103/carry[5] ),.IN2(N298),.Q(N309));
  XOR2X1 U743(.IN1(\add_90_I10_L14036_C103/carry[5] ),.IN2(N315),.Q(N326));
  XOR2X1 U744(.IN1(\add_90_I11_L14036_C103/carry[5] ),.IN2(N332),.Q(N343));
  XOR2X1 U745(.IN1(\add_90_I12_L14036_C103/carry[5] ),.IN2(N349),.Q(N360));
  XOR2X1 U746(.IN1(\add_90_I13_L14036_C103/carry[5] ),.IN2(N366),.Q(N377));
  XOR2X1 U747(.IN1(\add_90_I14_L14036_C103/carry[5] ),.IN2(N383),.Q(N394));
  XOR2X1 U748(.IN1(\add_90_I15_L14036_C103/carry[5] ),.IN2(N400),.Q(N411));
  XOR2X1 U749(.IN1(\add_90_I16_L14036_C103/carry[5] ),.IN2(N417),.Q(N428));
  XOR2X1 U750(.IN1(\add_90_I17_L14036_C103/carry[5] ),.IN2(N434),.Q(N445));
  XOR2X1 U751(.IN1(\add_90_I18_L14036_C103/carry[5] ),.IN2(N451),.Q(N462));
  XOR2X1 U752(.IN1(\add_90_I19_L14036_C103/carry[5] ),.IN2(N468),.Q(N479));
  XOR2X1 U753(.IN1(\add_90_I20_L14036_C103/carry[5] ),.IN2(N485),.Q(N496));
  XOR2X1 U754(.IN1(\add_90_I21_L14036_C103/carry[5] ),.IN2(N502),.Q(N513));
  XOR2X1 U755(.IN1(\add_90_I22_L14036_C103/carry[5] ),.IN2(N519),.Q(N530));
  XOR2X1 U756(.IN1(\add_90_I23_L14036_C103/carry[5] ),.IN2(N536),.Q(N547));
  XOR2X1 U757(.IN1(\add_90_I24_L14036_C103/carry[5] ),.IN2(N553),.Q(N564));
  XOR2X1 U758(.IN1(\add_90_I8_L14036_C104/carry[5] ),.IN2(n11),.Q(N955));
  XOR2X1 U759(.IN1(\add_90_I9_L14036_C104/carry[5] ),.IN2(N961),.Q(N972));
  XOR2X1 U760(.IN1(\add_90_I10_L14036_C104/carry[5] ),.IN2(N978),.Q(N989));
  XOR2X1 U761(.IN1(\add_90_I11_L14036_C104/carry[5] ),.IN2(N995),.Q(N1006));
  XOR2X1 U762(.IN1(\add_90_I12_L14036_C104/carry[5] ),.IN2(N1012),.Q(N1023));
  XOR2X1 U763(.IN1(\add_90_I13_L14036_C104/carry[5] ),.IN2(N1029),.Q(N1040));
  XOR2X1 U764(.IN1(\add_90_I14_L14036_C104/carry[5] ),.IN2(N1046),.Q(N1057));
  XOR2X1 U765(.IN1(\add_90_I15_L14036_C104/carry[5] ),.IN2(N1063),.Q(N1074));
  XOR2X1 U766(.IN1(\add_90_I16_L14036_C104/carry[5] ),.IN2(N1080),.Q(N1091));
  XOR2X1 U767(.IN1(\add_90_I17_L14036_C104/carry[5] ),.IN2(N1097),.Q(N1108));
  XOR2X1 U768(.IN1(\add_90_I18_L14036_C104/carry[5] ),.IN2(N1114),.Q(N1125));
  XOR2X1 U769(.IN1(\add_90_I19_L14036_C104/carry[5] ),.IN2(N1131),.Q(N1142));
  XOR2X1 U770(.IN1(\add_90_I20_L14036_C104/carry[5] ),.IN2(N1148),.Q(N1159));
  XOR2X1 U771(.IN1(\add_90_I21_L14036_C104/carry[5] ),.IN2(N1165),.Q(N1176));
  XOR2X1 U772(.IN1(\add_90_I22_L14036_C104/carry[5] ),.IN2(N1182),.Q(N1193));
  XOR2X1 U773(.IN1(\add_90_I23_L14036_C104/carry[5] ),.IN2(N1199),.Q(N1210));
  XOR2X1 U774(.IN1(\add_90_I24_L14036_C104/carry[5] ),.IN2(N1216),.Q(N1227));
  AND2X1 U775(.IN1(N257),.IN2(n48),.Q(N263));
  AND2X1 U776(.IN1(N920),.IN2(n385),.Q(N926));
  OR2X1 U781(.IN1(n409),.IN2(s_dvd_zeros[1:1]),.Q(n416));
  NOR3X0 U782(.IN1(n444),.IN2(n19),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[26:26]));
  MUX21X1 U783(.IN1(n25),.IN2(opa_i[2:2]),.S(n22),.Q(n408));
  MUX21X1 U784(.IN1(n409),.IN2(n70),.S(n92),.Q(n428));
  OR2X1 U785(.IN1(n428),.IN2(s_dvd_zeros[2:2]),.Q(n452));
  MUX21X1 U786(.IN1(n28),.IN2(opa_i[4:4]),.S(n22),.Q(n410));
  MUX21X1 U787(.IN1(n31),.IN2(opa_i[6:6]),.S(n22),.Q(n411));
  MUX21X1 U788(.IN1(n71),.IN2(n72),.S(n92),.Q(n427));
  MUX21X1 U789(.IN1(opa_i[7:7]),.IN2(n35),.S(n22),.Q(n412));
  MUX21X1 U790(.IN1(opa_i[9:9]),.IN2(n38),.S(n22),.Q(n413));
  MUX21X1 U791(.IN1(n73),.IN2(n74),.S(n92),.Q(n430));
  MUX21X1 U792(.IN1(n427),.IN2(n430),.S(n93),.Q(n456));
  MUX21X1 U793(.IN1(n452),.IN2(n456),.S(n94),.Q(n414));
  NOR3X0 U794(.IN1(n414),.IN2(n20),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[36:36]));
  MUX21X1 U795(.IN1(opa_i[0:0]),.IN2(n25),.S(n22),.Q(n418));
  MUX21X1 U796(.IN1(opa_i[2:2]),.IN2(n28),.S(n22),.Q(n420));
  MUX21X1 U797(.IN1(n418),.IN2(n420),.S(n92),.Q(n433));
  MUX21X1 U798(.IN1(opa_i[4:4]),.IN2(n31),.S(n22),.Q(n419));
  MUX21X1 U799(.IN1(opa_i[6:6]),.IN2(opa_i[7:7]),.S(n22),.Q(n423));
  MUX21X1 U800(.IN1(n419),.IN2(n423),.S(n92),.Q(n432));
  MUX21X1 U801(.IN1(n35),.IN2(opa_i[9:9]),.S(n22),.Q(n422));
  MUX21X1 U802(.IN1(n39),.IN2(n41),.S(n22),.Q(n425));
  MUX21X1 U803(.IN1(n81),.IN2(n425),.S(n92),.Q(n436));
  MUX21X1 U804(.IN1(n78),.IN2(n436),.S(n93),.Q(n463));
  MUX21X1 U805(.IN1(n459),.IN2(n463),.S(n94),.Q(n415));
  NOR3X0 U806(.IN1(n415),.IN2(n19),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[37:37]));
  MUX21X1 U807(.IN1(n70),.IN2(n71),.S(n92),.Q(n439));
  MUX21X1 U808(.IN1(n416),.IN2(n439),.S(n93),.Q(n467));
  MUX21X1 U809(.IN1(n72),.IN2(n73),.S(n92),.Q(n438));
  MUX21X1 U810(.IN1(n41),.IN2(n117),.S(n22),.Q(n429));
  MUX21X1 U811(.IN1(n74),.IN2(n429),.S(n92),.Q(n441));
  MUX21X1 U812(.IN1(n438),.IN2(n441),.S(n93),.Q(n472));
  MUX21X1 U813(.IN1(n467),.IN2(n472),.S(n94),.Q(n417));
  NOR3X0 U814(.IN1(n417),.IN2(n20),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[38:38]));
  MUX21X1 U815(.IN1(n420),.IN2(n419),.S(n92),.Q(n421));
  MUX21X1 U816(.IN1(n446),.IN2(n77),.S(n93),.Q(n475));
  MUX21X1 U817(.IN1(n423),.IN2(n422),.S(n92),.Q(n424));
  MUX21X1 U818(.IN1(n117),.IN2(n42),.S(n21),.Q(n435));
  MUX21X1 U819(.IN1(n425),.IN2(n435),.S(n92),.Q(n448));
  MUX21X1 U820(.IN1(n79),.IN2(n448),.S(n93),.Q(n480));
  MUX21X1 U821(.IN1(n475),.IN2(n480),.S(n94),.Q(n426));
  NOR3X0 U822(.IN1(n426),.IN2(s_dvd_zeros[5:5]),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[39:39]));
  MUX21X1 U823(.IN1(n428),.IN2(n427),.S(n93),.Q(n483));
  MUX21X1 U824(.IN1(opa_i[13:13]),.IN2(opa_i[14:14]),.S(n21),.Q(n440));
  MUX21X1 U825(.IN1(n429),.IN2(n82),.S(n92),.Q(n454));
  MUX21X1 U826(.IN1(n430),.IN2(n454),.S(n93),.Q(n489));
  MUX21X1 U827(.IN1(n483),.IN2(n489),.S(n94),.Q(n431));
  NOR3X0 U828(.IN1(s_dvd_zeros[4:4]),.IN2(n19),.IN3(n431),.QN(dvdnd_50_o[40:40]));
  MUX21X1 U829(.IN1(n433),.IN2(n432),.S(n93),.Q(n434));
  MUX21X1 U830(.IN1(opa_i[14:14]),.IN2(opa_i[15:15]),.S(n21),.Q(n447));
  MUX21X1 U831(.IN1(n435),.IN2(n85),.S(n92),.Q(n461));
  MUX21X1 U832(.IN1(n436),.IN2(n461),.S(n93),.Q(n492));
  MUX21X1 U833(.IN1(n75),.IN2(n492),.S(n94),.Q(n437));
  NOR3X0 U834(.IN1(s_dvd_zeros[4:4]),.IN2(n20),.IN3(n437),.QN(dvdnd_50_o[41:41]));
  MUX21X1 U835(.IN1(n439),.IN2(n438),.S(n93),.Q(n506));
  MUX21X1 U836(.IN1(opa_i[15:15]),.IN2(opa_i[16:16]),.S(n21),.Q(n453));
  MUX21X1 U837(.IN1(n440),.IN2(n453),.S(n92),.Q(n470));
  MUX21X1 U838(.IN1(n441),.IN2(n83),.S(n93),.Q(n442));
  MUX21X1 U839(.IN1(n506),.IN2(n442),.S(n94),.Q(n443));
  MUX21X1 U840(.IN1(n444),.IN2(n443),.S(n54),.Q(n445));
  MUX21X1 U841(.IN1(n77),.IN2(n79),.S(n93),.Q(n510));
  MUX21X1 U842(.IN1(opa_i[16:16]),.IN2(opa_i[17:17]),.S(n21),.Q(n460));
  MUX21X1 U843(.IN1(n447),.IN2(n460),.S(n92),.Q(n478));
  MUX21X1 U844(.IN1(n448),.IN2(n86),.S(n93),.Q(n449));
  MUX21X1 U845(.IN1(n510),.IN2(n449),.S(n94),.Q(n450));
  MUX21X1 U846(.IN1(n466),.IN2(n450),.S(n54),.Q(n451));
  OR2X1 U847(.IN1(n452),.IN2(s_dvd_zeros[3:3]),.Q(n500));
  MUX21X1 U848(.IN1(opa_i[17:17]),.IN2(n47),.S(n21),.Q(n468));
  MUX21X1 U849(.IN1(n453),.IN2(n468),.S(n92),.Q(n487));
  MUX21X1 U850(.IN1(n454),.IN2(n88),.S(n93),.Q(n455));
  MUX21X1 U851(.IN1(n456),.IN2(n455),.S(n94),.Q(n457));
  MUX21X1 U852(.IN1(n500),.IN2(n457),.S(n54),.Q(n458));
  OR2X1 U853(.IN1(n459),.IN2(s_dvd_zeros[3:3]),.Q(n501));
  MUX21X1 U854(.IN1(n47),.IN2(opa_i[19:19]),.S(n21),.Q(n476));
  MUX21X1 U855(.IN1(n460),.IN2(n476),.S(n92),.Q(n496));
  MUX21X1 U856(.IN1(n461),.IN2(n90),.S(n93),.Q(n462));
  MUX21X1 U857(.IN1(n463),.IN2(n462),.S(n94),.Q(n464));
  MUX21X1 U858(.IN1(n501),.IN2(n464),.S(n54),.Q(n465));
  NOR3X0 U859(.IN1(n466),.IN2(s_dvd_zeros[5:5]),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[27:27]));
  OR2X1 U860(.IN1(n467),.IN2(s_dvd_zeros[3:3]),.Q(n502));
  MUX21X1 U861(.IN1(opa_i[19:19]),.IN2(opa_i[20:20]),.S(n21),.Q(n485));
  MUX21X1 U862(.IN1(n468),.IN2(n485),.S(n92),.Q(n469));
  MUX21X1 U863(.IN1(n470),.IN2(n469),.S(n93),.Q(n471));
  MUX21X1 U864(.IN1(n472),.IN2(n84),.S(n94),.Q(n473));
  MUX21X1 U865(.IN1(n502),.IN2(n473),.S(n54),.Q(n474));
  OR2X1 U866(.IN1(n475),.IN2(s_dvd_zeros[3:3]),.Q(n503));
  MUX21X1 U867(.IN1(opa_i[20:20]),.IN2(opa_i[21:21]),.S(n21),.Q(n494));
  MUX21X1 U868(.IN1(n476),.IN2(n494),.S(n92),.Q(n477));
  MUX21X1 U869(.IN1(n478),.IN2(n477),.S(n93),.Q(n479));
  MUX21X1 U870(.IN1(n480),.IN2(n87),.S(n94),.Q(n481));
  MUX21X1 U871(.IN1(n503),.IN2(n481),.S(n54),.Q(n482));
  OR2X1 U872(.IN1(n483),.IN2(s_dvd_zeros[3:3]),.Q(n504));
  MUX21X1 U873(.IN1(opa_i[21:21]),.IN2(opa_i[22:22]),.S(n21),.Q(n484));
  MUX21X1 U874(.IN1(n485),.IN2(n484),.S(n92),.Q(n486));
  MUX21X1 U875(.IN1(n487),.IN2(n486),.S(n93),.Q(n488));
  MUX21X1 U876(.IN1(n489),.IN2(n89),.S(n94),.Q(n490));
  MUX21X1 U877(.IN1(n504),.IN2(n490),.S(n54),.Q(n491));
  MUX21X1 U878(.IN1(opa_i[22:22]),.IN2(N192),.S(n21),.Q(n493));
  MUX21X1 U879(.IN1(n494),.IN2(n493),.S(n92),.Q(n495));
  MUX21X1 U880(.IN1(n496),.IN2(n495),.S(n93),.Q(n497));
  MUX21X1 U881(.IN1(n80),.IN2(n497),.S(n94),.Q(n498));
  MUX21X1 U882(.IN1(n505),.IN2(n498),.S(n54),.Q(n499));
  AND2X1 U883(.IN1(n499),.IN2(n49),.Q(dvdnd_50_o[49:49]));
  NOR3X0 U884(.IN1(s_dvd_zeros[4:4]),.IN2(n19),.IN3(n500),.QN(dvdnd_50_o[28:28]));
  NOR3X0 U885(.IN1(s_dvd_zeros[4:4]),.IN2(n20),.IN3(n501),.QN(dvdnd_50_o[29:29]));
  NOR3X0 U886(.IN1(s_dvd_zeros[4:4]),.IN2(s_dvd_zeros[5:5]),.IN3(n502),.QN(dvdnd_50_o[30:30]));
  NOR3X0 U887(.IN1(n503),.IN2(n19),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[31:31]));
  NOR3X0 U888(.IN1(n504),.IN2(n20),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[32:32]));
  AND3X1 U889(.IN1(n505),.IN2(n49),.IN3(n54),.Q(dvdnd_50_o[33:33]));
  MUX21X1 U890(.IN1(n507),.IN2(n69),.S(n94),.Q(n508));
  AND3X1 U891(.IN1(n54),.IN2(n49),.IN3(n508),.Q(dvdnd_50_o[34:34]));
  MUX21X1 U892(.IN1(n76),.IN2(n510),.S(n94),.Q(n511));
  NOR3X0 U893(.IN1(n511),.IN2(s_dvd_zeros[5:5]),.IN3(s_dvd_zeros[4:4]),.QN(dvdnd_50_o[35:35]));
  OR2X1 U894(.IN1(n513),.IN2(s_div_zeros[1:1]),.Q(n520));
  NOR3X0 U895(.IN1(n548),.IN2(n17),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[0:0]));
  MUX21X1 U896(.IN1(opb_i[1:1]),.IN2(opb_i[2:2]),.S(n24),.Q(n512));
  MUX21X1 U897(.IN1(n513),.IN2(n120),.S(n142),.Q(n532));
  OR2X1 U898(.IN1(n532),.IN2(s_div_zeros[2:2]),.Q(n556));
  MUX21X1 U899(.IN1(opb_i[3:3]),.IN2(opb_i[4:4]),.S(n24),.Q(n514));
  MUX21X1 U900(.IN1(n13),.IN2(opb_i[6:6]),.S(n24),.Q(n515));
  MUX21X1 U901(.IN1(n121),.IN2(n122),.S(n142),.Q(n531));
  MUX21X1 U902(.IN1(opb_i[7:7]),.IN2(opb_i[8:8]),.S(n24),.Q(n516));
  MUX21X1 U903(.IN1(opb_i[9:9]),.IN2(opb_i[10:10]),.S(n24),.Q(n517));
  MUX21X1 U904(.IN1(n123),.IN2(n124),.S(n142),.Q(n534));
  MUX21X1 U905(.IN1(n531),.IN2(n534),.S(n143),.Q(n560));
  MUX21X1 U906(.IN1(n556),.IN2(n560),.S(n144),.Q(n518));
  NOR3X0 U907(.IN1(n518),.IN2(n18),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[10:10]));
  MUX21X1 U908(.IN1(opb_i[0:0]),.IN2(opb_i[1:1]),.S(n24),.Q(n522));
  MUX21X1 U909(.IN1(opb_i[2:2]),.IN2(opb_i[3:3]),.S(n24),.Q(n524));
  MUX21X1 U910(.IN1(n522),.IN2(n524),.S(n142),.Q(n537));
  MUX21X1 U911(.IN1(opb_i[4:4]),.IN2(n13),.S(n24),.Q(n523));
  MUX21X1 U912(.IN1(opb_i[6:6]),.IN2(opb_i[7:7]),.S(n24),.Q(n527));
  MUX21X1 U913(.IN1(n523),.IN2(n527),.S(n142),.Q(n536));
  MUX21X1 U914(.IN1(opb_i[8:8]),.IN2(opb_i[9:9]),.S(n24),.Q(n526));
  MUX21X1 U915(.IN1(n394),.IN2(n392),.S(n24),.Q(n529));
  MUX21X1 U916(.IN1(n131),.IN2(n529),.S(n142),.Q(n540));
  MUX21X1 U917(.IN1(n128),.IN2(n540),.S(n143),.Q(n567));
  MUX21X1 U918(.IN1(n563),.IN2(n567),.S(n144),.Q(n519));
  NOR3X0 U919(.IN1(n519),.IN2(n17),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[11:11]));
  MUX21X1 U920(.IN1(n120),.IN2(n121),.S(n142),.Q(n543));
  MUX21X1 U921(.IN1(n520),.IN2(n543),.S(n143),.Q(n571));
  MUX21X1 U922(.IN1(n122),.IN2(n123),.S(n142),.Q(n542));
  MUX21X1 U923(.IN1(n392),.IN2(n391),.S(n24),.Q(n533));
  MUX21X1 U924(.IN1(n124),.IN2(n533),.S(n142),.Q(n545));
  MUX21X1 U925(.IN1(n542),.IN2(n545),.S(n143),.Q(n576));
  MUX21X1 U926(.IN1(n571),.IN2(n576),.S(n144),.Q(n521));
  NOR3X0 U927(.IN1(n521),.IN2(n18),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[12:12]));
  MUX21X1 U928(.IN1(n524),.IN2(n523),.S(n142),.Q(n525));
  MUX21X1 U929(.IN1(n550),.IN2(n127),.S(n143),.Q(n579));
  MUX21X1 U930(.IN1(n527),.IN2(n526),.S(n142),.Q(n528));
  MUX21X1 U931(.IN1(n391),.IN2(n390),.S(n23),.Q(n539));
  MUX21X1 U932(.IN1(n529),.IN2(n539),.S(n142),.Q(n552));
  MUX21X1 U933(.IN1(n129),.IN2(n552),.S(n143),.Q(n584));
  MUX21X1 U934(.IN1(n579),.IN2(n584),.S(n144),.Q(n530));
  NOR3X0 U935(.IN1(n530),.IN2(s_div_zeros[5:5]),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[13:13]));
  MUX21X1 U936(.IN1(n532),.IN2(n531),.S(n143),.Q(n587));
  MUX21X1 U937(.IN1(opb_i[13:13]),.IN2(opb_i[14:14]),.S(n23),.Q(n544));
  MUX21X1 U938(.IN1(n533),.IN2(n132),.S(n142),.Q(n558));
  MUX21X1 U939(.IN1(n534),.IN2(n558),.S(n143),.Q(n593));
  MUX21X1 U940(.IN1(n587),.IN2(n593),.S(n144),.Q(n535));
  NOR3X0 U941(.IN1(s_div_zeros[4:4]),.IN2(n17),.IN3(n535),.QN(dvsor_27_o[14:14]));
  MUX21X1 U942(.IN1(n537),.IN2(n536),.S(n143),.Q(n538));
  MUX21X1 U943(.IN1(opb_i[14:14]),.IN2(opb_i[15:15]),.S(n23),.Q(n551));
  MUX21X1 U944(.IN1(n539),.IN2(n135),.S(n142),.Q(n565));
  MUX21X1 U945(.IN1(n540),.IN2(n565),.S(n143),.Q(n596));
  MUX21X1 U946(.IN1(n125),.IN2(n596),.S(n144),.Q(n541));
  NOR3X0 U947(.IN1(s_div_zeros[4:4]),.IN2(n18),.IN3(n541),.QN(dvsor_27_o[15:15]));
  MUX21X1 U948(.IN1(n543),.IN2(n542),.S(n143),.Q(n610));
  MUX21X1 U949(.IN1(opb_i[15:15]),.IN2(opb_i[16:16]),.S(n23),.Q(n557));
  MUX21X1 U950(.IN1(n544),.IN2(n557),.S(n142),.Q(n574));
  MUX21X1 U951(.IN1(n545),.IN2(n133),.S(n143),.Q(n546));
  MUX21X1 U952(.IN1(n610),.IN2(n546),.S(n144),.Q(n547));
  MUX21X1 U953(.IN1(n548),.IN2(n547),.S(n64),.Q(n549));
  MUX21X1 U954(.IN1(n127),.IN2(n129),.S(n143),.Q(n614));
  MUX21X1 U955(.IN1(opb_i[16:16]),.IN2(opb_i[17:17]),.S(n23),.Q(n564));
  MUX21X1 U956(.IN1(n551),.IN2(n564),.S(n142),.Q(n582));
  MUX21X1 U957(.IN1(n552),.IN2(n136),.S(n143),.Q(n553));
  MUX21X1 U958(.IN1(n614),.IN2(n553),.S(n144),.Q(n554));
  MUX21X1 U959(.IN1(n570),.IN2(n554),.S(n64),.Q(n555));
  OR2X1 U960(.IN1(n556),.IN2(s_div_zeros[3:3]),.Q(n604));
  MUX21X1 U961(.IN1(opb_i[17:17]),.IN2(n16),.S(n23),.Q(n572));
  MUX21X1 U962(.IN1(n557),.IN2(n572),.S(n142),.Q(n591));
  MUX21X1 U963(.IN1(n558),.IN2(n138),.S(n143),.Q(n559));
  MUX21X1 U964(.IN1(n560),.IN2(n559),.S(n144),.Q(n561));
  MUX21X1 U965(.IN1(n604),.IN2(n561),.S(n64),.Q(n562));
  OR2X1 U966(.IN1(n563),.IN2(s_div_zeros[3:3]),.Q(n605));
  MUX21X1 U967(.IN1(n16),.IN2(opb_i[19:19]),.S(n23),.Q(n580));
  MUX21X1 U968(.IN1(n564),.IN2(n580),.S(n142),.Q(n600));
  MUX21X1 U969(.IN1(n565),.IN2(n140),.S(n143),.Q(n566));
  MUX21X1 U970(.IN1(n567),.IN2(n566),.S(n144),.Q(n568));
  MUX21X1 U971(.IN1(n605),.IN2(n568),.S(n64),.Q(n569));
  NOR3X0 U972(.IN1(n570),.IN2(s_div_zeros[5:5]),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[1:1]));
  OR2X1 U973(.IN1(n571),.IN2(s_div_zeros[3:3]),.Q(n606));
  MUX21X1 U974(.IN1(opb_i[19:19]),.IN2(opb_i[20:20]),.S(n23),.Q(n589));
  MUX21X1 U975(.IN1(n572),.IN2(n589),.S(n142),.Q(n573));
  MUX21X1 U976(.IN1(n574),.IN2(n573),.S(n143),.Q(n575));
  MUX21X1 U977(.IN1(n576),.IN2(n134),.S(n144),.Q(n577));
  MUX21X1 U978(.IN1(n606),.IN2(n577),.S(n64),.Q(n578));
  OR2X1 U979(.IN1(n579),.IN2(s_div_zeros[3:3]),.Q(n607));
  MUX21X1 U980(.IN1(opb_i[20:20]),.IN2(opb_i[21:21]),.S(n23),.Q(n598));
  MUX21X1 U981(.IN1(n580),.IN2(n598),.S(n142),.Q(n581));
  MUX21X1 U982(.IN1(n582),.IN2(n581),.S(n143),.Q(n583));
  MUX21X1 U983(.IN1(n584),.IN2(n137),.S(n144),.Q(n585));
  MUX21X1 U984(.IN1(n607),.IN2(n585),.S(n64),.Q(n586));
  OR2X1 U985(.IN1(n587),.IN2(s_div_zeros[3:3]),.Q(n608));
  MUX21X1 U986(.IN1(opb_i[21:21]),.IN2(opb_i[22:22]),.S(n23),.Q(n588));
  MUX21X1 U987(.IN1(n589),.IN2(n588),.S(n142),.Q(n590));
  MUX21X1 U988(.IN1(n591),.IN2(n590),.S(n143),.Q(n592));
  MUX21X1 U989(.IN1(n593),.IN2(n139),.S(n144),.Q(n594));
  MUX21X1 U990(.IN1(n608),.IN2(n594),.S(n64),.Q(n595));
  MUX21X1 U991(.IN1(opb_i[22:22]),.IN2(N199),.S(n23),.Q(n597));
  MUX21X1 U992(.IN1(n598),.IN2(n597),.S(n142),.Q(n599));
  MUX21X1 U993(.IN1(n600),.IN2(n599),.S(n143),.Q(n601));
  MUX21X1 U994(.IN1(n130),.IN2(n601),.S(n144),.Q(n602));
  MUX21X1 U995(.IN1(n609),.IN2(n602),.S(n64),.Q(n603));
  AND2X1 U996(.IN1(n603),.IN2(n59),.Q(dvsor_27_o[23:23]));
  NOR3X0 U997(.IN1(s_div_zeros[4:4]),.IN2(n17),.IN3(n604),.QN(dvsor_27_o[2:2]));
  NOR3X0 U998(.IN1(s_div_zeros[4:4]),.IN2(n18),.IN3(n605),.QN(dvsor_27_o[3:3]));
  NOR3X0 U999(.IN1(s_div_zeros[4:4]),.IN2(s_div_zeros[5:5]),.IN3(n606),.QN(dvsor_27_o[4:4]));
  NOR3X0 U1000(.IN1(n607),.IN2(n17),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[5:5]));
  NOR3X0 U1001(.IN1(n608),.IN2(n18),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[6:6]));
  AND3X1 U1002(.IN1(n609),.IN2(n59),.IN3(n64),.Q(dvsor_27_o[7:7]));
  MUX21X1 U1003(.IN1(n611),.IN2(n119),.S(n144),.Q(n612));
  AND3X1 U1004(.IN1(n64),.IN2(n59),.IN3(n612),.Q(dvsor_27_o[8:8]));
  MUX21X1 U1005(.IN1(n126),.IN2(n614),.S(n144),.Q(n615));
  NOR3X0 U1006(.IN1(n615),.IN2(s_div_zeros[5:5]),.IN3(s_div_zeros[4:4]),.QN(dvsor_27_o[9:9]));
assign dvsor_27_o[24:24]=1'b0;
assign dvsor_27_o[25:25]=1'b0;
assign dvsor_27_o[26:26]=1'b0;
assign dvdnd_50_o[0:0]=1'b0;
assign dvdnd_50_o[1:1]=1'b0;
assign dvdnd_50_o[2:2]=1'b0;
assign dvdnd_50_o[3:3]=1'b0;
assign dvdnd_50_o[4:4]=1'b0;
assign dvdnd_50_o[5:5]=1'b0;
assign dvdnd_50_o[6:6]=1'b0;
assign dvdnd_50_o[7:7]=1'b0;
assign dvdnd_50_o[8:8]=1'b0;
assign dvdnd_50_o[9:9]=1'b0;
assign dvdnd_50_o[10:10]=1'b0;
assign dvdnd_50_o[11:11]=1'b0;
assign dvdnd_50_o[12:12]=1'b0;
assign dvdnd_50_o[13:13]=1'b0;
assign dvdnd_50_o[14:14]=1'b0;
assign dvdnd_50_o[15:15]=1'b0;
assign dvdnd_50_o[16:16]=1'b0;
assign dvdnd_50_o[17:17]=1'b0;
assign dvdnd_50_o[18:18]=1'b0;
assign dvdnd_50_o[19:19]=1'b0;
assign dvdnd_50_o[20:20]=1'b0;
assign dvdnd_50_o[21:21]=1'b0;
assign dvdnd_50_o[22:22]=1'b0;
assign dvdnd_50_o[23:23]=1'b0;
assign dvdnd_50_o[24:24]=1'b0;
assign dvdnd_50_o[25:25]=1'b0;
endmodule
module serial_div_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [26:0] A ;
input [26:0] B ;
output [26:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire [27:0] carry ;
// instances
  FADDX1 U2_25(.A(A[25:25]),.B(n3),.CI(carry[25:25]),.CO(carry[26:26]),.S(DIFF[25:25]));
  FADDX1 U2_24(.A(A[24:24]),.B(n4),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n5),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n6),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n7),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n8),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n9),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n10),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n11),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n12),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n13),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n14),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n15),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n16),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n17),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n18),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n19),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n20),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n21),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n22),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n23),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n24),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n25),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n26),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n27),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_26(.IN1(A[26:26]),.IN2(n2),.IN3(carry[26:26]),.Q(DIFF[26:26]));
  INVX0 U1(.INP(B[6:6]),.ZN(n22));
  INVX0 U2(.INP(B[10:10]),.ZN(n18));
  INVX0 U3(.INP(B[14:14]),.ZN(n14));
  INVX0 U4(.INP(B[18:18]),.ZN(n10));
  INVX0 U5(.INP(B[16:16]),.ZN(n12));
  INVX0 U6(.INP(B[20:20]),.ZN(n8));
  INVX0 U7(.INP(B[22:22]),.ZN(n6));
  INVX0 U8(.INP(B[2:2]),.ZN(n26));
  INVX0 U9(.INP(B[1:1]),.ZN(n27));
  NAND2X1 U10(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U11(.INP(A[0:0]),.ZN(n1));
  INVX0 U12(.INP(B[3:3]),.ZN(n25));
  INVX0 U13(.INP(B[4:4]),.ZN(n24));
  INVX0 U14(.INP(B[7:7]),.ZN(n21));
  INVX0 U15(.INP(B[8:8]),.ZN(n20));
  INVX0 U16(.INP(B[11:11]),.ZN(n17));
  INVX0 U17(.INP(B[12:12]),.ZN(n16));
  INVX0 U18(.INP(B[15:15]),.ZN(n13));
  INVX0 U19(.INP(B[17:17]),.ZN(n11));
  INVX0 U20(.INP(B[19:19]),.ZN(n9));
  INVX0 U21(.INP(B[21:21]),.ZN(n7));
  INVX0 U22(.INP(B[23:23]),.ZN(n5));
  INVX0 U23(.INP(B[5:5]),.ZN(n23));
  INVX0 U24(.INP(B[9:9]),.ZN(n19));
  INVX0 U25(.INP(B[13:13]),.ZN(n15));
  INVX0 U26(.INP(B[24:24]),.ZN(n4));
  INVX0 U27(.INP(B[25:25]),.ZN(n3));
  INVX0 U28(.INP(B[26:26]),.ZN(n2));
  XOR2X1 U29(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module serial_div_DW_cmp_0_inj (A,B,TC,GE_LT,GE_GT_EQ,GE_LT_GT_LE,EQ_NE);
input [26:0] A ;
input [26:0] B ;
input TC ;
input GE_LT ;
input GE_GT_EQ ;
output GE_LT_GT_LE ;
output EQ_NE ;
wire n1069 ;
wire n1070 ;
wire n1071 ;
wire n1072 ;
wire n1073 ;
wire n1074 ;
wire n1075 ;
wire n1076 ;
wire n1077 ;
wire n1078 ;
wire n1079 ;
wire n1080 ;
wire n1081 ;
wire n1082 ;
wire n1083 ;
wire n1084 ;
wire n1085 ;
wire n1086 ;
wire n1087 ;
wire n1088 ;
wire n1089 ;
wire n1090 ;
wire n1091 ;
wire n1092 ;
wire n1093 ;
wire n1094 ;
wire n1095 ;
wire n1096 ;
wire n1097 ;
wire n1098 ;
wire n1099 ;
wire n1100 ;
wire n1101 ;
wire n1102 ;
wire n1103 ;
wire n1104 ;
wire n1105 ;
wire n1106 ;
wire n1107 ;
wire n1108 ;
wire n1109 ;
wire n1110 ;
wire n1111 ;
wire n1112 ;
wire n1113 ;
wire n1114 ;
wire n1115 ;
wire n1116 ;
wire n1117 ;
wire n1118 ;
wire n1119 ;
wire n1120 ;
wire n1121 ;
wire n1122 ;
wire n1123 ;
wire n1124 ;
wire n1125 ;
wire n1126 ;
wire n1127 ;
wire n1128 ;
wire n1129 ;
wire n1130 ;
wire n1131 ;
wire n1132 ;
wire n1133 ;
wire n1134 ;
wire n1135 ;
wire n1136 ;
wire n1137 ;
wire n1138 ;
wire n1139 ;
wire n1140 ;
wire n1141 ;
wire n1142 ;
wire n1143 ;
wire n1144 ;
wire n1145 ;
wire n1146 ;
wire n1147 ;
wire n1148 ;
wire n1149 ;
wire n1150 ;
wire n1151 ;
wire n1152 ;
wire n1153 ;
wire n1154 ;
wire n1155 ;
wire n1156 ;
wire n1157 ;
wire n1158 ;
wire n1159 ;
wire n1160 ;
wire n1161 ;
wire n1162 ;
wire n1163 ;
wire n1164 ;
wire n1165 ;
wire n1166 ;
wire n1167 ;
wire n1168 ;
wire n1169 ;
wire n1170 ;
wire n1171 ;
wire n1172 ;
wire n1173 ;
// instances
  INVX0 U545(.INP(n1114),.ZN(n1075));
  INVX0 U546(.INP(A[12:12]),.ZN(n1080));
  INVX0 U547(.INP(A[8:8]),.ZN(n1083));
  INVX0 U548(.INP(A[4:4]),.ZN(n1086));
  INVX0 U549(.INP(A[21:21]),.ZN(n1072));
  INVX0 U550(.INP(A[17:17]),.ZN(n1076));
  INVX0 U551(.INP(A[3:3]),.ZN(n1087));
  INVX0 U552(.INP(A[23:23]),.ZN(n1070));
  INVX0 U553(.INP(A[19:19]),.ZN(n1074));
  INVX0 U554(.INP(A[11:11]),.ZN(n1082));
  INVX0 U555(.INP(A[7:7]),.ZN(n1085));
  INVX0 U556(.INP(A[15:15]),.ZN(n1079));
  INVX0 U557(.INP(A[25:25]),.ZN(n1102));
  INVX0 U558(.INP(A[26:26]),.ZN(n1103));
  INVX0 U559(.INP(n1109),.ZN(n1069));
  INVX0 U560(.INP(n1140),.ZN(n1084));
  INVX0 U561(.INP(n1156),.ZN(n1089));
  INVX0 U562(.INP(A[24:24]),.ZN(n1101));
  INVX0 U563(.INP(n1164),.ZN(n1071));
  INVX0 U564(.INP(B[20:20]),.ZN(n1091));
  INVX0 U565(.INP(n1129),.ZN(n1078));
  INVX0 U566(.INP(n1120),.ZN(n1081));
  INVX0 U567(.INP(n1119),.ZN(n1077));
  INVX0 U568(.INP(B[18:18]),.ZN(n1092));
  INVX0 U569(.INP(A[1:1]),.ZN(n1088));
  INVX0 U570(.INP(B[14:14]),.ZN(n1094));
  INVX0 U571(.INP(B[6:6]),.ZN(n1098));
  INVX0 U572(.INP(B[10:10]),.ZN(n1096));
  INVX0 U573(.INP(n1108),.ZN(n1073));
  INVX0 U574(.INP(B[2:2]),.ZN(n1100));
  INVX0 U575(.INP(B[22:22]),.ZN(n1090));
  INVX0 U576(.INP(B[13:13]),.ZN(n1095));
  INVX0 U577(.INP(B[9:9]),.ZN(n1097));
  INVX0 U578(.INP(B[5:5]),.ZN(n1099));
  INVX0 U579(.INP(B[16:16]),.ZN(n1093));
  AO21X1 U580(.IN1(n1104),.IN2(n1105),.IN3(n1106),.Q(GE_LT_GT_LE));
  NOR4X0 U581(.IN1(n1107),.IN2(n1108),.IN3(n1109),.IN4(n1110),.QN(n1106));
  NAND4X0 U582(.IN1(n1111),.IN2(n1112),.IN3(n1075),.IN4(n1113),.QN(n1107));
  NAND2X0 U583(.IN1(A[16:16]),.IN2(n1093),.QN(n1113));
  NAND2X0 U584(.IN1(n1115),.IN2(n1116),.QN(n1112));
  NAND4X0 U585(.IN1(n1081),.IN2(n1077),.IN3(n1117),.IN4(n1118),.QN(n1116));
  OR2X1 U586(.IN1(n1083),.IN2(B[8:8]),.Q(n1118));
  NAND3X0 U587(.IN1(n1121),.IN2(n1122),.IN3(n1115),.QN(n1111));
  AND2X1 U588(.IN1(n1123),.IN2(n1124),.Q(n1115));
  AO221X1 U589(.IN1(n1125),.IN2(n1120),.IN3(n1126),.IN4(n1125),.IN5(n1119),.Q(n1124));
  NAND3X0 U590(.IN1(n1127),.IN2(n1128),.IN3(n1078),.QN(n1119));
  OR2X1 U591(.IN1(n1080),.IN2(B[12:12]),.Q(n1128));
  OA21X1 U592(.IN1(A[9:9]),.IN2(n1097),.IN3(n1130),.Q(n1126));
  NAND3X0 U593(.IN1(n1117),.IN2(n1083),.IN3(B[8:8]),.QN(n1130));
  NAND2X0 U594(.IN1(A[9:9]),.IN2(n1097),.QN(n1117));
  AO21X1 U595(.IN1(A[10:10]),.IN2(n1096),.IN3(n1131),.Q(n1120));
  AOI22X1 U596(.IN1(B[11:11]),.IN2(n1082),.IN3(n1132),.IN4(B[10:10]),.QN(n1125));
  NOR2X0 U597(.IN1(A[10:10]),.IN2(n1131),.QN(n1132));
  NOR2X0 U598(.IN1(n1082),.IN2(B[11:11]),.QN(n1131));
  AO22X1 U599(.IN1(n1133),.IN2(n1134),.IN3(n1134),.IN4(n1129),.Q(n1123));
  AO21X1 U600(.IN1(A[14:14]),.IN2(n1094),.IN3(n1135),.Q(n1129));
  AOI22X1 U601(.IN1(B[15:15]),.IN2(n1079),.IN3(n1136),.IN4(B[14:14]),.QN(n1134));
  NOR2X0 U602(.IN1(A[14:14]),.IN2(n1135),.QN(n1136));
  NOR2X0 U603(.IN1(n1079),.IN2(B[15:15]),.QN(n1135));
  OA21X1 U604(.IN1(A[13:13]),.IN2(n1095),.IN3(n1137),.Q(n1133));
  NAND3X0 U605(.IN1(n1127),.IN2(n1080),.IN3(B[12:12]),.QN(n1137));
  NAND2X0 U606(.IN1(A[13:13]),.IN2(n1095),.QN(n1127));
  AO22X1 U607(.IN1(n1138),.IN2(n1139),.IN3(n1139),.IN4(n1140),.Q(n1122));
  AOI22X1 U608(.IN1(B[7:7]),.IN2(n1085),.IN3(n1141),.IN4(B[6:6]),.QN(n1139));
  NOR2X0 U609(.IN1(A[6:6]),.IN2(n1142),.QN(n1141));
  OA21X1 U610(.IN1(A[5:5]),.IN2(n1099),.IN3(n1143),.Q(n1138));
  NAND3X0 U611(.IN1(n1144),.IN2(n1086),.IN3(B[4:4]),.QN(n1143));
  NAND3X0 U612(.IN1(n1084),.IN2(n1145),.IN3(n1146),.QN(n1121));
  OA221X1 U613(.IN1(n1147),.IN2(n1148),.IN3(B[4:4]),.IN4(n1086),.IN5(n1144),.Q(n1146));
  NAND2X0 U614(.IN1(A[5:5]),.IN2(n1099),.QN(n1144));
  AOI21X1 U615(.IN1(n1100),.IN2(A[2:2]),.IN3(n1149),.QN(n1147));
  AO221X1 U616(.IN1(B[1:1]),.IN2(n1088),.IN3(n1150),.IN4(B[0:0]),.IN5(n1148),.Q(n1145));
  AO22X1 U617(.IN1(B[3:3]),.IN2(n1087),.IN3(n1151),.IN4(B[2:2]),.Q(n1148));
  NOR2X0 U618(.IN1(A[2:2]),.IN2(n1149),.QN(n1151));
  NOR2X0 U619(.IN1(n1087),.IN2(B[3:3]),.QN(n1149));
  NOR2X0 U620(.IN1(A[0:0]),.IN2(n1152),.QN(n1150));
  NOR2X0 U621(.IN1(B[1:1]),.IN2(n1088),.QN(n1152));
  AO21X1 U622(.IN1(A[6:6]),.IN2(n1098),.IN3(n1142),.Q(n1140));
  NOR2X0 U623(.IN1(n1085),.IN2(B[7:7]),.QN(n1142));
  NAND2X0 U624(.IN1(n1089),.IN2(n1110),.QN(n1105));
  OR3X1 U625(.IN1(n1153),.IN2(n1154),.IN3(n1155),.Q(n1110));
  NOR2X0 U626(.IN1(n1101),.IN2(B[24:24]),.QN(n1154));
  AO221X1 U627(.IN1(n1157),.IN2(n1158),.IN3(n1159),.IN4(n1069),.IN5(n1156),.Q(n1104));
  AO22X1 U628(.IN1(B[26:26]),.IN2(n1103),.IN3(n1160),.IN4(n1161),.Q(n1156));
  AO22X1 U629(.IN1(B[25:25]),.IN2(n1102),.IN3(B[24:24]),.IN4(n1101),.Q(n1161));
  NOR2X0 U630(.IN1(n1153),.IN2(n1155),.QN(n1160));
  NOR2X0 U631(.IN1(n1103),.IN2(B[26:26]),.QN(n1155));
  NOR2X0 U632(.IN1(n1102),.IN2(B[25:25]),.QN(n1153));
  NAND3X0 U633(.IN1(n1071),.IN2(n1162),.IN3(n1163),.QN(n1109));
  NAND2X0 U634(.IN1(A[20:20]),.IN2(n1091),.QN(n1162));
  OA21X1 U635(.IN1(n1073),.IN2(n1165),.IN3(n1166),.Q(n1159));
  AO221X1 U636(.IN1(B[17:17]),.IN2(n1076),.IN3(n1167),.IN4(B[16:16]),.IN5(n1165),.Q(n1166));
  NOR2X0 U637(.IN1(A[16:16]),.IN2(n1114),.QN(n1167));
  NOR2X0 U638(.IN1(n1076),.IN2(B[17:17]),.QN(n1114));
  AO22X1 U639(.IN1(B[19:19]),.IN2(n1074),.IN3(n1168),.IN4(B[18:18]),.Q(n1165));
  NOR2X0 U640(.IN1(A[18:18]),.IN2(n1169),.QN(n1168));
  AO21X1 U641(.IN1(A[18:18]),.IN2(n1092),.IN3(n1169),.Q(n1108));
  NOR2X0 U642(.IN1(n1074),.IN2(B[19:19]),.QN(n1169));
  OR2X1 U643(.IN1(n1170),.IN2(n1163),.Q(n1158));
  AOI21X1 U644(.IN1(A[22:22]),.IN2(n1090),.IN3(n1171),.QN(n1163));
  AO221X1 U645(.IN1(B[21:21]),.IN2(n1072),.IN3(n1172),.IN4(B[20:20]),.IN5(n1170),.Q(n1157));
  AO22X1 U646(.IN1(B[23:23]),.IN2(n1070),.IN3(n1173),.IN4(B[22:22]),.Q(n1170));
  NOR2X0 U647(.IN1(A[22:22]),.IN2(n1171),.QN(n1173));
  NOR2X0 U648(.IN1(n1070),.IN2(B[23:23]),.QN(n1171));
  NOR2X0 U649(.IN1(A[20:20]),.IN2(n1164),.QN(n1172));
  NOR2X0 U650(.IN1(n1072),.IN2(B[21:21]),.QN(n1164));
endmodule
module serial_div_inj (clk_i,dvdnd_i,dvsor_i,sign_dvd_i,sign_div_i,start_i,ready_o,qutnt_o,rmndr_o,sign_o,div_zero_o,p_desc1368_p_O_DFFX1,p_desc1369_p_O_DFFX1,p_desc1370_p_O_DFFX1,p_desc1371_p_O_DFFX1,p_desc1372_p_O_DFFX1,p_desc1373_p_O_DFFX1,p_desc1374_p_O_DFFX1,p_desc1375_p_O_DFFX1,p_desc1376_p_O_DFFX1,p_desc1377_p_O_DFFX1,p_desc1378_p_O_DFFX1,p_desc1379_p_O_DFFX1,p_desc1380_p_O_DFFX1,p_desc1381_p_O_DFFX1,p_desc1382_p_O_DFFX1,p_desc1383_p_O_DFFX1,p_desc1384_p_O_DFFX1,p_desc1385_p_O_DFFX1,p_desc1386_p_O_DFFX1,p_desc1387_p_O_DFFX1,p_desc1388_p_O_DFFX1,p_desc1389_p_O_DFFX1,p_desc1390_p_O_DFFX1,p_desc1391_p_O_DFFX1,p_desc1392_p_O_DFFX1,p_desc1393_p_O_DFFX1,p_desc1394_p_O_DFFX1,p_desc1395_p_O_DFFX1,p_desc1396_p_O_DFFX1,p_desc1397_p_O_DFFX1,p_desc1398_p_O_DFFX1,p_desc1399_p_O_DFFX1,p_desc1400_p_O_DFFX1,p_desc1401_p_O_DFFX1,p_desc1402_p_O_DFFX1,p_desc1403_p_O_DFFX1,p_desc1404_p_O_DFFX1,p_desc1405_p_O_DFFX1,p_desc1406_p_O_DFFX1,p_desc1407_p_O_DFFX1,p_desc1408_p_O_DFFX1,p_desc1409_p_O_DFFX1,p_desc1410_p_O_DFFX1,p_desc1411_p_O_DFFX1,p_desc1412_p_O_DFFX1,p_desc1413_p_O_DFFX1,p_desc1414_p_O_DFFX1,p_desc1415_p_O_DFFX1,p_desc1416_p_O_DFFX1,p_desc1417_p_O_DFFX1,p_desc1418_p_O_DFFX1,p_desc1419_p_O_DFFX1,p_desc1420_p_O_DFFX1,p_desc1421_p_O_DFFX1,p_desc1422_p_O_DFFX1,p_desc1423_p_O_DFFX1,p_desc1424_p_O_DFFX1,p_desc1425_p_O_DFFX1,p_desc1426_p_O_DFFX1,p_desc1427_p_O_DFFX1,p_desc1428_p_O_DFFX1,p_desc1429_p_O_DFFX1,p_desc1430_p_O_DFFX1,p_desc1431_p_O_DFFX1,p_desc1432_p_O_DFFX1,p_desc1433_p_O_DFFX1,p_desc1434_p_O_DFFX1,p_desc1435_p_O_DFFX1,p_desc1436_p_O_DFFX1,p_desc1437_p_O_DFFX1,p_desc1438_p_O_DFFX1,p_desc1439_p_O_DFFX1,p_desc1440_p_O_DFFX1,p_desc1441_p_O_DFFX1,p_desc1442_p_O_DFFX1,p_desc1443_p_O_DFFX1,p_desc1444_p_O_DFFX1,p_s_start_i_reg_p_O_DFFX1,p_s_ready_o_reg_p_O_DFFX1,p_desc1445_p_O_DFFX1,p_desc1446_p_O_DFFX1,p_desc1447_p_O_DFFX1,p_desc1448_p_O_DFFX1,p_desc1449_p_O_DFFX1,p_desc1450_p_O_DFFX1,p_desc1451_p_O_DFFX1,p_desc1452_p_O_DFFX1,p_desc1453_p_O_DFFX1,p_desc1454_p_O_DFFX1,p_desc1455_p_O_DFFX1,p_desc1456_p_O_DFFX1,p_desc1457_p_O_DFFX1,p_desc1458_p_O_DFFX1,p_desc1459_p_O_DFFX1,p_desc1460_p_O_DFFX1,p_desc1461_p_O_DFFX1,p_desc1462_p_O_DFFX1,p_desc1463_p_O_DFFX1,p_desc1464_p_O_DFFX1,p_desc1465_p_O_DFFX1,p_desc1466_p_O_DFFX1,p_desc1467_p_O_DFFX1,p_desc1468_p_O_DFFX1,p_desc1469_p_O_DFFX1,p_desc1470_p_O_DFFX1,p_desc1471_p_O_DFFX1,p_desc1472_p_O_DFFX1,p_desc1473_p_O_DFFX1,p_desc1474_p_O_DFFX1,p_desc1475_p_O_DFFX1,p_desc1476_p_O_DFFX1,p_desc1477_p_O_DFFX1,p_desc1478_p_O_DFFX1,p_desc1479_p_O_DFFX1,p_desc1480_p_O_DFFX1,p_desc1481_p_O_DFFX1,p_desc1482_p_O_DFFX1,p_desc1483_p_O_DFFX1,p_desc1484_p_O_DFFX1,p_desc1485_p_O_DFFX1,p_desc1486_p_O_DFFX1,p_desc1487_p_O_DFFX1,p_desc1488_p_O_DFFX1,p_desc1489_p_O_DFFX1,p_desc1490_p_O_DFFX1,p_desc1491_p_O_DFFX1,p_desc1492_p_O_DFFX1,p_desc1493_p_O_DFFX1,p_desc1494_p_O_DFFX1,p_desc1495_p_O_DFFX1,p_desc1496_p_O_DFFX1,p_desc1497_p_O_DFFX1,p_desc1498_p_O_DFFX1,p_desc1499_p_O_DFFX1,p_desc1500_p_O_DFFX1,p_desc1501_p_O_DFFX1,p_desc1502_p_O_DFFX1,p_desc1503_p_O_DFFX1,p_desc1504_p_O_DFFX1,p_desc1505_p_O_DFFX1,p_desc1506_p_O_DFFX1,p_desc1507_p_O_DFFX1,p_desc1508_p_O_DFFX1,p_desc1509_p_O_DFFX1,p_desc1510_p_O_DFFX1,p_desc1511_p_O_DFFX1,p_desc1512_p_O_DFFX1,p_desc1513_p_O_DFFX1,p_desc1514_p_O_DFFX1,p_desc1515_p_O_DFFX1,p_desc1516_p_O_DFFX1,p_desc1517_p_O_DFFX1,p_desc1518_p_O_DFFX1,p_desc1519_p_O_DFFX1,p_desc1520_p_O_DFFX1,p_desc1521_p_O_DFFX1,p_desc1522_p_O_DFFX1,p_desc1523_p_O_DFFX1,p_desc1524_p_O_DFFX1,p_desc1525_p_O_DFFX1,p_desc1526_p_O_DFFX1,p_desc1527_p_O_DFFX1,p_desc1528_p_O_DFFX1,p_s_state_reg_p_O_DFFX1,p_desc1529_p_O_DFFX1);
input [49:0] dvdnd_i ;
input [26:0] dvsor_i ;
output [26:0] qutnt_o ;
output [26:0] rmndr_o ;
input clk_i ;
input sign_dvd_i ;
input sign_div_i ;
input start_i ;
output ready_o ;
output sign_o ;
output div_zero_o ;
wire s_start_i ;
wire N102 ;
wire s_state ;
wire N110 ;
wire N111 ;
wire N112 ;
wire N113 ;
wire N132 ;
wire N133 ;
wire N134 ;
wire N135 ;
wire N136 ;
wire N137 ;
wire N138 ;
wire N139 ;
wire N140 ;
wire N141 ;
wire N142 ;
wire N143 ;
wire N144 ;
wire N145 ;
wire N146 ;
wire N147 ;
wire N148 ;
wire N149 ;
wire N150 ;
wire N151 ;
wire N152 ;
wire N153 ;
wire N154 ;
wire N155 ;
wire N156 ;
wire N157 ;
wire N158 ;
wire N160 ;
wire N161 ;
wire N162 ;
wire N163 ;
wire N164 ;
wire N165 ;
wire N166 ;
wire N167 ;
wire N168 ;
wire N169 ;
wire N170 ;
wire N171 ;
wire N172 ;
wire N173 ;
wire N174 ;
wire N175 ;
wire N176 ;
wire N177 ;
wire N178 ;
wire N179 ;
wire N180 ;
wire N181 ;
wire N182 ;
wire N183 ;
wire N184 ;
wire N185 ;
wire N186 ;
wire n8 ;
wire n38 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n39 ;
wire n40 ;
wire n47 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire [49:0] s_dvdnd_i ;
wire [26:0] s_dvsor_i ;
wire [4:0] s_count ;
wire [26:0] s_dvd ;
input p_desc1368_p_O_DFFX1 ;
input p_desc1369_p_O_DFFX1 ;
input p_desc1370_p_O_DFFX1 ;
input p_desc1371_p_O_DFFX1 ;
input p_desc1372_p_O_DFFX1 ;
input p_desc1373_p_O_DFFX1 ;
input p_desc1374_p_O_DFFX1 ;
input p_desc1375_p_O_DFFX1 ;
input p_desc1376_p_O_DFFX1 ;
input p_desc1377_p_O_DFFX1 ;
input p_desc1378_p_O_DFFX1 ;
input p_desc1379_p_O_DFFX1 ;
input p_desc1380_p_O_DFFX1 ;
input p_desc1381_p_O_DFFX1 ;
input p_desc1382_p_O_DFFX1 ;
input p_desc1383_p_O_DFFX1 ;
input p_desc1384_p_O_DFFX1 ;
input p_desc1385_p_O_DFFX1 ;
input p_desc1386_p_O_DFFX1 ;
input p_desc1387_p_O_DFFX1 ;
input p_desc1388_p_O_DFFX1 ;
input p_desc1389_p_O_DFFX1 ;
input p_desc1390_p_O_DFFX1 ;
input p_desc1391_p_O_DFFX1 ;
input p_desc1392_p_O_DFFX1 ;
input p_desc1393_p_O_DFFX1 ;
input p_desc1394_p_O_DFFX1 ;
input p_desc1395_p_O_DFFX1 ;
input p_desc1396_p_O_DFFX1 ;
input p_desc1397_p_O_DFFX1 ;
input p_desc1398_p_O_DFFX1 ;
input p_desc1399_p_O_DFFX1 ;
input p_desc1400_p_O_DFFX1 ;
input p_desc1401_p_O_DFFX1 ;
input p_desc1402_p_O_DFFX1 ;
input p_desc1403_p_O_DFFX1 ;
input p_desc1404_p_O_DFFX1 ;
input p_desc1405_p_O_DFFX1 ;
input p_desc1406_p_O_DFFX1 ;
input p_desc1407_p_O_DFFX1 ;
input p_desc1408_p_O_DFFX1 ;
input p_desc1409_p_O_DFFX1 ;
input p_desc1410_p_O_DFFX1 ;
input p_desc1411_p_O_DFFX1 ;
input p_desc1412_p_O_DFFX1 ;
input p_desc1413_p_O_DFFX1 ;
input p_desc1414_p_O_DFFX1 ;
input p_desc1415_p_O_DFFX1 ;
input p_desc1416_p_O_DFFX1 ;
input p_desc1417_p_O_DFFX1 ;
input p_desc1418_p_O_DFFX1 ;
input p_desc1419_p_O_DFFX1 ;
input p_desc1420_p_O_DFFX1 ;
input p_desc1421_p_O_DFFX1 ;
input p_desc1422_p_O_DFFX1 ;
input p_desc1423_p_O_DFFX1 ;
input p_desc1424_p_O_DFFX1 ;
input p_desc1425_p_O_DFFX1 ;
input p_desc1426_p_O_DFFX1 ;
input p_desc1427_p_O_DFFX1 ;
input p_desc1428_p_O_DFFX1 ;
input p_desc1429_p_O_DFFX1 ;
input p_desc1430_p_O_DFFX1 ;
input p_desc1431_p_O_DFFX1 ;
input p_desc1432_p_O_DFFX1 ;
input p_desc1433_p_O_DFFX1 ;
input p_desc1434_p_O_DFFX1 ;
input p_desc1435_p_O_DFFX1 ;
input p_desc1436_p_O_DFFX1 ;
input p_desc1437_p_O_DFFX1 ;
input p_desc1438_p_O_DFFX1 ;
input p_desc1439_p_O_DFFX1 ;
input p_desc1440_p_O_DFFX1 ;
input p_desc1441_p_O_DFFX1 ;
input p_desc1442_p_O_DFFX1 ;
input p_desc1443_p_O_DFFX1 ;
input p_desc1444_p_O_DFFX1 ;
input p_s_start_i_reg_p_O_DFFX1 ;
input p_s_ready_o_reg_p_O_DFFX1 ;
input p_desc1445_p_O_DFFX1 ;
input p_desc1446_p_O_DFFX1 ;
input p_desc1447_p_O_DFFX1 ;
input p_desc1448_p_O_DFFX1 ;
input p_desc1449_p_O_DFFX1 ;
input p_desc1450_p_O_DFFX1 ;
input p_desc1451_p_O_DFFX1 ;
input p_desc1452_p_O_DFFX1 ;
input p_desc1453_p_O_DFFX1 ;
input p_desc1454_p_O_DFFX1 ;
input p_desc1455_p_O_DFFX1 ;
input p_desc1456_p_O_DFFX1 ;
input p_desc1457_p_O_DFFX1 ;
input p_desc1458_p_O_DFFX1 ;
input p_desc1459_p_O_DFFX1 ;
input p_desc1460_p_O_DFFX1 ;
input p_desc1461_p_O_DFFX1 ;
input p_desc1462_p_O_DFFX1 ;
input p_desc1463_p_O_DFFX1 ;
input p_desc1464_p_O_DFFX1 ;
input p_desc1465_p_O_DFFX1 ;
input p_desc1466_p_O_DFFX1 ;
input p_desc1467_p_O_DFFX1 ;
input p_desc1468_p_O_DFFX1 ;
input p_desc1469_p_O_DFFX1 ;
input p_desc1470_p_O_DFFX1 ;
input p_desc1471_p_O_DFFX1 ;
input p_desc1472_p_O_DFFX1 ;
input p_desc1473_p_O_DFFX1 ;
input p_desc1474_p_O_DFFX1 ;
input p_desc1475_p_O_DFFX1 ;
input p_desc1476_p_O_DFFX1 ;
input p_desc1477_p_O_DFFX1 ;
input p_desc1478_p_O_DFFX1 ;
input p_desc1479_p_O_DFFX1 ;
input p_desc1480_p_O_DFFX1 ;
input p_desc1481_p_O_DFFX1 ;
input p_desc1482_p_O_DFFX1 ;
input p_desc1483_p_O_DFFX1 ;
input p_desc1484_p_O_DFFX1 ;
input p_desc1485_p_O_DFFX1 ;
input p_desc1486_p_O_DFFX1 ;
input p_desc1487_p_O_DFFX1 ;
input p_desc1488_p_O_DFFX1 ;
input p_desc1489_p_O_DFFX1 ;
input p_desc1490_p_O_DFFX1 ;
input p_desc1491_p_O_DFFX1 ;
input p_desc1492_p_O_DFFX1 ;
input p_desc1493_p_O_DFFX1 ;
input p_desc1494_p_O_DFFX1 ;
input p_desc1495_p_O_DFFX1 ;
input p_desc1496_p_O_DFFX1 ;
input p_desc1497_p_O_DFFX1 ;
input p_desc1498_p_O_DFFX1 ;
input p_desc1499_p_O_DFFX1 ;
input p_desc1500_p_O_DFFX1 ;
input p_desc1501_p_O_DFFX1 ;
input p_desc1502_p_O_DFFX1 ;
input p_desc1503_p_O_DFFX1 ;
input p_desc1504_p_O_DFFX1 ;
input p_desc1505_p_O_DFFX1 ;
input p_desc1506_p_O_DFFX1 ;
input p_desc1507_p_O_DFFX1 ;
input p_desc1508_p_O_DFFX1 ;
input p_desc1509_p_O_DFFX1 ;
input p_desc1510_p_O_DFFX1 ;
input p_desc1511_p_O_DFFX1 ;
input p_desc1512_p_O_DFFX1 ;
input p_desc1513_p_O_DFFX1 ;
input p_desc1514_p_O_DFFX1 ;
input p_desc1515_p_O_DFFX1 ;
input p_desc1516_p_O_DFFX1 ;
input p_desc1517_p_O_DFFX1 ;
input p_desc1518_p_O_DFFX1 ;
input p_desc1519_p_O_DFFX1 ;
input p_desc1520_p_O_DFFX1 ;
input p_desc1521_p_O_DFFX1 ;
input p_desc1522_p_O_DFFX1 ;
input p_desc1523_p_O_DFFX1 ;
input p_desc1524_p_O_DFFX1 ;
input p_desc1525_p_O_DFFX1 ;
input p_desc1526_p_O_DFFX1 ;
input p_desc1527_p_O_DFFX1 ;
input p_desc1528_p_O_DFFX1 ;
input p_s_state_reg_p_O_DFFX1 ;
input p_desc1529_p_O_DFFX1 ;
// instances
  p_O_DFFX1 desc1368(.D(dvdnd_i[49:49]),.CLK(clk_i),.Q(s_dvdnd_i[49:49]),.QN(n8),.E(p_desc1368_p_O_DFFX1));
  p_O_DFFX1 desc1369(.D(dvdnd_i[48:48]),.CLK(clk_i),.Q(s_dvdnd_i[48:48]),.E(p_desc1369_p_O_DFFX1));
  p_O_DFFX1 desc1370(.D(dvdnd_i[47:47]),.CLK(clk_i),.Q(s_dvdnd_i[47:47]),.E(p_desc1370_p_O_DFFX1));
  p_O_DFFX1 desc1371(.D(dvdnd_i[46:46]),.CLK(clk_i),.Q(s_dvdnd_i[46:46]),.E(p_desc1371_p_O_DFFX1));
  p_O_DFFX1 desc1372(.D(dvdnd_i[45:45]),.CLK(clk_i),.Q(s_dvdnd_i[45:45]),.E(p_desc1372_p_O_DFFX1));
  p_O_DFFX1 desc1373(.D(dvdnd_i[44:44]),.CLK(clk_i),.Q(s_dvdnd_i[44:44]),.E(p_desc1373_p_O_DFFX1));
  p_O_DFFX1 desc1374(.D(dvdnd_i[43:43]),.CLK(clk_i),.Q(s_dvdnd_i[43:43]),.E(p_desc1374_p_O_DFFX1));
  p_O_DFFX1 desc1375(.D(dvdnd_i[42:42]),.CLK(clk_i),.Q(s_dvdnd_i[42:42]),.E(p_desc1375_p_O_DFFX1));
  p_O_DFFX1 desc1376(.D(dvdnd_i[41:41]),.CLK(clk_i),.Q(s_dvdnd_i[41:41]),.E(p_desc1376_p_O_DFFX1));
  p_O_DFFX1 desc1377(.D(dvdnd_i[40:40]),.CLK(clk_i),.Q(s_dvdnd_i[40:40]),.E(p_desc1377_p_O_DFFX1));
  p_O_DFFX1 desc1378(.D(dvdnd_i[39:39]),.CLK(clk_i),.Q(s_dvdnd_i[39:39]),.E(p_desc1378_p_O_DFFX1));
  p_O_DFFX1 desc1379(.D(dvdnd_i[38:38]),.CLK(clk_i),.Q(s_dvdnd_i[38:38]),.E(p_desc1379_p_O_DFFX1));
  p_O_DFFX1 desc1380(.D(dvdnd_i[37:37]),.CLK(clk_i),.Q(s_dvdnd_i[37:37]),.E(p_desc1380_p_O_DFFX1));
  p_O_DFFX1 desc1381(.D(dvdnd_i[36:36]),.CLK(clk_i),.Q(s_dvdnd_i[36:36]),.E(p_desc1381_p_O_DFFX1));
  p_O_DFFX1 desc1382(.D(dvdnd_i[35:35]),.CLK(clk_i),.Q(s_dvdnd_i[35:35]),.E(p_desc1382_p_O_DFFX1));
  p_O_DFFX1 desc1383(.D(dvdnd_i[34:34]),.CLK(clk_i),.Q(s_dvdnd_i[34:34]),.E(p_desc1383_p_O_DFFX1));
  p_O_DFFX1 desc1384(.D(dvdnd_i[33:33]),.CLK(clk_i),.Q(s_dvdnd_i[33:33]),.E(p_desc1384_p_O_DFFX1));
  p_O_DFFX1 desc1385(.D(dvdnd_i[32:32]),.CLK(clk_i),.Q(s_dvdnd_i[32:32]),.E(p_desc1385_p_O_DFFX1));
  p_O_DFFX1 desc1386(.D(dvdnd_i[31:31]),.CLK(clk_i),.Q(s_dvdnd_i[31:31]),.E(p_desc1386_p_O_DFFX1));
  p_O_DFFX1 desc1387(.D(dvdnd_i[30:30]),.CLK(clk_i),.Q(s_dvdnd_i[30:30]),.E(p_desc1387_p_O_DFFX1));
  p_O_DFFX1 desc1388(.D(dvdnd_i[29:29]),.CLK(clk_i),.Q(s_dvdnd_i[29:29]),.E(p_desc1388_p_O_DFFX1));
  p_O_DFFX1 desc1389(.D(dvdnd_i[28:28]),.CLK(clk_i),.Q(s_dvdnd_i[28:28]),.E(p_desc1389_p_O_DFFX1));
  p_O_DFFX1 desc1390(.D(dvdnd_i[27:27]),.CLK(clk_i),.Q(s_dvdnd_i[27:27]),.E(p_desc1390_p_O_DFFX1));
  p_O_DFFX1 desc1391(.D(dvdnd_i[26:26]),.CLK(clk_i),.Q(s_dvdnd_i[26:26]),.E(p_desc1391_p_O_DFFX1));
  p_O_DFFX1 desc1392(.D(dvdnd_i[25:25]),.CLK(clk_i),.Q(s_dvdnd_i[25:25]),.E(p_desc1392_p_O_DFFX1));
  p_O_DFFX1 desc1393(.D(dvdnd_i[24:24]),.CLK(clk_i),.Q(s_dvdnd_i[24:24]),.E(p_desc1393_p_O_DFFX1));
  p_O_DFFX1 desc1394(.D(dvdnd_i[23:23]),.CLK(clk_i),.Q(s_dvdnd_i[23:23]),.E(p_desc1394_p_O_DFFX1));
  p_O_DFFX1 desc1395(.D(dvdnd_i[22:22]),.CLK(clk_i),.Q(s_dvdnd_i[22:22]),.E(p_desc1395_p_O_DFFX1));
  p_O_DFFX1 desc1396(.D(dvdnd_i[21:21]),.CLK(clk_i),.Q(s_dvdnd_i[21:21]),.E(p_desc1396_p_O_DFFX1));
  p_O_DFFX1 desc1397(.D(dvdnd_i[20:20]),.CLK(clk_i),.Q(s_dvdnd_i[20:20]),.E(p_desc1397_p_O_DFFX1));
  p_O_DFFX1 desc1398(.D(dvdnd_i[19:19]),.CLK(clk_i),.Q(s_dvdnd_i[19:19]),.E(p_desc1398_p_O_DFFX1));
  p_O_DFFX1 desc1399(.D(dvdnd_i[18:18]),.CLK(clk_i),.Q(s_dvdnd_i[18:18]),.E(p_desc1399_p_O_DFFX1));
  p_O_DFFX1 desc1400(.D(dvdnd_i[17:17]),.CLK(clk_i),.Q(s_dvdnd_i[17:17]),.E(p_desc1400_p_O_DFFX1));
  p_O_DFFX1 desc1401(.D(dvdnd_i[16:16]),.CLK(clk_i),.Q(s_dvdnd_i[16:16]),.E(p_desc1401_p_O_DFFX1));
  p_O_DFFX1 desc1402(.D(dvdnd_i[15:15]),.CLK(clk_i),.Q(s_dvdnd_i[15:15]),.E(p_desc1402_p_O_DFFX1));
  p_O_DFFX1 desc1403(.D(dvdnd_i[14:14]),.CLK(clk_i),.Q(s_dvdnd_i[14:14]),.E(p_desc1403_p_O_DFFX1));
  p_O_DFFX1 desc1404(.D(dvdnd_i[13:13]),.CLK(clk_i),.Q(s_dvdnd_i[13:13]),.E(p_desc1404_p_O_DFFX1));
  p_O_DFFX1 desc1405(.D(dvdnd_i[12:12]),.CLK(clk_i),.Q(s_dvdnd_i[12:12]),.E(p_desc1405_p_O_DFFX1));
  p_O_DFFX1 desc1406(.D(dvdnd_i[11:11]),.CLK(clk_i),.Q(s_dvdnd_i[11:11]),.E(p_desc1406_p_O_DFFX1));
  p_O_DFFX1 desc1407(.D(dvdnd_i[10:10]),.CLK(clk_i),.Q(s_dvdnd_i[10:10]),.E(p_desc1407_p_O_DFFX1));
  p_O_DFFX1 desc1408(.D(dvdnd_i[9:9]),.CLK(clk_i),.Q(s_dvdnd_i[9:9]),.E(p_desc1408_p_O_DFFX1));
  p_O_DFFX1 desc1409(.D(dvdnd_i[8:8]),.CLK(clk_i),.Q(s_dvdnd_i[8:8]),.E(p_desc1409_p_O_DFFX1));
  p_O_DFFX1 desc1410(.D(dvdnd_i[7:7]),.CLK(clk_i),.Q(s_dvdnd_i[7:7]),.E(p_desc1410_p_O_DFFX1));
  p_O_DFFX1 desc1411(.D(dvdnd_i[6:6]),.CLK(clk_i),.Q(s_dvdnd_i[6:6]),.E(p_desc1411_p_O_DFFX1));
  p_O_DFFX1 desc1412(.D(dvdnd_i[5:5]),.CLK(clk_i),.Q(s_dvdnd_i[5:5]),.E(p_desc1412_p_O_DFFX1));
  p_O_DFFX1 desc1413(.D(dvdnd_i[4:4]),.CLK(clk_i),.Q(s_dvdnd_i[4:4]),.E(p_desc1413_p_O_DFFX1));
  p_O_DFFX1 desc1414(.D(dvdnd_i[3:3]),.CLK(clk_i),.Q(s_dvdnd_i[3:3]),.E(p_desc1414_p_O_DFFX1));
  p_O_DFFX1 desc1415(.D(dvdnd_i[2:2]),.CLK(clk_i),.Q(s_dvdnd_i[2:2]),.E(p_desc1415_p_O_DFFX1));
  p_O_DFFX1 desc1416(.D(dvdnd_i[1:1]),.CLK(clk_i),.Q(s_dvdnd_i[1:1]),.E(p_desc1416_p_O_DFFX1));
  p_O_DFFX1 desc1417(.D(dvdnd_i[0:0]),.CLK(clk_i),.Q(s_dvdnd_i[0:0]),.E(p_desc1417_p_O_DFFX1));
  p_O_DFFX1 desc1418(.D(dvsor_i[26:26]),.CLK(clk_i),.Q(s_dvsor_i[26:26]),.E(p_desc1418_p_O_DFFX1));
  p_O_DFFX1 desc1419(.D(dvsor_i[25:25]),.CLK(clk_i),.Q(s_dvsor_i[25:25]),.E(p_desc1419_p_O_DFFX1));
  p_O_DFFX1 desc1420(.D(dvsor_i[24:24]),.CLK(clk_i),.Q(s_dvsor_i[24:24]),.E(p_desc1420_p_O_DFFX1));
  p_O_DFFX1 desc1421(.D(dvsor_i[23:23]),.CLK(clk_i),.Q(s_dvsor_i[23:23]),.E(p_desc1421_p_O_DFFX1));
  p_O_DFFX1 desc1422(.D(dvsor_i[22:22]),.CLK(clk_i),.Q(s_dvsor_i[22:22]),.E(p_desc1422_p_O_DFFX1));
  p_O_DFFX1 desc1423(.D(dvsor_i[21:21]),.CLK(clk_i),.Q(s_dvsor_i[21:21]),.E(p_desc1423_p_O_DFFX1));
  p_O_DFFX1 desc1424(.D(dvsor_i[20:20]),.CLK(clk_i),.Q(s_dvsor_i[20:20]),.E(p_desc1424_p_O_DFFX1));
  p_O_DFFX1 desc1425(.D(dvsor_i[19:19]),.CLK(clk_i),.Q(s_dvsor_i[19:19]),.E(p_desc1425_p_O_DFFX1));
  p_O_DFFX1 desc1426(.D(dvsor_i[18:18]),.CLK(clk_i),.Q(s_dvsor_i[18:18]),.E(p_desc1426_p_O_DFFX1));
  p_O_DFFX1 desc1427(.D(dvsor_i[17:17]),.CLK(clk_i),.Q(s_dvsor_i[17:17]),.E(p_desc1427_p_O_DFFX1));
  p_O_DFFX1 desc1428(.D(dvsor_i[16:16]),.CLK(clk_i),.Q(s_dvsor_i[16:16]),.E(p_desc1428_p_O_DFFX1));
  p_O_DFFX1 desc1429(.D(dvsor_i[15:15]),.CLK(clk_i),.Q(s_dvsor_i[15:15]),.E(p_desc1429_p_O_DFFX1));
  p_O_DFFX1 desc1430(.D(dvsor_i[14:14]),.CLK(clk_i),.Q(s_dvsor_i[14:14]),.E(p_desc1430_p_O_DFFX1));
  p_O_DFFX1 desc1431(.D(dvsor_i[13:13]),.CLK(clk_i),.Q(s_dvsor_i[13:13]),.E(p_desc1431_p_O_DFFX1));
  p_O_DFFX1 desc1432(.D(dvsor_i[12:12]),.CLK(clk_i),.Q(s_dvsor_i[12:12]),.E(p_desc1432_p_O_DFFX1));
  p_O_DFFX1 desc1433(.D(dvsor_i[11:11]),.CLK(clk_i),.Q(s_dvsor_i[11:11]),.E(p_desc1433_p_O_DFFX1));
  p_O_DFFX1 desc1434(.D(dvsor_i[10:10]),.CLK(clk_i),.Q(s_dvsor_i[10:10]),.E(p_desc1434_p_O_DFFX1));
  p_O_DFFX1 desc1435(.D(dvsor_i[9:9]),.CLK(clk_i),.Q(s_dvsor_i[9:9]),.E(p_desc1435_p_O_DFFX1));
  p_O_DFFX1 desc1436(.D(dvsor_i[8:8]),.CLK(clk_i),.Q(s_dvsor_i[8:8]),.E(p_desc1436_p_O_DFFX1));
  p_O_DFFX1 desc1437(.D(dvsor_i[7:7]),.CLK(clk_i),.Q(s_dvsor_i[7:7]),.E(p_desc1437_p_O_DFFX1));
  p_O_DFFX1 desc1438(.D(dvsor_i[6:6]),.CLK(clk_i),.Q(s_dvsor_i[6:6]),.E(p_desc1438_p_O_DFFX1));
  p_O_DFFX1 desc1439(.D(dvsor_i[5:5]),.CLK(clk_i),.Q(s_dvsor_i[5:5]),.E(p_desc1439_p_O_DFFX1));
  p_O_DFFX1 desc1440(.D(dvsor_i[4:4]),.CLK(clk_i),.Q(s_dvsor_i[4:4]),.E(p_desc1440_p_O_DFFX1));
  p_O_DFFX1 desc1441(.D(dvsor_i[3:3]),.CLK(clk_i),.Q(s_dvsor_i[3:3]),.E(p_desc1441_p_O_DFFX1));
  p_O_DFFX1 desc1442(.D(dvsor_i[2:2]),.CLK(clk_i),.Q(s_dvsor_i[2:2]),.E(p_desc1442_p_O_DFFX1));
  p_O_DFFX1 desc1443(.D(dvsor_i[1:1]),.CLK(clk_i),.Q(s_dvsor_i[1:1]),.E(p_desc1443_p_O_DFFX1));
  p_O_DFFX1 desc1444(.D(dvsor_i[0:0]),.CLK(clk_i),.Q(s_dvsor_i[0:0]),.E(p_desc1444_p_O_DFFX1));
  p_O_DFFX1 s_start_i_reg(.D(start_i),.CLK(clk_i),.Q(s_start_i),.QN(n38),.E(p_s_start_i_reg_p_O_DFFX1));
  p_O_DFFX1 s_ready_o_reg(.D(n234),.CLK(clk_i),.Q(ready_o),.E(p_s_ready_o_reg_p_O_DFFX1));
  p_O_DFFX1 desc1445(.D(n236),.CLK(clk_i),.Q(s_count[4:4]),.E(p_desc1445_p_O_DFFX1));
  p_O_DFFX1 desc1446(.D(n233),.CLK(clk_i),.Q(s_count[1:1]),.QN(n43),.E(p_desc1446_p_O_DFFX1));
  p_O_DFFX1 desc1447(.D(n232),.CLK(clk_i),.Q(s_count[2:2]),.QN(n42),.E(p_desc1447_p_O_DFFX1));
  p_O_DFFX1 desc1448(.D(n231),.CLK(clk_i),.Q(s_count[3:3]),.QN(n41),.E(p_desc1448_p_O_DFFX1));
  p_O_DFFX1 desc1449(.D(n177),.CLK(clk_i),.Q(rmndr_o[0:0]),.E(p_desc1449_p_O_DFFX1));
  p_O_DFFX1 desc1450(.D(n203),.CLK(clk_i),.Q(s_dvd[1:1]),.E(p_desc1450_p_O_DFFX1));
  p_O_DFFX1 desc1451(.D(n176),.CLK(clk_i),.Q(rmndr_o[1:1]),.E(p_desc1451_p_O_DFFX1));
  p_O_DFFX1 desc1452(.D(n202),.CLK(clk_i),.Q(s_dvd[2:2]),.E(p_desc1452_p_O_DFFX1));
  p_O_DFFX1 desc1453(.D(n175),.CLK(clk_i),.Q(rmndr_o[2:2]),.E(p_desc1453_p_O_DFFX1));
  p_O_DFFX1 desc1454(.D(n201),.CLK(clk_i),.Q(s_dvd[3:3]),.E(p_desc1454_p_O_DFFX1));
  p_O_DFFX1 desc1455(.D(n174),.CLK(clk_i),.Q(rmndr_o[3:3]),.E(p_desc1455_p_O_DFFX1));
  p_O_DFFX1 desc1456(.D(n200),.CLK(clk_i),.Q(s_dvd[4:4]),.E(p_desc1456_p_O_DFFX1));
  p_O_DFFX1 desc1457(.D(n173),.CLK(clk_i),.Q(rmndr_o[4:4]),.E(p_desc1457_p_O_DFFX1));
  p_O_DFFX1 desc1458(.D(n199),.CLK(clk_i),.Q(s_dvd[5:5]),.E(p_desc1458_p_O_DFFX1));
  p_O_DFFX1 desc1459(.D(n172),.CLK(clk_i),.Q(rmndr_o[5:5]),.E(p_desc1459_p_O_DFFX1));
  p_O_DFFX1 desc1460(.D(n198),.CLK(clk_i),.Q(s_dvd[6:6]),.E(p_desc1460_p_O_DFFX1));
  p_O_DFFX1 desc1461(.D(n171),.CLK(clk_i),.Q(rmndr_o[6:6]),.E(p_desc1461_p_O_DFFX1));
  p_O_DFFX1 desc1462(.D(n197),.CLK(clk_i),.Q(s_dvd[7:7]),.E(p_desc1462_p_O_DFFX1));
  p_O_DFFX1 desc1463(.D(n170),.CLK(clk_i),.Q(rmndr_o[7:7]),.E(p_desc1463_p_O_DFFX1));
  p_O_DFFX1 desc1464(.D(n196),.CLK(clk_i),.Q(s_dvd[8:8]),.E(p_desc1464_p_O_DFFX1));
  p_O_DFFX1 desc1465(.D(n169),.CLK(clk_i),.Q(rmndr_o[8:8]),.E(p_desc1465_p_O_DFFX1));
  p_O_DFFX1 desc1466(.D(n195),.CLK(clk_i),.Q(s_dvd[9:9]),.E(p_desc1466_p_O_DFFX1));
  p_O_DFFX1 desc1467(.D(n168),.CLK(clk_i),.Q(rmndr_o[9:9]),.E(p_desc1467_p_O_DFFX1));
  p_O_DFFX1 desc1468(.D(n194),.CLK(clk_i),.Q(s_dvd[10:10]),.E(p_desc1468_p_O_DFFX1));
  p_O_DFFX1 desc1469(.D(n167),.CLK(clk_i),.Q(rmndr_o[10:10]),.E(p_desc1469_p_O_DFFX1));
  p_O_DFFX1 desc1470(.D(n193),.CLK(clk_i),.Q(s_dvd[11:11]),.E(p_desc1470_p_O_DFFX1));
  p_O_DFFX1 desc1471(.D(n166),.CLK(clk_i),.Q(rmndr_o[11:11]),.E(p_desc1471_p_O_DFFX1));
  p_O_DFFX1 desc1472(.D(n192),.CLK(clk_i),.Q(s_dvd[12:12]),.E(p_desc1472_p_O_DFFX1));
  p_O_DFFX1 desc1473(.D(n165),.CLK(clk_i),.Q(rmndr_o[12:12]),.E(p_desc1473_p_O_DFFX1));
  p_O_DFFX1 desc1474(.D(n191),.CLK(clk_i),.Q(s_dvd[13:13]),.E(p_desc1474_p_O_DFFX1));
  p_O_DFFX1 desc1475(.D(n164),.CLK(clk_i),.Q(rmndr_o[13:13]),.E(p_desc1475_p_O_DFFX1));
  p_O_DFFX1 desc1476(.D(n190),.CLK(clk_i),.Q(s_dvd[14:14]),.E(p_desc1476_p_O_DFFX1));
  p_O_DFFX1 desc1477(.D(n163),.CLK(clk_i),.Q(rmndr_o[14:14]),.E(p_desc1477_p_O_DFFX1));
  p_O_DFFX1 desc1478(.D(n189),.CLK(clk_i),.Q(s_dvd[15:15]),.E(p_desc1478_p_O_DFFX1));
  p_O_DFFX1 desc1479(.D(n162),.CLK(clk_i),.Q(rmndr_o[15:15]),.E(p_desc1479_p_O_DFFX1));
  p_O_DFFX1 desc1480(.D(n188),.CLK(clk_i),.Q(s_dvd[16:16]),.E(p_desc1480_p_O_DFFX1));
  p_O_DFFX1 desc1481(.D(n161),.CLK(clk_i),.Q(rmndr_o[16:16]),.E(p_desc1481_p_O_DFFX1));
  p_O_DFFX1 desc1482(.D(n187),.CLK(clk_i),.Q(s_dvd[17:17]),.E(p_desc1482_p_O_DFFX1));
  p_O_DFFX1 desc1483(.D(n160),.CLK(clk_i),.Q(rmndr_o[17:17]),.E(p_desc1483_p_O_DFFX1));
  p_O_DFFX1 desc1484(.D(n186),.CLK(clk_i),.Q(s_dvd[18:18]),.E(p_desc1484_p_O_DFFX1));
  p_O_DFFX1 desc1485(.D(n159),.CLK(clk_i),.Q(rmndr_o[18:18]),.E(p_desc1485_p_O_DFFX1));
  p_O_DFFX1 desc1486(.D(n185),.CLK(clk_i),.Q(s_dvd[19:19]),.E(p_desc1486_p_O_DFFX1));
  p_O_DFFX1 desc1487(.D(n158),.CLK(clk_i),.Q(rmndr_o[19:19]),.E(p_desc1487_p_O_DFFX1));
  p_O_DFFX1 desc1488(.D(n184),.CLK(clk_i),.Q(s_dvd[20:20]),.E(p_desc1488_p_O_DFFX1));
  p_O_DFFX1 desc1489(.D(n157),.CLK(clk_i),.Q(rmndr_o[20:20]),.E(p_desc1489_p_O_DFFX1));
  p_O_DFFX1 desc1490(.D(n183),.CLK(clk_i),.Q(s_dvd[21:21]),.E(p_desc1490_p_O_DFFX1));
  p_O_DFFX1 desc1491(.D(n156),.CLK(clk_i),.Q(rmndr_o[21:21]),.E(p_desc1491_p_O_DFFX1));
  p_O_DFFX1 desc1492(.D(n182),.CLK(clk_i),.Q(s_dvd[22:22]),.E(p_desc1492_p_O_DFFX1));
  p_O_DFFX1 desc1493(.D(n155),.CLK(clk_i),.Q(rmndr_o[22:22]),.E(p_desc1493_p_O_DFFX1));
  p_O_DFFX1 desc1494(.D(n181),.CLK(clk_i),.Q(s_dvd[23:23]),.E(p_desc1494_p_O_DFFX1));
  p_O_DFFX1 desc1495(.D(n154),.CLK(clk_i),.Q(rmndr_o[23:23]),.E(p_desc1495_p_O_DFFX1));
  p_O_DFFX1 desc1496(.D(n180),.CLK(clk_i),.Q(s_dvd[24:24]),.E(p_desc1496_p_O_DFFX1));
  p_O_DFFX1 desc1497(.D(n153),.CLK(clk_i),.Q(rmndr_o[24:24]),.E(p_desc1497_p_O_DFFX1));
  p_O_DFFX1 desc1498(.D(n179),.CLK(clk_i),.Q(s_dvd[25:25]),.E(p_desc1498_p_O_DFFX1));
  p_O_DFFX1 desc1499(.D(n152),.CLK(clk_i),.Q(rmndr_o[25:25]),.E(p_desc1499_p_O_DFFX1));
  p_O_DFFX1 desc1500(.D(n178),.CLK(clk_i),.Q(s_dvd[26:26]),.E(p_desc1500_p_O_DFFX1));
  p_O_DFFX1 desc1501(.D(n204),.CLK(clk_i),.Q(qutnt_o[26:26]),.E(p_desc1501_p_O_DFFX1));
  p_O_DFFX1 desc1502(.D(n205),.CLK(clk_i),.Q(qutnt_o[25:25]),.E(p_desc1502_p_O_DFFX1));
  p_O_DFFX1 desc1503(.D(n206),.CLK(clk_i),.Q(qutnt_o[24:24]),.E(p_desc1503_p_O_DFFX1));
  p_O_DFFX1 desc1504(.D(n207),.CLK(clk_i),.Q(qutnt_o[23:23]),.E(p_desc1504_p_O_DFFX1));
  p_O_DFFX1 desc1505(.D(n208),.CLK(clk_i),.Q(qutnt_o[22:22]),.E(p_desc1505_p_O_DFFX1));
  p_O_DFFX1 desc1506(.D(n209),.CLK(clk_i),.Q(qutnt_o[21:21]),.E(p_desc1506_p_O_DFFX1));
  p_O_DFFX1 desc1507(.D(n210),.CLK(clk_i),.Q(qutnt_o[20:20]),.E(p_desc1507_p_O_DFFX1));
  p_O_DFFX1 desc1508(.D(n211),.CLK(clk_i),.Q(qutnt_o[19:19]),.E(p_desc1508_p_O_DFFX1));
  p_O_DFFX1 desc1509(.D(n212),.CLK(clk_i),.Q(qutnt_o[18:18]),.E(p_desc1509_p_O_DFFX1));
  p_O_DFFX1 desc1510(.D(n213),.CLK(clk_i),.Q(qutnt_o[17:17]),.E(p_desc1510_p_O_DFFX1));
  p_O_DFFX1 desc1511(.D(n214),.CLK(clk_i),.Q(qutnt_o[16:16]),.E(p_desc1511_p_O_DFFX1));
  p_O_DFFX1 desc1512(.D(n215),.CLK(clk_i),.Q(qutnt_o[15:15]),.E(p_desc1512_p_O_DFFX1));
  p_O_DFFX1 desc1513(.D(n216),.CLK(clk_i),.Q(qutnt_o[14:14]),.E(p_desc1513_p_O_DFFX1));
  p_O_DFFX1 desc1514(.D(n217),.CLK(clk_i),.Q(qutnt_o[13:13]),.E(p_desc1514_p_O_DFFX1));
  p_O_DFFX1 desc1515(.D(n218),.CLK(clk_i),.Q(qutnt_o[12:12]),.E(p_desc1515_p_O_DFFX1));
  p_O_DFFX1 desc1516(.D(n219),.CLK(clk_i),.Q(qutnt_o[11:11]),.E(p_desc1516_p_O_DFFX1));
  p_O_DFFX1 desc1517(.D(n220),.CLK(clk_i),.Q(qutnt_o[10:10]),.E(p_desc1517_p_O_DFFX1));
  p_O_DFFX1 desc1518(.D(n221),.CLK(clk_i),.Q(qutnt_o[9:9]),.E(p_desc1518_p_O_DFFX1));
  p_O_DFFX1 desc1519(.D(n222),.CLK(clk_i),.Q(qutnt_o[8:8]),.E(p_desc1519_p_O_DFFX1));
  p_O_DFFX1 desc1520(.D(n223),.CLK(clk_i),.Q(qutnt_o[7:7]),.E(p_desc1520_p_O_DFFX1));
  p_O_DFFX1 desc1521(.D(n224),.CLK(clk_i),.Q(qutnt_o[6:6]),.E(p_desc1521_p_O_DFFX1));
  p_O_DFFX1 desc1522(.D(n225),.CLK(clk_i),.Q(qutnt_o[5:5]),.E(p_desc1522_p_O_DFFX1));
  p_O_DFFX1 desc1523(.D(n226),.CLK(clk_i),.Q(qutnt_o[4:4]),.E(p_desc1523_p_O_DFFX1));
  p_O_DFFX1 desc1524(.D(n227),.CLK(clk_i),.Q(qutnt_o[3:3]),.E(p_desc1524_p_O_DFFX1));
  p_O_DFFX1 desc1525(.D(n228),.CLK(clk_i),.Q(qutnt_o[2:2]),.E(p_desc1525_p_O_DFFX1));
  p_O_DFFX1 desc1526(.D(n229),.CLK(clk_i),.Q(qutnt_o[1:1]),.E(p_desc1526_p_O_DFFX1));
  p_O_DFFX1 desc1527(.D(n230),.CLK(clk_i),.Q(qutnt_o[0:0]),.E(p_desc1527_p_O_DFFX1));
  p_O_DFFX1 desc1528(.D(n151),.CLK(clk_i),.Q(rmndr_o[26:26]),.E(p_desc1528_p_O_DFFX1));
  XOR2X1 U50(.IN1(sign_dvd_i),.IN2(sign_div_i),.Q(sign_o));
  AO222X1 U51(.IN1(n45),.IN2(N186),.IN3(n46),.IN4(N158),.IN5(rmndr_o[26:26]),.IN6(n24),.Q(n151));
  AND2X1 U52(.IN1(n23),.IN2(N157),.Q(n46));
  AND2X1 U53(.IN1(n4),.IN2(n18),.Q(n45));
  AO22X1 U54(.IN1(rmndr_o[25:25]),.IN2(n24),.IN3(n23),.IN4(n50),.Q(n152));
  AO22X1 U55(.IN1(rmndr_o[24:24]),.IN2(n24),.IN3(n23),.IN4(n51),.Q(n153));
  AO22X1 U56(.IN1(rmndr_o[23:23]),.IN2(n24),.IN3(n22),.IN4(n52),.Q(n154));
  AO22X1 U57(.IN1(rmndr_o[22:22]),.IN2(n24),.IN3(n22),.IN4(n53),.Q(n155));
  AO22X1 U58(.IN1(rmndr_o[21:21]),.IN2(n24),.IN3(n22),.IN4(n54),.Q(n156));
  AO22X1 U59(.IN1(rmndr_o[20:20]),.IN2(n24),.IN3(n22),.IN4(n55),.Q(n157));
  AO22X1 U60(.IN1(rmndr_o[19:19]),.IN2(n24),.IN3(n22),.IN4(n56),.Q(n158));
  AO22X1 U61(.IN1(rmndr_o[18:18]),.IN2(n24),.IN3(n22),.IN4(n57),.Q(n159));
  AO22X1 U62(.IN1(rmndr_o[17:17]),.IN2(n24),.IN3(n22),.IN4(n58),.Q(n160));
  AO22X1 U63(.IN1(rmndr_o[16:16]),.IN2(n24),.IN3(n22),.IN4(n59),.Q(n161));
  AO22X1 U64(.IN1(rmndr_o[15:15]),.IN2(n24),.IN3(n22),.IN4(n60),.Q(n162));
  AO22X1 U65(.IN1(rmndr_o[14:14]),.IN2(n24),.IN3(n22),.IN4(n61),.Q(n163));
  AO22X1 U66(.IN1(rmndr_o[13:13]),.IN2(n24),.IN3(n22),.IN4(n62),.Q(n164));
  AO22X1 U67(.IN1(rmndr_o[12:12]),.IN2(n24),.IN3(n22),.IN4(n63),.Q(n165));
  AO22X1 U68(.IN1(rmndr_o[11:11]),.IN2(n24),.IN3(n21),.IN4(n64),.Q(n166));
  AO22X1 U69(.IN1(rmndr_o[10:10]),.IN2(n24),.IN3(n21),.IN4(n65),.Q(n167));
  AO22X1 U70(.IN1(rmndr_o[9:9]),.IN2(n24),.IN3(n21),.IN4(n66),.Q(n168));
  AO22X1 U71(.IN1(rmndr_o[8:8]),.IN2(n24),.IN3(n21),.IN4(n67),.Q(n169));
  AO22X1 U72(.IN1(rmndr_o[7:7]),.IN2(n24),.IN3(n21),.IN4(n68),.Q(n170));
  AO22X1 U73(.IN1(rmndr_o[6:6]),.IN2(n24),.IN3(n21),.IN4(n69),.Q(n171));
  AO22X1 U74(.IN1(rmndr_o[5:5]),.IN2(n24),.IN3(n21),.IN4(n70),.Q(n172));
  AO22X1 U75(.IN1(rmndr_o[4:4]),.IN2(n24),.IN3(n21),.IN4(n71),.Q(n173));
  AO22X1 U76(.IN1(rmndr_o[3:3]),.IN2(n24),.IN3(n21),.IN4(n72),.Q(n174));
  AO22X1 U77(.IN1(rmndr_o[2:2]),.IN2(n24),.IN3(n21),.IN4(n73),.Q(n175));
  AO22X1 U78(.IN1(rmndr_o[1:1]),.IN2(n24),.IN3(n21),.IN4(n74),.Q(n176));
  AO22X1 U79(.IN1(rmndr_o[0:0]),.IN2(n24),.IN3(n21),.IN4(n75),.Q(n177));
  AO22X1 U80(.IN1(s_dvd[26:26]),.IN2(n15),.IN3(n16),.IN4(n50),.Q(n178));
  AO22X1 U81(.IN1(N185),.IN2(n25),.IN3(N156),.IN4(N158),.Q(n50));
  AO22X1 U82(.IN1(s_dvd[25:25]),.IN2(n15),.IN3(n17),.IN4(n51),.Q(n179));
  AO22X1 U83(.IN1(N184),.IN2(n25),.IN3(N155),.IN4(N158),.Q(n51));
  AO22X1 U84(.IN1(s_dvd[24:24]),.IN2(n15),.IN3(n17),.IN4(n52),.Q(n180));
  AO22X1 U85(.IN1(N183),.IN2(n25),.IN3(N158),.IN4(N154),.Q(n52));
  AO22X1 U86(.IN1(s_dvd[23:23]),.IN2(n15),.IN3(n17),.IN4(n53),.Q(n181));
  AO22X1 U87(.IN1(N182),.IN2(n25),.IN3(N158),.IN4(N153),.Q(n53));
  AO22X1 U88(.IN1(s_dvd[22:22]),.IN2(n15),.IN3(n17),.IN4(n54),.Q(n182));
  AO22X1 U89(.IN1(N181),.IN2(n25),.IN3(N158),.IN4(N152),.Q(n54));
  AO22X1 U90(.IN1(s_dvd[21:21]),.IN2(n15),.IN3(n17),.IN4(n55),.Q(n183));
  AO22X1 U91(.IN1(N180),.IN2(n25),.IN3(N158),.IN4(N151),.Q(n55));
  AO22X1 U92(.IN1(s_dvd[20:20]),.IN2(n15),.IN3(n17),.IN4(n56),.Q(n184));
  AO22X1 U93(.IN1(N179),.IN2(n26),.IN3(N158),.IN4(N150),.Q(n56));
  AO22X1 U94(.IN1(s_dvd[19:19]),.IN2(n15),.IN3(n17),.IN4(n57),.Q(n185));
  AO22X1 U95(.IN1(N178),.IN2(n26),.IN3(N158),.IN4(N149),.Q(n57));
  AO22X1 U96(.IN1(s_dvd[18:18]),.IN2(n14),.IN3(n17),.IN4(n58),.Q(n186));
  AO22X1 U97(.IN1(N177),.IN2(n26),.IN3(N158),.IN4(N148),.Q(n58));
  AO22X1 U98(.IN1(s_dvd[17:17]),.IN2(n14),.IN3(n17),.IN4(n59),.Q(n187));
  AO22X1 U99(.IN1(N176),.IN2(n26),.IN3(N158),.IN4(N147),.Q(n59));
  AO22X1 U100(.IN1(s_dvd[16:16]),.IN2(n14),.IN3(n17),.IN4(n60),.Q(n188));
  AO22X1 U101(.IN1(N175),.IN2(n26),.IN3(N158),.IN4(N146),.Q(n60));
  AO22X1 U102(.IN1(s_dvd[15:15]),.IN2(n14),.IN3(n17),.IN4(n61),.Q(n189));
  AO22X1 U103(.IN1(N174),.IN2(n26),.IN3(N158),.IN4(N145),.Q(n61));
  AO22X1 U104(.IN1(s_dvd[14:14]),.IN2(n14),.IN3(n17),.IN4(n62),.Q(n190));
  AO22X1 U105(.IN1(N173),.IN2(n26),.IN3(N158),.IN4(N144),.Q(n62));
  AO22X1 U106(.IN1(s_dvd[13:13]),.IN2(n14),.IN3(n17),.IN4(n63),.Q(n191));
  AO22X1 U107(.IN1(N172),.IN2(n26),.IN3(N158),.IN4(N143),.Q(n63));
  AO22X1 U108(.IN1(s_dvd[12:12]),.IN2(n14),.IN3(n16),.IN4(n64),.Q(n192));
  AO22X1 U109(.IN1(N171),.IN2(n26),.IN3(N158),.IN4(N142),.Q(n64));
  AO22X1 U110(.IN1(s_dvd[11:11]),.IN2(n13),.IN3(n16),.IN4(n65),.Q(n193));
  AO22X1 U111(.IN1(N170),.IN2(n26),.IN3(N158),.IN4(N141),.Q(n65));
  AO22X1 U112(.IN1(s_dvd[10:10]),.IN2(n13),.IN3(n16),.IN4(n66),.Q(n194));
  AO22X1 U113(.IN1(N169),.IN2(n26),.IN3(N158),.IN4(N140),.Q(n66));
  AO22X1 U114(.IN1(s_dvd[9:9]),.IN2(n13),.IN3(n16),.IN4(n67),.Q(n195));
  AO22X1 U115(.IN1(N168),.IN2(n26),.IN3(N158),.IN4(N139),.Q(n67));
  AO22X1 U116(.IN1(s_dvd[8:8]),.IN2(n13),.IN3(n16),.IN4(n68),.Q(n196));
  AO22X1 U117(.IN1(N167),.IN2(n26),.IN3(N158),.IN4(N138),.Q(n68));
  AO22X1 U118(.IN1(s_dvd[7:7]),.IN2(n13),.IN3(n16),.IN4(n69),.Q(n197));
  AO22X1 U119(.IN1(N166),.IN2(n26),.IN3(N158),.IN4(N137),.Q(n69));
  AO22X1 U120(.IN1(s_dvd[6:6]),.IN2(n13),.IN3(n16),.IN4(n70),.Q(n198));
  AO22X1 U121(.IN1(N165),.IN2(n26),.IN3(N158),.IN4(N136),.Q(n70));
  AO22X1 U122(.IN1(s_dvd[5:5]),.IN2(n13),.IN3(n16),.IN4(n71),.Q(n199));
  AO22X1 U123(.IN1(N164),.IN2(n26),.IN3(N158),.IN4(N135),.Q(n71));
  AO22X1 U124(.IN1(s_dvd[4:4]),.IN2(n12),.IN3(n16),.IN4(n72),.Q(n200));
  AO22X1 U125(.IN1(N163),.IN2(n26),.IN3(N158),.IN4(N134),.Q(n72));
  AO22X1 U126(.IN1(s_dvd[3:3]),.IN2(n12),.IN3(n16),.IN4(n73),.Q(n201));
  AO22X1 U127(.IN1(N162),.IN2(n26),.IN3(N158),.IN4(N133),.Q(n73));
  AO22X1 U128(.IN1(s_dvd[2:2]),.IN2(n12),.IN3(n16),.IN4(n74),.Q(n202));
  AO22X1 U129(.IN1(N161),.IN2(n26),.IN3(N158),.IN4(N132),.Q(n74));
  AO22X1 U130(.IN1(s_dvd[1:1]),.IN2(n12),.IN3(n16),.IN4(n75),.Q(n203));
  AO22X1 U131(.IN1(N160),.IN2(n26),.IN3(N158),.IN4(n5),.Q(n75));
  AO22X1 U132(.IN1(n18),.IN2(n77),.IN3(qutnt_o[26:26]),.IN4(n36),.Q(n204));
  AO21X1 U133(.IN1(s_state),.IN2(n11),.IN3(n27),.Q(n77));
  AO22X1 U134(.IN1(n18),.IN2(n78),.IN3(qutnt_o[25:25]),.IN4(n35),.Q(n205));
  NAND3X0 U135(.IN1(s_count[4:4]),.IN2(s_count[3:3]),.IN3(n80),.QN(n79));
  AO22X1 U136(.IN1(n18),.IN2(n81),.IN3(qutnt_o[24:24]),.IN4(n34),.Q(n206));
  NAND3X0 U137(.IN1(s_count[4:4]),.IN2(s_count[3:3]),.IN3(n83),.QN(n82));
  AO22X1 U138(.IN1(n18),.IN2(n84),.IN3(qutnt_o[23:23]),.IN4(n37),.Q(n207));
  AO21X1 U139(.IN1(n85),.IN2(n86),.IN3(n27),.Q(n84));
  AO22X1 U140(.IN1(n18),.IN2(n87),.IN3(qutnt_o[22:22]),.IN4(n39),.Q(n208));
  AO21X1 U141(.IN1(n88),.IN2(n85),.IN3(n27),.Q(n87));
  AO22X1 U142(.IN1(n18),.IN2(n89),.IN3(qutnt_o[21:21]),.IN4(n40),.Q(n209));
  AO21X1 U143(.IN1(n90),.IN2(n85),.IN3(n27),.Q(n89));
  AO22X1 U144(.IN1(n18),.IN2(n91),.IN3(qutnt_o[20:20]),.IN4(n47),.Q(n210));
  AO21X1 U145(.IN1(n92),.IN2(n85),.IN3(n27),.Q(n91));
  AO22X1 U146(.IN1(n18),.IN2(n93),.IN3(qutnt_o[19:19]),.IN4(n238),.Q(n211));
  AO21X1 U147(.IN1(n94),.IN2(n85),.IN3(n27),.Q(n93));
  AO22X1 U148(.IN1(n18),.IN2(n95),.IN3(qutnt_o[18:18]),.IN4(n239),.Q(n212));
  AO21X1 U149(.IN1(n96),.IN2(n85),.IN3(n27),.Q(n95));
  AO22X1 U150(.IN1(n18),.IN2(n97),.IN3(qutnt_o[17:17]),.IN4(n240),.Q(n213));
  AO21X1 U151(.IN1(n85),.IN2(n80),.IN3(n27),.Q(n97));
  AO22X1 U152(.IN1(n18),.IN2(n98),.IN3(qutnt_o[16:16]),.IN4(n241),.Q(n214));
  AO21X1 U153(.IN1(n85),.IN2(n83),.IN3(n27),.Q(n98));
  AND2X1 U154(.IN1(s_count[4:4]),.IN2(n41),.Q(n85));
  AO22X1 U155(.IN1(n18),.IN2(n99),.IN3(qutnt_o[15:15]),.IN4(n242),.Q(n215));
  AO21X1 U156(.IN1(n100),.IN2(n86),.IN3(n27),.Q(n99));
  AO22X1 U157(.IN1(n19),.IN2(n101),.IN3(qutnt_o[14:14]),.IN4(n243),.Q(n216));
  AO21X1 U158(.IN1(n100),.IN2(n88),.IN3(n27),.Q(n101));
  AO22X1 U159(.IN1(n19),.IN2(n102),.IN3(qutnt_o[13:13]),.IN4(n244),.Q(n217));
  AO21X1 U160(.IN1(n100),.IN2(n90),.IN3(n27),.Q(n102));
  AO22X1 U161(.IN1(n19),.IN2(n103),.IN3(qutnt_o[12:12]),.IN4(n245),.Q(n218));
  AO21X1 U162(.IN1(n100),.IN2(n92),.IN3(n27),.Q(n103));
  AO22X1 U163(.IN1(n19),.IN2(n104),.IN3(qutnt_o[11:11]),.IN4(n246),.Q(n219));
  AO21X1 U164(.IN1(n100),.IN2(n94),.IN3(n27),.Q(n104));
  AO22X1 U165(.IN1(n19),.IN2(n105),.IN3(qutnt_o[10:10]),.IN4(n247),.Q(n220));
  AO21X1 U166(.IN1(n100),.IN2(n96),.IN3(n27),.Q(n105));
  AO22X1 U167(.IN1(n19),.IN2(n106),.IN3(qutnt_o[9:9]),.IN4(n248),.Q(n221));
  AO21X1 U168(.IN1(n100),.IN2(n80),.IN3(n27),.Q(n106));
  AO22X1 U169(.IN1(n19),.IN2(n107),.IN3(qutnt_o[8:8]),.IN4(n249),.Q(n222));
  AO21X1 U170(.IN1(n100),.IN2(n83),.IN3(n27),.Q(n107));
  AO22X1 U171(.IN1(n19),.IN2(n108),.IN3(qutnt_o[7:7]),.IN4(n250),.Q(n223));
  AO21X1 U172(.IN1(n109),.IN2(n86),.IN3(n27),.Q(n108));
  AND2X1 U173(.IN1(n110),.IN2(s_count[0:0]),.Q(n86));
  AO22X1 U174(.IN1(n19),.IN2(n111),.IN3(qutnt_o[6:6]),.IN4(n251),.Q(n224));
  AO21X1 U175(.IN1(n109),.IN2(n88),.IN3(n27),.Q(n111));
  AND2X1 U176(.IN1(n110),.IN2(n44),.Q(n88));
  AND2X1 U177(.IN1(n112),.IN2(s_count[1:1]),.Q(n110));
  AO22X1 U178(.IN1(n19),.IN2(n113),.IN3(qutnt_o[5:5]),.IN4(n252),.Q(n225));
  AO21X1 U179(.IN1(n109),.IN2(n90),.IN3(n27),.Q(n113));
  AND2X1 U180(.IN1(n114),.IN2(s_count[0:0]),.Q(n90));
  AO22X1 U181(.IN1(n19),.IN2(n115),.IN3(qutnt_o[4:4]),.IN4(n253),.Q(n226));
  AO21X1 U182(.IN1(n109),.IN2(n92),.IN3(n27),.Q(n115));
  AND2X1 U183(.IN1(n114),.IN2(n44),.Q(n92));
  AND2X1 U184(.IN1(n112),.IN2(n43),.Q(n114));
  AND2X1 U185(.IN1(s_count[2:2]),.IN2(s_state),.Q(n112));
  AO22X1 U186(.IN1(n19),.IN2(n116),.IN3(qutnt_o[3:3]),.IN4(n254),.Q(n227));
  AO21X1 U187(.IN1(n109),.IN2(n94),.IN3(n27),.Q(n116));
  AND4X1 U188(.IN1(s_count[0:0]),.IN2(s_state),.IN3(s_count[1:1]),.IN4(n42),.Q(n94));
  AO22X1 U189(.IN1(n19),.IN2(n117),.IN3(qutnt_o[2:2]),.IN4(n255),.Q(n228));
  AO21X1 U190(.IN1(n109),.IN2(n96),.IN3(n27),.Q(n117));
  AND2X1 U191(.IN1(s_state),.IN2(n118),.Q(n96));
  AO22X1 U192(.IN1(n20),.IN2(n119),.IN3(qutnt_o[1:1]),.IN4(n256),.Q(n229));
  AO21X1 U193(.IN1(n109),.IN2(n80),.IN3(n27),.Q(n119));
  AND4X1 U194(.IN1(s_count[0:0]),.IN2(s_state),.IN3(n43),.IN4(n42),.Q(n80));
  AO22X1 U195(.IN1(n20),.IN2(n120),.IN3(qutnt_o[0:0]),.IN4(n33),.Q(n230));
  AO221X1 U196(.IN1(n24),.IN2(s_count[3:3]),.IN3(N112),.IN4(n4),.IN5(n120),.Q(n231));
  AO22X1 U197(.IN1(s_count[2:2]),.IN2(n24),.IN3(N111),.IN4(n121),.Q(n232));
  AO221X1 U198(.IN1(n24),.IN2(s_count[1:1]),.IN3(N110),.IN4(n4),.IN5(n120),.Q(n233));
  AO22X1 U199(.IN1(n257),.IN2(n38),.IN3(ready_o),.IN4(n4),.Q(n234));
  AO21X1 U200(.IN1(s_state),.IN2(n122),.IN3(n27),.Q(n235));
  AO221X1 U201(.IN1(n24),.IN2(s_count[4:4]),.IN3(N113),.IN4(n4),.IN5(n120),.Q(n236));
  AO22X1 U202(.IN1(s_count[0:0]),.IN2(n24),.IN3(n44),.IN4(n121),.Q(n237));
  NOR3X0 U203(.IN1(n257),.IN2(n27),.IN3(n24),.QN(n121));
  AND4X1 U204(.IN1(s_state),.IN2(n44),.IN3(n43),.IN4(n42),.Q(n83));
  AND2X1 U205(.IN1(s_dvd[26:26]),.IN2(n6),.Q(N157));
  AND2X1 U206(.IN1(s_dvd[25:25]),.IN2(n6),.Q(N156));
  AND2X1 U207(.IN1(s_dvd[24:24]),.IN2(n6),.Q(N155));
  AO22X1 U208(.IN1(s_dvd[23:23]),.IN2(n6),.IN3(s_dvdnd_i[49:49]),.IN4(n11),.Q(N154));
  AO22X1 U209(.IN1(s_dvd[22:22]),.IN2(n10),.IN3(s_dvdnd_i[48:48]),.IN4(n11),.Q(N153));
  AO22X1 U210(.IN1(s_dvd[21:21]),.IN2(n10),.IN3(s_dvdnd_i[47:47]),.IN4(n11),.Q(N152));
  AO22X1 U211(.IN1(s_dvd[20:20]),.IN2(n10),.IN3(s_dvdnd_i[46:46]),.IN4(n11),.Q(N151));
  AO22X1 U212(.IN1(s_dvd[19:19]),.IN2(n10),.IN3(s_dvdnd_i[45:45]),.IN4(n11),.Q(N150));
  AO22X1 U213(.IN1(s_dvd[18:18]),.IN2(n10),.IN3(s_dvdnd_i[44:44]),.IN4(n11),.Q(N149));
  AO22X1 U214(.IN1(s_dvd[17:17]),.IN2(n10),.IN3(s_dvdnd_i[43:43]),.IN4(n11),.Q(N148));
  AO22X1 U215(.IN1(s_dvd[16:16]),.IN2(n9),.IN3(s_dvdnd_i[42:42]),.IN4(n11),.Q(N147));
  AO22X1 U216(.IN1(s_dvd[15:15]),.IN2(n9),.IN3(s_dvdnd_i[41:41]),.IN4(n11),.Q(N146));
  AO22X1 U217(.IN1(s_dvd[14:14]),.IN2(n9),.IN3(s_dvdnd_i[40:40]),.IN4(n11),.Q(N145));
  AO22X1 U218(.IN1(s_dvd[13:13]),.IN2(n9),.IN3(s_dvdnd_i[39:39]),.IN4(n11),.Q(N144));
  AO22X1 U219(.IN1(s_dvd[12:12]),.IN2(n9),.IN3(s_dvdnd_i[38:38]),.IN4(n11),.Q(N143));
  AO22X1 U220(.IN1(s_dvd[11:11]),.IN2(n9),.IN3(s_dvdnd_i[37:37]),.IN4(n11),.Q(N142));
  AO22X1 U221(.IN1(s_dvd[10:10]),.IN2(n7),.IN3(s_dvdnd_i[36:36]),.IN4(n11),.Q(N141));
  AO22X1 U222(.IN1(s_dvd[9:9]),.IN2(n7),.IN3(s_dvdnd_i[35:35]),.IN4(n11),.Q(N140));
  AO22X1 U223(.IN1(s_dvd[8:8]),.IN2(n7),.IN3(s_dvdnd_i[34:34]),.IN4(n11),.Q(N139));
  AO22X1 U224(.IN1(s_dvd[7:7]),.IN2(n7),.IN3(s_dvdnd_i[33:33]),.IN4(n11),.Q(N138));
  AO22X1 U225(.IN1(s_dvd[6:6]),.IN2(n9),.IN3(s_dvdnd_i[32:32]),.IN4(n11),.Q(N137));
  AO22X1 U226(.IN1(s_dvd[5:5]),.IN2(n7),.IN3(s_dvdnd_i[31:31]),.IN4(n11),.Q(N136));
  AO22X1 U227(.IN1(s_dvd[4:4]),.IN2(n7),.IN3(s_dvdnd_i[30:30]),.IN4(n11),.Q(N135));
  AO22X1 U228(.IN1(s_dvd[3:3]),.IN2(n7),.IN3(s_dvdnd_i[29:29]),.IN4(n11),.Q(N134));
  AO22X1 U229(.IN1(s_dvd[2:2]),.IN2(n6),.IN3(s_dvdnd_i[28:28]),.IN4(n11),.Q(N133));
  AO22X1 U230(.IN1(s_dvd[1:1]),.IN2(n6),.IN3(s_dvdnd_i[27:27]),.IN4(n11),.Q(N132));
  NAND3X0 U232(.IN1(s_count[3:3]),.IN2(n118),.IN3(s_count[4:4]),.QN(n123));
  NOR3X0 U233(.IN1(s_count[0:0]),.IN2(s_count[2:2]),.IN3(n43),.QN(n118));
  AND4X1 U234(.IN1(n124),.IN2(n125),.IN3(n126),.IN4(n127),.Q(N102));
  NOR4X0 U235(.IN1(n128),.IN2(s_dvsor_i[3:3]),.IN3(s_dvsor_i[5:5]),.IN4(s_dvsor_i[4:4]),.QN(n127));
  OR4X1 U236(.IN1(s_dvsor_i[7:7]),.IN2(s_dvsor_i[6:6]),.IN3(s_dvsor_i[9:9]),.IN4(s_dvsor_i[8:8]),.Q(n128));
  NOR4X0 U237(.IN1(n129),.IN2(s_dvsor_i[21:21]),.IN3(s_dvsor_i[23:23]),.IN4(s_dvsor_i[22:22]),.QN(n126));
  OR4X1 U238(.IN1(s_dvsor_i[25:25]),.IN2(s_dvsor_i[24:24]),.IN3(s_dvsor_i[2:2]),.IN4(s_dvsor_i[26:26]),.Q(n129));
  NOR4X0 U239(.IN1(n130),.IN2(s_dvsor_i[15:15]),.IN3(s_dvsor_i[17:17]),.IN4(s_dvsor_i[16:16]),.QN(n125));
  OR4X1 U240(.IN1(s_dvsor_i[19:19]),.IN2(s_dvsor_i[18:18]),.IN3(s_dvsor_i[20:20]),.IN4(s_dvsor_i[1:1]),.Q(n130));
  NOR4X0 U241(.IN1(n131),.IN2(n132),.IN3(s_dvsor_i[10:10]),.IN4(s_dvsor_i[0:0]),.QN(n124));
  NOR4X0 U242(.IN1(n133),.IN2(n134),.IN3(n135),.IN4(n136),.QN(n132));
  OR4X1 U243(.IN1(s_dvdnd_i[33:33]),.IN2(s_dvdnd_i[34:34]),.IN3(s_dvdnd_i[32:32]),.IN4(n137),.Q(n136));
  OR3X1 U244(.IN1(s_dvdnd_i[35:35]),.IN2(s_dvdnd_i[37:37]),.IN3(s_dvdnd_i[36:36]),.Q(n137));
  OR4X1 U245(.IN1(s_dvdnd_i[41:41]),.IN2(s_dvdnd_i[42:42]),.IN3(s_dvdnd_i[40:40]),.IN4(n138),.Q(n135));
  OR3X1 U246(.IN1(s_dvdnd_i[38:38]),.IN2(s_dvdnd_i[3:3]),.IN3(s_dvdnd_i[39:39]),.Q(n138));
  NAND4X0 U247(.IN1(n139),.IN2(n8),.IN3(n140),.IN4(n141),.QN(n134));
  NOR4X0 U248(.IN1(n142),.IN2(s_dvdnd_i[43:43]),.IN3(s_dvdnd_i[45:45]),.IN4(s_dvdnd_i[44:44]),.QN(n141));
  OR3X1 U249(.IN1(s_dvdnd_i[47:47]),.IN2(s_dvdnd_i[48:48]),.IN3(s_dvdnd_i[46:46]),.Q(n142));
  NOR4X0 U250(.IN1(s_dvdnd_i[9:9]),.IN2(s_dvdnd_i[8:8]),.IN3(s_dvdnd_i[7:7]),.IN4(s_dvdnd_i[6:6]),.QN(n140));
  NAND4X0 U251(.IN1(n143),.IN2(n144),.IN3(n145),.IN4(n146),.QN(n133));
  NOR4X0 U252(.IN1(n147),.IN2(s_dvdnd_i[26:26]),.IN3(s_dvdnd_i[28:28]),.IN4(s_dvdnd_i[27:27]),.QN(n146));
  OR4X1 U253(.IN1(s_dvdnd_i[2:2]),.IN2(s_dvdnd_i[29:29]),.IN3(s_dvdnd_i[31:31]),.IN4(s_dvdnd_i[30:30]),.Q(n147));
  NOR4X0 U254(.IN1(n148),.IN2(s_dvdnd_i[20:20]),.IN3(s_dvdnd_i[22:22]),.IN4(s_dvdnd_i[21:21]),.QN(n145));
  OR3X1 U255(.IN1(s_dvdnd_i[25:25]),.IN2(s_dvdnd_i[24:24]),.IN3(s_dvdnd_i[23:23]),.Q(n148));
  NOR4X0 U256(.IN1(n149),.IN2(s_dvdnd_i[15:15]),.IN3(s_dvdnd_i[17:17]),.IN4(s_dvdnd_i[16:16]),.QN(n144));
  OR3X1 U257(.IN1(s_dvdnd_i[1:1]),.IN2(s_dvdnd_i[19:19]),.IN3(s_dvdnd_i[18:18]),.Q(n149));
  NOR4X0 U258(.IN1(n150),.IN2(s_dvdnd_i[0:0]),.IN3(s_dvdnd_i[11:11]),.IN4(s_dvdnd_i[10:10]),.QN(n143));
  OR3X1 U259(.IN1(s_dvdnd_i[14:14]),.IN2(s_dvdnd_i[13:13]),.IN3(s_dvdnd_i[12:12]),.Q(n150));
  OR4X1 U260(.IN1(s_dvsor_i[12:12]),.IN2(s_dvsor_i[11:11]),.IN3(s_dvsor_i[14:14]),.IN4(s_dvsor_i[13:13]),.Q(n131));
  serial_div_DW01_sub_0_inj sub_154(.A({N157,N156,N155,N154,N153,N152,N151,N150,N149,N148,N147,N146,N145,N144,N143,N142,N141,N140,N139,N138,N137,N136,N135,N134,N133,N132,n5}),.B(s_dvsor_i),.CI(1'b0),.DIFF({N186,N185,N184,N183,N182,N181,N180,N179,N178,N177,N176,N175,N174,N173,N172,N171,N170,N169,N168,N167,N166,N165,N164,N163,N162,N161,N160}));
  serial_div_DW_cmp_0_inj lt_150(.A({N157,N156,N155,N154,N153,N152,N151,N150,N149,N148,N147,N146,N145,N144,N143,N142,N141,N140,N139,N138,N137,N136,N135,N134,N133,N132,n5}),.B(s_dvsor_i),.TC(1'b0),.GE_LT(1'b1),.GE_GT_EQ(1'b0),.GE_LT_GT_LE(N158));
  p_O_DFFX1 s_state_reg(.D(n235),.CLK(clk_i),.Q(s_state),.E(p_s_state_reg_p_O_DFFX1));
  p_O_DFFX1 desc1529(.D(n237),.CLK(clk_i),.Q(s_count[0:0]),.QN(n44),.E(p_desc1529_p_O_DFFX1));
  OR2X1 U3(.IN1(s_state),.IN2(n27),.Q(n4));
  INVX0 U4(.INP(n6),.ZN(n11));
  NBUFFX2 U5(.INP(n49),.Z(n18));
  NBUFFX2 U9(.INP(n49),.Z(n19));
  INVX0 U10(.INP(N158),.ZN(n25));
  NBUFFX2 U11(.INP(n49),.Z(n20));
  INVX0 U12(.INP(n4),.ZN(n24));
  NBUFFX2 U13(.INP(n48),.Z(n22));
  NBUFFX2 U14(.INP(n48),.Z(n21));
  INVX0 U15(.INP(N158),.ZN(n26));
  NBUFFX2 U16(.INP(n48),.Z(n23));
  INVX0 U17(.INP(n122),.ZN(n257));
  NBUFFX2 U18(.INP(n123),.Z(n6));
  NBUFFX2 U19(.INP(n123),.Z(n7));
  NBUFFX2 U20(.INP(n123),.Z(n9));
  NOR2X0 U21(.IN1(N158),.IN2(n27),.QN(n49));
  NBUFFX2 U22(.INP(n123),.Z(n10));
  NOR2X0 U23(.IN1(n24),.IN2(n27),.QN(n48));
  NBUFFX2 U24(.INP(n76),.Z(n12));
  NAND2X1 U25(.IN1(n109),.IN2(n83),.QN(n122));
  INVX0 U26(.INP(n29),.ZN(n32));
  INVX0 U27(.INP(n28),.ZN(n31));
  NBUFFX2 U28(.INP(n76),.Z(n15));
  NBUFFX2 U29(.INP(n76),.Z(n14));
  NBUFFX2 U30(.INP(n76),.Z(n13));
  NOR2X0 U31(.IN1(s_dvdnd_i[5:5]),.IN2(s_dvdnd_i[4:4]),.QN(n139));
  AND2X1 U32(.IN1(s_dvdnd_i[26:26]),.IN2(n11),.Q(n5));
  INVX0 U33(.INP(n99),.ZN(n242));
  INVX0 U34(.INP(n98),.ZN(n241));
  INVX0 U35(.INP(n97),.ZN(n240));
  INVX0 U36(.INP(n95),.ZN(n239));
  INVX0 U37(.INP(n93),.ZN(n238));
  INVX0 U38(.INP(n91),.ZN(n47));
  INVX0 U39(.INP(n89),.ZN(n40));
  INVX0 U40(.INP(n87),.ZN(n39));
  INVX0 U41(.INP(n84),.ZN(n37));
  INVX0 U42(.INP(n81),.ZN(n34));
  NAND2X1 U43(.IN1(n38),.IN2(n82),.QN(n81));
  INVX0 U44(.INP(n78),.ZN(n35));
  NAND2X1 U45(.IN1(n38),.IN2(n79),.QN(n78));
  INVX0 U46(.INP(n77),.ZN(n36));
  INVX0 U47(.INP(n117),.ZN(n255));
  INVX0 U48(.INP(n116),.ZN(n254));
  INVX0 U49(.INP(n115),.ZN(n253));
  INVX0 U231(.INP(n113),.ZN(n252));
  INVX0 U261(.INP(n111),.ZN(n251));
  INVX0 U262(.INP(n108),.ZN(n250));
  INVX0 U263(.INP(n107),.ZN(n249));
  INVX0 U264(.INP(n106),.ZN(n248));
  INVX0 U265(.INP(n105),.ZN(n247));
  INVX0 U266(.INP(n104),.ZN(n246));
  INVX0 U267(.INP(n103),.ZN(n245));
  INVX0 U268(.INP(n102),.ZN(n244));
  INVX0 U269(.INP(n101),.ZN(n243));
  INVX0 U270(.INP(n120),.ZN(n33));
  INVX0 U271(.INP(n119),.ZN(n256));
  NOR2X0 U272(.IN1(s_count[3:3]),.IN2(s_count[4:4]),.QN(n109));
  NAND2X1 U273(.IN1(n38),.IN2(n122),.QN(n120));
  NAND2X1 U274(.IN1(s_state),.IN2(n38),.QN(n76));
  NOR2X0 U275(.IN1(n41),.IN2(s_count[4:4]),.QN(n100));
  NBUFFX4 U276(.INP(s_start_i),.Z(n27));
  INVX0 U277(.INP(n12),.ZN(n16));
  INVX0 U278(.INP(n12),.ZN(n17));
  NOR2X0 U279(.IN1(s_count[1:1]),.IN2(s_count[0:0]),.QN(n28));
  AO21X1 U280(.IN1(s_count[1:1]),.IN2(s_count[0:0]),.IN3(n28),.Q(N110));
  NOR2X0 U281(.IN1(n31),.IN2(s_count[2:2]),.QN(n29));
  AO21X1 U282(.IN1(s_count[2:2]),.IN2(n31),.IN3(n29),.Q(N111));
  XNOR2X1 U283(.IN1(s_count[3:3]),.IN2(n32),.Q(N112));
  NOR2X0 U284(.IN1(s_count[3:3]),.IN2(n32),.QN(n30));
  XOR2X1 U285(.IN1(s_count[4:4]),.IN2(n30),.Q(N113));
assign div_zero_o=N102;
endmodule
module post_norm_div_DW01_inc_0_inj (A,SUM);
input [8:0] A ;
output [8:0] SUM ;
wire [8:2] carry ;
// instances
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[8:8]),.IN2(A[8:8]),.Q(SUM[8:8]));
endmodule
module post_norm_div_DW01_inc_1_inj (A,SUM);
input [24:0] A ;
output [24:0] SUM ;
wire [24:2] carry ;
// instances
  HADDX1 U1_1_23(.A0(A[23:23]),.B0(carry[23:23]),.C1(SUM[24:24]),.SO(SUM[23:23]));
  HADDX1 U1_1_22(.A0(A[22:22]),.B0(carry[22:22]),.C1(carry[23:23]),.SO(SUM[22:22]));
  HADDX1 U1_1_21(.A0(A[21:21]),.B0(carry[21:21]),.C1(carry[22:22]),.SO(SUM[21:21]));
  HADDX1 U1_1_20(.A0(A[20:20]),.B0(carry[20:20]),.C1(carry[21:21]),.SO(SUM[20:20]));
  HADDX1 U1_1_19(.A0(A[19:19]),.B0(carry[19:19]),.C1(carry[20:20]),.SO(SUM[19:19]));
  HADDX1 U1_1_18(.A0(A[18:18]),.B0(carry[18:18]),.C1(carry[19:19]),.SO(SUM[18:18]));
  HADDX1 U1_1_17(.A0(A[17:17]),.B0(carry[17:17]),.C1(carry[18:18]),.SO(SUM[17:17]));
  HADDX1 U1_1_16(.A0(A[16:16]),.B0(carry[16:16]),.C1(carry[17:17]),.SO(SUM[16:16]));
  HADDX1 U1_1_15(.A0(A[15:15]),.B0(carry[15:15]),.C1(carry[16:16]),.SO(SUM[15:15]));
  HADDX1 U1_1_14(.A0(A[14:14]),.B0(carry[14:14]),.C1(carry[15:15]),.SO(SUM[14:14]));
  HADDX1 U1_1_13(.A0(A[13:13]),.B0(carry[13:13]),.C1(carry[14:14]),.SO(SUM[13:13]));
  HADDX1 U1_1_12(.A0(A[12:12]),.B0(carry[12:12]),.C1(carry[13:13]),.SO(SUM[12:12]));
  HADDX1 U1_1_11(.A0(A[11:11]),.B0(carry[11:11]),.C1(carry[12:12]),.SO(SUM[11:11]));
  HADDX1 U1_1_10(.A0(A[10:10]),.B0(carry[10:10]),.C1(carry[11:11]),.SO(SUM[10:10]));
  HADDX1 U1_1_9(.A0(A[9:9]),.B0(carry[9:9]),.C1(carry[10:10]),.SO(SUM[9:9]));
  HADDX1 U1_1_8(.A0(A[8:8]),.B0(carry[8:8]),.C1(carry[9:9]),.SO(SUM[8:8]));
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
endmodule
module post_norm_div_inj (clk_i,opa_i,opb_i,qutnt_i,rmndr_i,exp_10_i,sign_i,rmode_i,output_o,ine_o,p_desc1530_p_O_DFFX1,p_desc1531_p_O_DFFX1,p_desc1532_p_O_DFFX1,p_desc1533_p_O_DFFX1,p_desc1534_p_O_DFFX1,p_desc1535_p_O_DFFX1,p_desc1536_p_O_DFFX1,p_desc1537_p_O_DFFX1,p_desc1538_p_O_DFFX1,p_desc1539_p_O_DFFX1,p_desc1540_p_O_DFFX1,p_desc1541_p_O_DFFX1,p_desc1542_p_O_DFFX1,p_desc1543_p_O_DFFX1,p_desc1544_p_O_DFFX1,p_desc1545_p_O_DFFX1,p_desc1546_p_O_DFFX1,p_desc1547_p_O_DFFX1,p_desc1548_p_O_DFFX1,p_desc1549_p_O_DFFX1,p_desc1550_p_O_DFFX1,p_desc1551_p_O_DFFX1,p_desc1552_p_O_DFFX1,p_desc1553_p_O_DFFX1,p_desc1554_p_O_DFFX1,p_desc1555_p_O_DFFX1,p_desc1556_p_O_DFFX1,p_desc1557_p_O_DFFX1,p_desc1558_p_O_DFFX1,p_desc1559_p_O_DFFX1,p_desc1560_p_O_DFFX1,p_desc1561_p_O_DFFX1,p_desc1562_p_O_DFFX1,p_desc1563_p_O_DFFX1,p_desc1564_p_O_DFFX1,p_desc1565_p_O_DFFX1,p_desc1566_p_O_DFFX1,p_desc1567_p_O_DFFX1,p_desc1568_p_O_DFFX1,p_desc1569_p_O_DFFX1,p_desc1570_p_O_DFFX1,p_desc1571_p_O_DFFX1,p_desc1572_p_O_DFFX1,p_desc1573_p_O_DFFX1,p_desc1574_p_O_DFFX1,p_desc1575_p_O_DFFX1,p_desc1576_p_O_DFFX1,p_desc1577_p_O_DFFX1,p_desc1578_p_O_DFFX1,p_desc1579_p_O_DFFX1,p_desc1580_p_O_DFFX1,p_desc1581_p_O_DFFX1,p_desc1582_p_O_DFFX1,p_desc1583_p_O_DFFX1,p_desc1584_p_O_DFFX1,p_desc1585_p_O_DFFX1,p_desc1586_p_O_DFFX1,p_desc1587_p_O_DFFX1,p_desc1588_p_O_DFFX1,p_desc1589_p_O_DFFX1,p_desc1590_p_O_DFFX1,p_desc1591_p_O_DFFX1,p_desc1592_p_O_DFFX1,p_desc1593_p_O_DFFX1,p_desc1594_p_O_DFFX1,p_desc1595_p_O_DFFX1,p_desc1596_p_O_DFFX1,p_desc1597_p_O_DFFX1,p_desc1598_p_O_DFFX1,p_desc1599_p_O_DFFX1,p_desc1600_p_O_DFFX1,p_desc1601_p_O_DFFX1,p_desc1602_p_O_DFFX1,p_desc1603_p_O_DFFX1,p_desc1604_p_O_DFFX1,p_desc1605_p_O_DFFX1,p_desc1606_p_O_DFFX1,p_desc1607_p_O_DFFX1,p_desc1608_p_O_DFFX1,p_desc1609_p_O_DFFX1,p_desc1610_p_O_DFFX1,p_desc1611_p_O_DFFX1,p_desc1612_p_O_DFFX1,p_desc1613_p_O_DFFX1,p_desc1614_p_O_DFFX1,p_desc1615_p_O_DFFX1,p_desc1616_p_O_DFFX1,p_desc1617_p_O_DFFX1,p_desc1618_p_O_DFFX1,p_desc1619_p_O_DFFX1,p_desc1620_p_O_DFFX1,p_desc1621_p_O_DFFX1,p_desc1622_p_O_DFFX1,p_desc1623_p_O_DFFX1,p_desc1624_p_O_DFFX1,p_desc1625_p_O_DFFX1,p_desc1626_p_O_DFFX1,p_desc1627_p_O_DFFX1,p_desc1628_p_O_DFFX1,p_desc1629_p_O_DFFX1,p_desc1630_p_O_DFFX1,p_desc1631_p_O_DFFX1,p_desc1632_p_O_DFFX1,p_desc1633_p_O_DFFX1,p_desc1634_p_O_DFFX1,p_desc1635_p_O_DFFX1,p_desc1636_p_O_DFFX1,p_desc1637_p_O_DFFX1,p_desc1638_p_O_DFFX1,p_desc1639_p_O_DFFX1,p_desc1640_p_O_DFFX1,p_desc1641_p_O_DFFX1,p_desc1642_p_O_DFFX1,p_desc1643_p_O_DFFX1,p_desc1644_p_O_DFFX1,p_desc1645_p_O_DFFX1,p_desc1646_p_O_DFFX1,p_desc1647_p_O_DFFX1,p_desc1648_p_O_DFFX1,p_desc1649_p_O_DFFX1,p_desc1650_p_O_DFFX1,p_desc1651_p_O_DFFX1,p_s_sign_i_reg_p_O_DFFX1,p_desc1652_p_O_DFFX1,p_desc1653_p_O_DFFX1,p_desc1654_p_O_DFFX1,p_desc1658_p_O_DFFX1,p_desc1659_p_O_DFFX1,p_desc1663_p_O_DFFX1,p_desc1664_p_O_DFFX1,p_desc1665_p_O_DFFX1,p_desc1666_p_O_DFFX1,p_desc1667_p_O_DFFX1,p_desc1668_p_O_DFFX1,p_desc1669_p_O_DFFX1,p_desc1670_p_O_DFFX1,p_desc1671_p_O_DFFX1,p_desc1672_p_O_DFFX1,p_desc1673_p_O_DFFX1,p_desc1674_p_O_DFFX1,p_desc1675_p_O_DFFX1,p_desc1676_p_O_DFFX1,p_desc1677_p_O_DFFX1,p_desc1678_p_O_DFFX1,p_desc1679_p_O_DFFX1,p_desc1680_p_O_DFFX1,p_desc1681_p_O_DFFX1,p_desc1682_p_O_DFFX1,p_desc1683_p_O_DFFX1,p_desc1684_p_O_DFFX1,p_desc1685_p_O_DFFX1,p_desc1686_p_O_DFFX1,p_desc1687_p_O_DFFX1,p_desc1688_p_O_DFFX1,p_desc1689_p_O_DFFX1,p_desc1690_p_O_DFFX1,p_desc1691_p_O_DFFX1,p_desc1692_p_O_DFFX1,p_desc1693_p_O_DFFX1,p_desc1694_p_O_DFFX1,p_desc1695_p_O_DFFX1,p_desc1696_p_O_DFFX1,p_desc1697_p_O_DFFX1,p_desc1698_p_O_DFFX1,p_desc1699_p_O_DFFX1,p_desc1700_p_O_DFFX1,p_desc1701_p_O_DFFX1,p_desc1702_p_O_DFFX1,p_desc1703_p_O_DFFX1,p_desc1704_p_O_DFFX1,p_desc1705_p_O_DFFX1,p_desc1706_p_O_DFFX1,p_desc1707_p_O_DFFX1,p_desc1708_p_O_DFFX1,p_desc1709_p_O_DFFX1,p_desc1710_p_O_DFFX1,p_desc1711_p_O_DFFX1,p_desc1712_p_O_DFFX1,p_desc1713_p_O_DFFX1,p_desc1714_p_O_DFFX1,p_desc1715_p_O_DFFX1,p_desc1716_p_O_DFFX1,p_desc1717_p_O_DFFX1,p_desc1718_p_O_DFFX1,p_desc1719_p_O_DFFX1,p_desc1720_p_O_DFFX1,p_desc1721_p_O_DFFX1,p_desc1722_p_O_DFFX1,p_desc1723_p_O_DFFX1,p_desc1724_p_O_DFFX1,p_desc1725_p_O_DFFX1,p_desc1726_p_O_DFFX1,p_desc1727_p_O_DFFX1,p_desc1728_p_O_DFFX1,p_ine_o_reg_p_O_DFFX1,p_desc1729_p_O_DFFX1,p_desc1737_p_O_DFFX1,p_desc1738_p_O_DFFX1,p_desc1739_p_O_DFFX1,p_desc1740_p_O_DFFX1,p_desc1741_p_O_DFFX1,p_desc1742_p_O_DFFX1,p_desc1743_p_O_DFFX1,p_desc1744_p_O_DFFX1,p_desc1745_p_O_DFFX1,p_desc1746_p_O_DFFX1,p_desc1747_p_O_DFFX1,p_desc1748_p_O_DFFX1,p_desc1749_p_O_DFFX1,p_desc1750_p_O_DFFX1,p_desc1751_p_O_DFFX1,p_desc1752_p_O_DFFX1,p_desc1753_p_O_DFFX1,p_desc1754_p_O_DFFX1,p_desc1755_p_O_DFFX1,p_desc1756_p_O_DFFX1,p_desc1757_p_O_DFFX1,p_desc1758_p_O_DFFX1,p_desc1849_p_O_DFFX1,p_desc1850_p_O_DFFX1,p_desc1851_p_O_DFFX1,p_desc1852_p_O_DFFX1,p_desc1853_p_O_DFFX1,p_desc1854_p_O_DFFX1,p_desc1855_p_O_DFFX1,p_desc1856_p_O_DFFX1,p_desc1857_p_O_DFFX1,p_desc1858_p_O_DFFX1,p_desc1859_p_O_DFFX1,p_desc1860_p_O_DFFX1,p_desc1861_p_O_DFFX1,p_desc1862_p_O_DFFX1,p_desc1863_p_O_DFFX1,p_desc1864_p_O_DFFX1,p_desc1865_p_O_DFFX1,p_desc1866_p_O_DFFX1,p_desc1867_p_O_DFFX1,p_desc1868_p_O_DFFX1,p_desc1869_p_O_DFFX1);
input [31:0] opa_i ;
input [31:0] opb_i ;
input [26:0] qutnt_i ;
input [26:0] rmndr_i ;
input [9:0] exp_10_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input clk_i ;
input sign_i ;
output ine_o ;
wire s_sign_i ;
wire \s_rmode_i[1]  ;
wire N145 ;
wire N146 ;
wire N147 ;
wire N148 ;
wire N149 ;
wire N150 ;
wire N151 ;
wire N161 ;
wire N162 ;
wire N166 ;
wire N167 ;
wire N172 ;
wire N173 ;
wire N174 ;
wire N175 ;
wire N176 ;
wire N177 ;
wire \s_shl1[0]  ;
wire N184 ;
wire N185 ;
wire N186 ;
wire N187 ;
wire N188 ;
wire N189 ;
wire N190 ;
wire N191 ;
wire N192 ;
wire N193 ;
wire N194 ;
wire N195 ;
wire N196 ;
wire N197 ;
wire N198 ;
wire N199 ;
wire N200 ;
wire N201 ;
wire N202 ;
wire N203 ;
wire N204 ;
wire N205 ;
wire N206 ;
wire N207 ;
wire N208 ;
wire N209 ;
wire N210 ;
wire N211 ;
wire N212 ;
wire N213 ;
wire N214 ;
wire N215 ;
wire N216 ;
wire N217 ;
wire N218 ;
wire N219 ;
wire N220 ;
wire N221 ;
wire N222 ;
wire N223 ;
wire N224 ;
wire N225 ;
wire N226 ;
wire N227 ;
wire N228 ;
wire N229 ;
wire N230 ;
wire N231 ;
wire N232 ;
wire N233 ;
wire N234 ;
wire N235 ;
wire N236 ;
wire N237 ;
wire N238 ;
wire N239 ;
wire N240 ;
wire N241 ;
wire N242 ;
wire N243 ;
wire N244 ;
wire N245 ;
wire N246 ;
wire N247 ;
wire N248 ;
wire N249 ;
wire N250 ;
wire N251 ;
wire N252 ;
wire N253 ;
wire N254 ;
wire N255 ;
wire N256 ;
wire N257 ;
wire N258 ;
wire N259 ;
wire N260 ;
wire N261 ;
wire N262 ;
wire N263 ;
wire N264 ;
wire N295 ;
wire N297 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N319 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N325 ;
wire N326 ;
wire N327 ;
wire N328 ;
wire N329 ;
wire N336 ;
wire N337 ;
wire N338 ;
wire N339 ;
wire N340 ;
wire N341 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N345 ;
wire N346 ;
wire N353 ;
wire N354 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N361 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N370 ;
wire N371 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N377 ;
wire N378 ;
wire N379 ;
wire N380 ;
wire N381 ;
wire N387 ;
wire N388 ;
wire N389 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N394 ;
wire N395 ;
wire N396 ;
wire N397 ;
wire N398 ;
wire N404 ;
wire N405 ;
wire N406 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N411 ;
wire N412 ;
wire N413 ;
wire N414 ;
wire N415 ;
wire N421 ;
wire N422 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N438 ;
wire N439 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N455 ;
wire N456 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N462 ;
wire N463 ;
wire N464 ;
wire N465 ;
wire N466 ;
wire N472 ;
wire N473 ;
wire N474 ;
wire N475 ;
wire N476 ;
wire N477 ;
wire N478 ;
wire N479 ;
wire N480 ;
wire N481 ;
wire N482 ;
wire N483 ;
wire N489 ;
wire N490 ;
wire N491 ;
wire N492 ;
wire N493 ;
wire N494 ;
wire N495 ;
wire N496 ;
wire N497 ;
wire N498 ;
wire N499 ;
wire N500 ;
wire N506 ;
wire N507 ;
wire N508 ;
wire N509 ;
wire N510 ;
wire N511 ;
wire N512 ;
wire N513 ;
wire N514 ;
wire N515 ;
wire N516 ;
wire N517 ;
wire N523 ;
wire N524 ;
wire N525 ;
wire N526 ;
wire N527 ;
wire N528 ;
wire N529 ;
wire N530 ;
wire N531 ;
wire N532 ;
wire N533 ;
wire N534 ;
wire N540 ;
wire N541 ;
wire N542 ;
wire N543 ;
wire N544 ;
wire N545 ;
wire N546 ;
wire N547 ;
wire N548 ;
wire N549 ;
wire N550 ;
wire N551 ;
wire N557 ;
wire N558 ;
wire N559 ;
wire N560 ;
wire N561 ;
wire N562 ;
wire N563 ;
wire N564 ;
wire N565 ;
wire N566 ;
wire N567 ;
wire N568 ;
wire N574 ;
wire N575 ;
wire N576 ;
wire N577 ;
wire N578 ;
wire N579 ;
wire N580 ;
wire N581 ;
wire N582 ;
wire N583 ;
wire N584 ;
wire N585 ;
wire N592 ;
wire N593 ;
wire N594 ;
wire N595 ;
wire N596 ;
wire N597 ;
wire N598 ;
wire N599 ;
wire N600 ;
wire N601 ;
wire N602 ;
wire N608 ;
wire N609 ;
wire N610 ;
wire N611 ;
wire N612 ;
wire N613 ;
wire N614 ;
wire N615 ;
wire N616 ;
wire N617 ;
wire N618 ;
wire N619 ;
wire N625 ;
wire N626 ;
wire N627 ;
wire N628 ;
wire N629 ;
wire N630 ;
wire N631 ;
wire N632 ;
wire N633 ;
wire N634 ;
wire N635 ;
wire N636 ;
wire N642 ;
wire N643 ;
wire N644 ;
wire N645 ;
wire N646 ;
wire N647 ;
wire N648 ;
wire N649 ;
wire N650 ;
wire N651 ;
wire N652 ;
wire N653 ;
wire N659 ;
wire N660 ;
wire N661 ;
wire N662 ;
wire N663 ;
wire N664 ;
wire N665 ;
wire N666 ;
wire N667 ;
wire N668 ;
wire N669 ;
wire N670 ;
wire N676 ;
wire N677 ;
wire N678 ;
wire N679 ;
wire N680 ;
wire N681 ;
wire N1019 ;
wire N1020 ;
wire N1021 ;
wire N1022 ;
wire N1023 ;
wire N1024 ;
wire N1025 ;
wire N1065 ;
wire N1066 ;
wire N1067 ;
wire N1068 ;
wire N1069 ;
wire N1070 ;
wire N1071 ;
wire N1072 ;
wire N1073 ;
wire N1074 ;
wire N1075 ;
wire N1076 ;
wire N1077 ;
wire N1078 ;
wire N1079 ;
wire N1080 ;
wire N1081 ;
wire N1082 ;
wire N1083 ;
wire N1084 ;
wire N1085 ;
wire N1086 ;
wire N1087 ;
wire N1088 ;
wire N1089 ;
wire N1091 ;
wire N1092 ;
wire N1093 ;
wire N1094 ;
wire N1095 ;
wire N1096 ;
wire N1097 ;
wire N1098 ;
wire N1099 ;
wire N1100 ;
wire N1101 ;
wire N1102 ;
wire N1103 ;
wire N1104 ;
wire N1105 ;
wire N1106 ;
wire N1107 ;
wire N1108 ;
wire N1109 ;
wire N1110 ;
wire N1111 ;
wire N1112 ;
wire N1113 ;
wire N1114 ;
wire N1115 ;
wire N1116 ;
wire N1117 ;
wire N1118 ;
wire N1119 ;
wire N1120 ;
wire N1121 ;
wire N1122 ;
wire N1123 ;
wire N1124 ;
wire N1125 ;
wire N1126 ;
wire N1127 ;
wire N1128 ;
wire N1129 ;
wire N1130 ;
wire N1131 ;
wire N1386 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n71 ;
wire n79 ;
wire n86 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n108 ;
wire n112 ;
wire n113 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire \add_194/carry[5]  ;
wire \add_194/carry[4]  ;
wire \add_194/carry[3]  ;
wire \add_194/carry[2]  ;
wire \add_194/carry[1]  ;
wire \add_194/B[0]  ;
wire \add_105_I27_L14036_C191/carry[5]  ;
wire \add_105_I27_L14036_C191/carry[4]  ;
wire \add_105_I27_L14036_C191/carry[3]  ;
wire \add_105_I27_L14036_C191/carry[2]  ;
wire \add_105_I26_L14036_C191/carry[5]  ;
wire \add_105_I26_L14036_C191/carry[4]  ;
wire \add_105_I26_L14036_C191/carry[3]  ;
wire \add_105_I26_L14036_C191/carry[2]  ;
wire \add_105_I25_L14036_C191/carry[5]  ;
wire \add_105_I25_L14036_C191/carry[4]  ;
wire \add_105_I25_L14036_C191/carry[3]  ;
wire \add_105_I25_L14036_C191/carry[2]  ;
wire \add_105_I24_L14036_C191/carry[5]  ;
wire \add_105_I24_L14036_C191/carry[4]  ;
wire \add_105_I24_L14036_C191/carry[3]  ;
wire \add_105_I24_L14036_C191/carry[2]  ;
wire \add_105_I23_L14036_C191/carry[5]  ;
wire \add_105_I23_L14036_C191/carry[4]  ;
wire \add_105_I23_L14036_C191/carry[3]  ;
wire \add_105_I23_L14036_C191/carry[2]  ;
wire \add_105_I22_L14036_C191/carry[5]  ;
wire \add_105_I22_L14036_C191/carry[4]  ;
wire \add_105_I22_L14036_C191/carry[3]  ;
wire \add_105_I22_L14036_C191/carry[2]  ;
wire \add_105_I21_L14036_C191/carry[5]  ;
wire \add_105_I21_L14036_C191/carry[4]  ;
wire \add_105_I21_L14036_C191/carry[3]  ;
wire \add_105_I21_L14036_C191/carry[2]  ;
wire \add_105_I20_L14036_C191/carry[5]  ;
wire \add_105_I20_L14036_C191/carry[4]  ;
wire \add_105_I20_L14036_C191/carry[3]  ;
wire \add_105_I20_L14036_C191/carry[2]  ;
wire \add_105_I19_L14036_C191/carry[5]  ;
wire \add_105_I19_L14036_C191/carry[4]  ;
wire \add_105_I19_L14036_C191/carry[3]  ;
wire \add_105_I19_L14036_C191/carry[2]  ;
wire \add_105_I18_L14036_C191/carry[5]  ;
wire \add_105_I18_L14036_C191/carry[4]  ;
wire \add_105_I18_L14036_C191/carry[3]  ;
wire \add_105_I18_L14036_C191/carry[2]  ;
wire \add_105_I17_L14036_C191/carry[5]  ;
wire \add_105_I17_L14036_C191/carry[4]  ;
wire \add_105_I17_L14036_C191/carry[3]  ;
wire \add_105_I17_L14036_C191/carry[2]  ;
wire \add_105_I16_L14036_C191/carry[5]  ;
wire \add_105_I16_L14036_C191/carry[4]  ;
wire \add_105_I16_L14036_C191/carry[3]  ;
wire \add_105_I16_L14036_C191/carry[2]  ;
wire \add_105_I15_L14036_C191/carry[5]  ;
wire \add_105_I15_L14036_C191/carry[4]  ;
wire \add_105_I15_L14036_C191/carry[3]  ;
wire \add_105_I15_L14036_C191/carry[2]  ;
wire \add_105_I14_L14036_C191/carry[5]  ;
wire \add_105_I14_L14036_C191/carry[4]  ;
wire \add_105_I14_L14036_C191/carry[3]  ;
wire \add_105_I14_L14036_C191/carry[2]  ;
wire \add_105_I13_L14036_C191/carry[5]  ;
wire \add_105_I13_L14036_C191/carry[4]  ;
wire \add_105_I13_L14036_C191/carry[3]  ;
wire \add_105_I13_L14036_C191/carry[2]  ;
wire \add_105_I12_L14036_C191/carry[5]  ;
wire \add_105_I12_L14036_C191/carry[4]  ;
wire \add_105_I12_L14036_C191/carry[3]  ;
wire \add_105_I12_L14036_C191/carry[2]  ;
wire \add_105_I11_L14036_C191/carry[5]  ;
wire \add_105_I11_L14036_C191/carry[4]  ;
wire \add_105_I11_L14036_C191/carry[3]  ;
wire \add_105_I11_L14036_C191/carry[2]  ;
wire \add_105_I10_L14036_C191/carry[5]  ;
wire \add_105_I10_L14036_C191/carry[4]  ;
wire \add_105_I10_L14036_C191/carry[3]  ;
wire \add_105_I10_L14036_C191/carry[2]  ;
wire \add_105_I9_L14036_C191/carry[5]  ;
wire \add_105_I9_L14036_C191/carry[4]  ;
wire \add_105_I9_L14036_C191/carry[3]  ;
wire \add_105_I9_L14036_C191/carry[2]  ;
wire \add_105_I8_L14036_C191/carry[5]  ;
wire \add_105_I8_L14036_C191/carry[4]  ;
wire \add_105_I8_L14036_C191/carry[3]  ;
wire \add_105_I8_L14036_C191/carry[2]  ;
wire \add_105_I7_L14036_C191/carry[4]  ;
wire \add_105_I7_L14036_C191/carry[3]  ;
wire \add_105_I7_L14036_C191/carry[2]  ;
wire \add_105_I6_L14036_C191/carry[2]  ;
wire \add_105_I6_L14036_C191/carry[3]  ;
wire \add_105_I5_L14036_C191/carry[2]  ;
wire \add_105_I5_L14036_C191/A[1]  ;
wire \sub_188_aco/carry[8]  ;
wire \sub_188_aco/carry[7]  ;
wire \sub_188_aco/carry[6]  ;
wire \sub_188_aco/carry[5]  ;
wire \sub_188_aco/carry[4]  ;
wire \sub_188_aco/carry[3]  ;
wire \sub_188_aco/carry[2]  ;
wire \sub_188_aco/carry[1]  ;
wire \sub_1_root_sub_150_2/carry[5]  ;
wire \sub_1_root_sub_150_2/carry[4]  ;
wire \sub_1_root_sub_150_2/carry[3]  ;
wire \sub_1_root_sub_150_2/carry[2]  ;
wire \sub_1_root_sub_150_2/carry[1]  ;
wire \sub_1_root_sub_150_2/CI  ;
wire \sub_141/carry[9]  ;
wire \sub_141/carry[8]  ;
wire \sub_141/carry[7]  ;
wire \sub_141/carry[6]  ;
wire \sub_141/carry[5]  ;
wire \sub_141/carry[4]  ;
wire \sub_141/carry[3]  ;
wire \sub_141/carry[2]  ;
wire \sub_141/carry[1]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n102 ;
wire n107 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n120 ;
wire n121 ;
wire n125 ;
wire n299 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n381 ;
wire n382 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n404 ;
wire n405 ;
wire n406 ;
wire n407 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n416 ;
wire n417 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire n429 ;
wire n430 ;
wire n431 ;
wire n432 ;
wire n433 ;
wire n434 ;
wire n435 ;
wire n436 ;
wire n437 ;
wire n438 ;
wire n439 ;
wire n440 ;
wire n441 ;
wire n442 ;
wire n443 ;
wire n444 ;
wire n445 ;
wire n446 ;
wire n447 ;
wire n448 ;
wire [30:0] s_opa_i ;
wire [30:0] s_opb_i ;
wire [7:0] s_expa ;
wire [7:0] s_expb ;
wire [26:0] s_qutnt_i ;
wire [26:0] s_rmndr_i ;
wire [9:0] s_exp_10_i ;
wire [31:0] s_output_o ;
wire [9:0] s_exp_10b ;
wire [8:0] s_expo1 ;
wire [5:0] s_shr1 ;
wire [26:0] s_fraco1 ;
wire [8:0] s_expo2 ;
wire [5:0] s_r_zeros ;
wire [8:0] s_expo3 ;
wire [22:0] s_fraco2 ;
input p_desc1530_p_O_DFFX1 ;
input p_desc1531_p_O_DFFX1 ;
input p_desc1532_p_O_DFFX1 ;
input p_desc1533_p_O_DFFX1 ;
input p_desc1534_p_O_DFFX1 ;
input p_desc1535_p_O_DFFX1 ;
input p_desc1536_p_O_DFFX1 ;
input p_desc1537_p_O_DFFX1 ;
input p_desc1538_p_O_DFFX1 ;
input p_desc1539_p_O_DFFX1 ;
input p_desc1540_p_O_DFFX1 ;
input p_desc1541_p_O_DFFX1 ;
input p_desc1542_p_O_DFFX1 ;
input p_desc1543_p_O_DFFX1 ;
input p_desc1544_p_O_DFFX1 ;
input p_desc1545_p_O_DFFX1 ;
input p_desc1546_p_O_DFFX1 ;
input p_desc1547_p_O_DFFX1 ;
input p_desc1548_p_O_DFFX1 ;
input p_desc1549_p_O_DFFX1 ;
input p_desc1550_p_O_DFFX1 ;
input p_desc1551_p_O_DFFX1 ;
input p_desc1552_p_O_DFFX1 ;
input p_desc1553_p_O_DFFX1 ;
input p_desc1554_p_O_DFFX1 ;
input p_desc1555_p_O_DFFX1 ;
input p_desc1556_p_O_DFFX1 ;
input p_desc1557_p_O_DFFX1 ;
input p_desc1558_p_O_DFFX1 ;
input p_desc1559_p_O_DFFX1 ;
input p_desc1560_p_O_DFFX1 ;
input p_desc1561_p_O_DFFX1 ;
input p_desc1562_p_O_DFFX1 ;
input p_desc1563_p_O_DFFX1 ;
input p_desc1564_p_O_DFFX1 ;
input p_desc1565_p_O_DFFX1 ;
input p_desc1566_p_O_DFFX1 ;
input p_desc1567_p_O_DFFX1 ;
input p_desc1568_p_O_DFFX1 ;
input p_desc1569_p_O_DFFX1 ;
input p_desc1570_p_O_DFFX1 ;
input p_desc1571_p_O_DFFX1 ;
input p_desc1572_p_O_DFFX1 ;
input p_desc1573_p_O_DFFX1 ;
input p_desc1574_p_O_DFFX1 ;
input p_desc1575_p_O_DFFX1 ;
input p_desc1576_p_O_DFFX1 ;
input p_desc1577_p_O_DFFX1 ;
input p_desc1578_p_O_DFFX1 ;
input p_desc1579_p_O_DFFX1 ;
input p_desc1580_p_O_DFFX1 ;
input p_desc1581_p_O_DFFX1 ;
input p_desc1582_p_O_DFFX1 ;
input p_desc1583_p_O_DFFX1 ;
input p_desc1584_p_O_DFFX1 ;
input p_desc1585_p_O_DFFX1 ;
input p_desc1586_p_O_DFFX1 ;
input p_desc1587_p_O_DFFX1 ;
input p_desc1588_p_O_DFFX1 ;
input p_desc1589_p_O_DFFX1 ;
input p_desc1590_p_O_DFFX1 ;
input p_desc1591_p_O_DFFX1 ;
input p_desc1592_p_O_DFFX1 ;
input p_desc1593_p_O_DFFX1 ;
input p_desc1594_p_O_DFFX1 ;
input p_desc1595_p_O_DFFX1 ;
input p_desc1596_p_O_DFFX1 ;
input p_desc1597_p_O_DFFX1 ;
input p_desc1598_p_O_DFFX1 ;
input p_desc1599_p_O_DFFX1 ;
input p_desc1600_p_O_DFFX1 ;
input p_desc1601_p_O_DFFX1 ;
input p_desc1602_p_O_DFFX1 ;
input p_desc1603_p_O_DFFX1 ;
input p_desc1604_p_O_DFFX1 ;
input p_desc1605_p_O_DFFX1 ;
input p_desc1606_p_O_DFFX1 ;
input p_desc1607_p_O_DFFX1 ;
input p_desc1608_p_O_DFFX1 ;
input p_desc1609_p_O_DFFX1 ;
input p_desc1610_p_O_DFFX1 ;
input p_desc1611_p_O_DFFX1 ;
input p_desc1612_p_O_DFFX1 ;
input p_desc1613_p_O_DFFX1 ;
input p_desc1614_p_O_DFFX1 ;
input p_desc1615_p_O_DFFX1 ;
input p_desc1616_p_O_DFFX1 ;
input p_desc1617_p_O_DFFX1 ;
input p_desc1618_p_O_DFFX1 ;
input p_desc1619_p_O_DFFX1 ;
input p_desc1620_p_O_DFFX1 ;
input p_desc1621_p_O_DFFX1 ;
input p_desc1622_p_O_DFFX1 ;
input p_desc1623_p_O_DFFX1 ;
input p_desc1624_p_O_DFFX1 ;
input p_desc1625_p_O_DFFX1 ;
input p_desc1626_p_O_DFFX1 ;
input p_desc1627_p_O_DFFX1 ;
input p_desc1628_p_O_DFFX1 ;
input p_desc1629_p_O_DFFX1 ;
input p_desc1630_p_O_DFFX1 ;
input p_desc1631_p_O_DFFX1 ;
input p_desc1632_p_O_DFFX1 ;
input p_desc1633_p_O_DFFX1 ;
input p_desc1634_p_O_DFFX1 ;
input p_desc1635_p_O_DFFX1 ;
input p_desc1636_p_O_DFFX1 ;
input p_desc1637_p_O_DFFX1 ;
input p_desc1638_p_O_DFFX1 ;
input p_desc1639_p_O_DFFX1 ;
input p_desc1640_p_O_DFFX1 ;
input p_desc1641_p_O_DFFX1 ;
input p_desc1642_p_O_DFFX1 ;
input p_desc1643_p_O_DFFX1 ;
input p_desc1644_p_O_DFFX1 ;
input p_desc1645_p_O_DFFX1 ;
input p_desc1646_p_O_DFFX1 ;
input p_desc1647_p_O_DFFX1 ;
input p_desc1648_p_O_DFFX1 ;
input p_desc1649_p_O_DFFX1 ;
input p_desc1650_p_O_DFFX1 ;
input p_desc1651_p_O_DFFX1 ;
input p_s_sign_i_reg_p_O_DFFX1 ;
input p_desc1652_p_O_DFFX1 ;
input p_desc1653_p_O_DFFX1 ;
input p_desc1654_p_O_DFFX1 ;
input p_desc1658_p_O_DFFX1 ;
input p_desc1659_p_O_DFFX1 ;
input p_desc1663_p_O_DFFX1 ;
input p_desc1664_p_O_DFFX1 ;
input p_desc1665_p_O_DFFX1 ;
input p_desc1666_p_O_DFFX1 ;
input p_desc1667_p_O_DFFX1 ;
input p_desc1668_p_O_DFFX1 ;
input p_desc1669_p_O_DFFX1 ;
input p_desc1670_p_O_DFFX1 ;
input p_desc1671_p_O_DFFX1 ;
input p_desc1672_p_O_DFFX1 ;
input p_desc1673_p_O_DFFX1 ;
input p_desc1674_p_O_DFFX1 ;
input p_desc1675_p_O_DFFX1 ;
input p_desc1676_p_O_DFFX1 ;
input p_desc1677_p_O_DFFX1 ;
input p_desc1678_p_O_DFFX1 ;
input p_desc1679_p_O_DFFX1 ;
input p_desc1680_p_O_DFFX1 ;
input p_desc1681_p_O_DFFX1 ;
input p_desc1682_p_O_DFFX1 ;
input p_desc1683_p_O_DFFX1 ;
input p_desc1684_p_O_DFFX1 ;
input p_desc1685_p_O_DFFX1 ;
input p_desc1686_p_O_DFFX1 ;
input p_desc1687_p_O_DFFX1 ;
input p_desc1688_p_O_DFFX1 ;
input p_desc1689_p_O_DFFX1 ;
input p_desc1690_p_O_DFFX1 ;
input p_desc1691_p_O_DFFX1 ;
input p_desc1692_p_O_DFFX1 ;
input p_desc1693_p_O_DFFX1 ;
input p_desc1694_p_O_DFFX1 ;
input p_desc1695_p_O_DFFX1 ;
input p_desc1696_p_O_DFFX1 ;
input p_desc1697_p_O_DFFX1 ;
input p_desc1698_p_O_DFFX1 ;
input p_desc1699_p_O_DFFX1 ;
input p_desc1700_p_O_DFFX1 ;
input p_desc1701_p_O_DFFX1 ;
input p_desc1702_p_O_DFFX1 ;
input p_desc1703_p_O_DFFX1 ;
input p_desc1704_p_O_DFFX1 ;
input p_desc1705_p_O_DFFX1 ;
input p_desc1706_p_O_DFFX1 ;
input p_desc1707_p_O_DFFX1 ;
input p_desc1708_p_O_DFFX1 ;
input p_desc1709_p_O_DFFX1 ;
input p_desc1710_p_O_DFFX1 ;
input p_desc1711_p_O_DFFX1 ;
input p_desc1712_p_O_DFFX1 ;
input p_desc1713_p_O_DFFX1 ;
input p_desc1714_p_O_DFFX1 ;
input p_desc1715_p_O_DFFX1 ;
input p_desc1716_p_O_DFFX1 ;
input p_desc1717_p_O_DFFX1 ;
input p_desc1718_p_O_DFFX1 ;
input p_desc1719_p_O_DFFX1 ;
input p_desc1720_p_O_DFFX1 ;
input p_desc1721_p_O_DFFX1 ;
input p_desc1722_p_O_DFFX1 ;
input p_desc1723_p_O_DFFX1 ;
input p_desc1724_p_O_DFFX1 ;
input p_desc1725_p_O_DFFX1 ;
input p_desc1726_p_O_DFFX1 ;
input p_desc1727_p_O_DFFX1 ;
input p_desc1728_p_O_DFFX1 ;
input p_ine_o_reg_p_O_DFFX1 ;
input p_desc1729_p_O_DFFX1 ;
input p_desc1737_p_O_DFFX1 ;
input p_desc1738_p_O_DFFX1 ;
input p_desc1739_p_O_DFFX1 ;
input p_desc1740_p_O_DFFX1 ;
input p_desc1741_p_O_DFFX1 ;
input p_desc1742_p_O_DFFX1 ;
input p_desc1743_p_O_DFFX1 ;
input p_desc1744_p_O_DFFX1 ;
input p_desc1745_p_O_DFFX1 ;
input p_desc1746_p_O_DFFX1 ;
input p_desc1747_p_O_DFFX1 ;
input p_desc1748_p_O_DFFX1 ;
input p_desc1749_p_O_DFFX1 ;
input p_desc1750_p_O_DFFX1 ;
input p_desc1751_p_O_DFFX1 ;
input p_desc1752_p_O_DFFX1 ;
input p_desc1753_p_O_DFFX1 ;
input p_desc1754_p_O_DFFX1 ;
input p_desc1755_p_O_DFFX1 ;
input p_desc1756_p_O_DFFX1 ;
input p_desc1757_p_O_DFFX1 ;
input p_desc1758_p_O_DFFX1 ;
input p_desc1849_p_O_DFFX1 ;
input p_desc1850_p_O_DFFX1 ;
input p_desc1851_p_O_DFFX1 ;
input p_desc1852_p_O_DFFX1 ;
input p_desc1853_p_O_DFFX1 ;
input p_desc1854_p_O_DFFX1 ;
input p_desc1855_p_O_DFFX1 ;
input p_desc1856_p_O_DFFX1 ;
input p_desc1857_p_O_DFFX1 ;
input p_desc1858_p_O_DFFX1 ;
input p_desc1859_p_O_DFFX1 ;
input p_desc1860_p_O_DFFX1 ;
input p_desc1861_p_O_DFFX1 ;
input p_desc1862_p_O_DFFX1 ;
input p_desc1863_p_O_DFFX1 ;
input p_desc1864_p_O_DFFX1 ;
input p_desc1865_p_O_DFFX1 ;
input p_desc1866_p_O_DFFX1 ;
input p_desc1867_p_O_DFFX1 ;
input p_desc1868_p_O_DFFX1 ;
input p_desc1869_p_O_DFFX1 ;
// instances
  p_O_DFFX1 desc1530(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_opa_i[30:30]),.E(p_desc1530_p_O_DFFX1));
  p_O_DFFX1 desc1531(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_opa_i[29:29]),.E(p_desc1531_p_O_DFFX1));
  p_O_DFFX1 desc1532(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_opa_i[28:28]),.E(p_desc1532_p_O_DFFX1));
  p_O_DFFX1 desc1533(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_opa_i[27:27]),.E(p_desc1533_p_O_DFFX1));
  p_O_DFFX1 desc1534(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_opa_i[26:26]),.E(p_desc1534_p_O_DFFX1));
  p_O_DFFX1 desc1535(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_opa_i[25:25]),.E(p_desc1535_p_O_DFFX1));
  p_O_DFFX1 desc1536(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_opa_i[24:24]),.E(p_desc1536_p_O_DFFX1));
  p_O_DFFX1 desc1537(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_opa_i[23:23]),.E(p_desc1537_p_O_DFFX1));
  p_O_DFFX1 desc1538(.D(opa_i[22:22]),.CLK(clk_i),.Q(s_opa_i[22:22]),.E(p_desc1538_p_O_DFFX1));
  p_O_DFFX1 desc1539(.D(opa_i[21:21]),.CLK(clk_i),.Q(s_opa_i[21:21]),.E(p_desc1539_p_O_DFFX1));
  p_O_DFFX1 desc1540(.D(opa_i[20:20]),.CLK(clk_i),.Q(s_opa_i[20:20]),.E(p_desc1540_p_O_DFFX1));
  p_O_DFFX1 desc1541(.D(opa_i[19:19]),.CLK(clk_i),.Q(s_opa_i[19:19]),.E(p_desc1541_p_O_DFFX1));
  p_O_DFFX1 desc1542(.D(opa_i[18:18]),.CLK(clk_i),.Q(s_opa_i[18:18]),.E(p_desc1542_p_O_DFFX1));
  p_O_DFFX1 desc1543(.D(opa_i[17:17]),.CLK(clk_i),.Q(s_opa_i[17:17]),.E(p_desc1543_p_O_DFFX1));
  p_O_DFFX1 desc1544(.D(opa_i[16:16]),.CLK(clk_i),.Q(s_opa_i[16:16]),.E(p_desc1544_p_O_DFFX1));
  p_O_DFFX1 desc1545(.D(opa_i[15:15]),.CLK(clk_i),.Q(s_opa_i[15:15]),.E(p_desc1545_p_O_DFFX1));
  p_O_DFFX1 desc1546(.D(opa_i[14:14]),.CLK(clk_i),.Q(s_opa_i[14:14]),.E(p_desc1546_p_O_DFFX1));
  p_O_DFFX1 desc1547(.D(opa_i[13:13]),.CLK(clk_i),.Q(s_opa_i[13:13]),.E(p_desc1547_p_O_DFFX1));
  p_O_DFFX1 desc1548(.D(opa_i[12:12]),.CLK(clk_i),.Q(s_opa_i[12:12]),.E(p_desc1548_p_O_DFFX1));
  p_O_DFFX1 desc1549(.D(opa_i[11:11]),.CLK(clk_i),.Q(s_opa_i[11:11]),.E(p_desc1549_p_O_DFFX1));
  p_O_DFFX1 desc1550(.D(opa_i[10:10]),.CLK(clk_i),.Q(s_opa_i[10:10]),.E(p_desc1550_p_O_DFFX1));
  p_O_DFFX1 desc1551(.D(opa_i[9:9]),.CLK(clk_i),.Q(s_opa_i[9:9]),.E(p_desc1551_p_O_DFFX1));
  p_O_DFFX1 desc1552(.D(opa_i[8:8]),.CLK(clk_i),.Q(s_opa_i[8:8]),.E(p_desc1552_p_O_DFFX1));
  p_O_DFFX1 desc1553(.D(opa_i[7:7]),.CLK(clk_i),.Q(s_opa_i[7:7]),.E(p_desc1553_p_O_DFFX1));
  p_O_DFFX1 desc1554(.D(opa_i[6:6]),.CLK(clk_i),.Q(s_opa_i[6:6]),.E(p_desc1554_p_O_DFFX1));
  p_O_DFFX1 desc1555(.D(opa_i[5:5]),.CLK(clk_i),.Q(s_opa_i[5:5]),.E(p_desc1555_p_O_DFFX1));
  p_O_DFFX1 desc1556(.D(opa_i[4:4]),.CLK(clk_i),.Q(s_opa_i[4:4]),.E(p_desc1556_p_O_DFFX1));
  p_O_DFFX1 desc1557(.D(opa_i[3:3]),.CLK(clk_i),.Q(s_opa_i[3:3]),.E(p_desc1557_p_O_DFFX1));
  p_O_DFFX1 desc1558(.D(opa_i[2:2]),.CLK(clk_i),.Q(s_opa_i[2:2]),.E(p_desc1558_p_O_DFFX1));
  p_O_DFFX1 desc1559(.D(opa_i[1:1]),.CLK(clk_i),.Q(s_opa_i[1:1]),.E(p_desc1559_p_O_DFFX1));
  p_O_DFFX1 desc1560(.D(opa_i[0:0]),.CLK(clk_i),.Q(s_opa_i[0:0]),.E(p_desc1560_p_O_DFFX1));
  p_O_DFFX1 desc1561(.D(opb_i[30:30]),.CLK(clk_i),.Q(s_opb_i[30:30]),.E(p_desc1561_p_O_DFFX1));
  p_O_DFFX1 desc1562(.D(opb_i[29:29]),.CLK(clk_i),.Q(s_opb_i[29:29]),.E(p_desc1562_p_O_DFFX1));
  p_O_DFFX1 desc1563(.D(opb_i[28:28]),.CLK(clk_i),.Q(s_opb_i[28:28]),.E(p_desc1563_p_O_DFFX1));
  p_O_DFFX1 desc1564(.D(opb_i[27:27]),.CLK(clk_i),.Q(s_opb_i[27:27]),.E(p_desc1564_p_O_DFFX1));
  p_O_DFFX1 desc1565(.D(opb_i[26:26]),.CLK(clk_i),.Q(s_opb_i[26:26]),.E(p_desc1565_p_O_DFFX1));
  p_O_DFFX1 desc1566(.D(opb_i[25:25]),.CLK(clk_i),.Q(s_opb_i[25:25]),.E(p_desc1566_p_O_DFFX1));
  p_O_DFFX1 desc1567(.D(opb_i[24:24]),.CLK(clk_i),.Q(s_opb_i[24:24]),.E(p_desc1567_p_O_DFFX1));
  p_O_DFFX1 desc1568(.D(opb_i[23:23]),.CLK(clk_i),.Q(s_opb_i[23:23]),.E(p_desc1568_p_O_DFFX1));
  p_O_DFFX1 desc1569(.D(opb_i[22:22]),.CLK(clk_i),.Q(s_opb_i[22:22]),.E(p_desc1569_p_O_DFFX1));
  p_O_DFFX1 desc1570(.D(opb_i[21:21]),.CLK(clk_i),.Q(s_opb_i[21:21]),.E(p_desc1570_p_O_DFFX1));
  p_O_DFFX1 desc1571(.D(opb_i[20:20]),.CLK(clk_i),.Q(s_opb_i[20:20]),.E(p_desc1571_p_O_DFFX1));
  p_O_DFFX1 desc1572(.D(opb_i[19:19]),.CLK(clk_i),.Q(s_opb_i[19:19]),.E(p_desc1572_p_O_DFFX1));
  p_O_DFFX1 desc1573(.D(opb_i[18:18]),.CLK(clk_i),.Q(s_opb_i[18:18]),.E(p_desc1573_p_O_DFFX1));
  p_O_DFFX1 desc1574(.D(opb_i[17:17]),.CLK(clk_i),.Q(s_opb_i[17:17]),.E(p_desc1574_p_O_DFFX1));
  p_O_DFFX1 desc1575(.D(opb_i[16:16]),.CLK(clk_i),.Q(s_opb_i[16:16]),.E(p_desc1575_p_O_DFFX1));
  p_O_DFFX1 desc1576(.D(opb_i[15:15]),.CLK(clk_i),.Q(s_opb_i[15:15]),.E(p_desc1576_p_O_DFFX1));
  p_O_DFFX1 desc1577(.D(opb_i[14:14]),.CLK(clk_i),.Q(s_opb_i[14:14]),.E(p_desc1577_p_O_DFFX1));
  p_O_DFFX1 desc1578(.D(opb_i[13:13]),.CLK(clk_i),.Q(s_opb_i[13:13]),.E(p_desc1578_p_O_DFFX1));
  p_O_DFFX1 desc1579(.D(opb_i[12:12]),.CLK(clk_i),.Q(s_opb_i[12:12]),.E(p_desc1579_p_O_DFFX1));
  p_O_DFFX1 desc1580(.D(opb_i[11:11]),.CLK(clk_i),.Q(s_opb_i[11:11]),.E(p_desc1580_p_O_DFFX1));
  p_O_DFFX1 desc1581(.D(opb_i[10:10]),.CLK(clk_i),.Q(s_opb_i[10:10]),.E(p_desc1581_p_O_DFFX1));
  p_O_DFFX1 desc1582(.D(opb_i[9:9]),.CLK(clk_i),.Q(s_opb_i[9:9]),.E(p_desc1582_p_O_DFFX1));
  p_O_DFFX1 desc1583(.D(opb_i[8:8]),.CLK(clk_i),.Q(s_opb_i[8:8]),.E(p_desc1583_p_O_DFFX1));
  p_O_DFFX1 desc1584(.D(opb_i[7:7]),.CLK(clk_i),.Q(s_opb_i[7:7]),.E(p_desc1584_p_O_DFFX1));
  p_O_DFFX1 desc1585(.D(opb_i[6:6]),.CLK(clk_i),.Q(s_opb_i[6:6]),.E(p_desc1585_p_O_DFFX1));
  p_O_DFFX1 desc1586(.D(opb_i[5:5]),.CLK(clk_i),.Q(s_opb_i[5:5]),.E(p_desc1586_p_O_DFFX1));
  p_O_DFFX1 desc1587(.D(opb_i[4:4]),.CLK(clk_i),.Q(s_opb_i[4:4]),.E(p_desc1587_p_O_DFFX1));
  p_O_DFFX1 desc1588(.D(opb_i[3:3]),.CLK(clk_i),.Q(s_opb_i[3:3]),.E(p_desc1588_p_O_DFFX1));
  p_O_DFFX1 desc1589(.D(opb_i[2:2]),.CLK(clk_i),.Q(s_opb_i[2:2]),.E(p_desc1589_p_O_DFFX1));
  p_O_DFFX1 desc1590(.D(opb_i[1:1]),.CLK(clk_i),.Q(s_opb_i[1:1]),.E(p_desc1590_p_O_DFFX1));
  p_O_DFFX1 desc1591(.D(opb_i[0:0]),.CLK(clk_i),.Q(s_opb_i[0:0]),.E(p_desc1591_p_O_DFFX1));
  p_O_DFFX1 desc1592(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_expa[7:7]),.E(p_desc1592_p_O_DFFX1));
  p_O_DFFX1 desc1593(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_expa[6:6]),.E(p_desc1593_p_O_DFFX1));
  p_O_DFFX1 desc1594(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_expa[5:5]),.E(p_desc1594_p_O_DFFX1));
  p_O_DFFX1 desc1595(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_expa[4:4]),.E(p_desc1595_p_O_DFFX1));
  p_O_DFFX1 desc1596(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_expa[3:3]),.E(p_desc1596_p_O_DFFX1));
  p_O_DFFX1 desc1597(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_expa[2:2]),.E(p_desc1597_p_O_DFFX1));
  p_O_DFFX1 desc1598(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_expa[1:1]),.E(p_desc1598_p_O_DFFX1));
  p_O_DFFX1 desc1599(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_expa[0:0]),.E(p_desc1599_p_O_DFFX1));
  p_O_DFFX1 desc1600(.D(opb_i[30:30]),.CLK(clk_i),.Q(s_expb[7:7]),.E(p_desc1600_p_O_DFFX1));
  p_O_DFFX1 desc1601(.D(opb_i[29:29]),.CLK(clk_i),.Q(s_expb[6:6]),.E(p_desc1601_p_O_DFFX1));
  p_O_DFFX1 desc1602(.D(opb_i[28:28]),.CLK(clk_i),.Q(s_expb[5:5]),.E(p_desc1602_p_O_DFFX1));
  p_O_DFFX1 desc1603(.D(opb_i[27:27]),.CLK(clk_i),.Q(s_expb[4:4]),.E(p_desc1603_p_O_DFFX1));
  p_O_DFFX1 desc1604(.D(opb_i[26:26]),.CLK(clk_i),.Q(s_expb[3:3]),.E(p_desc1604_p_O_DFFX1));
  p_O_DFFX1 desc1605(.D(opb_i[25:25]),.CLK(clk_i),.Q(s_expb[2:2]),.E(p_desc1605_p_O_DFFX1));
  p_O_DFFX1 desc1606(.D(opb_i[24:24]),.CLK(clk_i),.Q(s_expb[1:1]),.E(p_desc1606_p_O_DFFX1));
  p_O_DFFX1 desc1607(.D(opb_i[23:23]),.CLK(clk_i),.Q(s_expb[0:0]),.E(p_desc1607_p_O_DFFX1));
  p_O_DFFX1 desc1608(.D(qutnt_i[26:26]),.CLK(clk_i),.Q(s_qutnt_i[26:26]),.QN(\sub_1_root_sub_150_2/CI ),.E(p_desc1608_p_O_DFFX1));
  p_O_DFFX1 desc1609(.D(qutnt_i[5:5]),.CLK(clk_i),.Q(s_qutnt_i[5:5]),.QN(n106),.E(p_desc1609_p_O_DFFX1));
  p_O_DFFX1 desc1610(.D(qutnt_i[4:4]),.CLK(clk_i),.Q(s_qutnt_i[4:4]),.QN(n108),.E(p_desc1610_p_O_DFFX1));
  p_O_DFFX1 desc1611(.D(qutnt_i[3:3]),.CLK(clk_i),.Q(s_qutnt_i[3:3]),.E(p_desc1611_p_O_DFFX1));
  p_O_DFFX1 desc1612(.D(qutnt_i[2:2]),.CLK(clk_i),.Q(s_qutnt_i[2:2]),.QN(n112),.E(p_desc1612_p_O_DFFX1));
  p_O_DFFX1 desc1613(.D(qutnt_i[1:1]),.CLK(clk_i),.Q(s_qutnt_i[1:1]),.E(p_desc1613_p_O_DFFX1));
  p_O_DFFX1 desc1614(.D(qutnt_i[0:0]),.CLK(clk_i),.Q(s_qutnt_i[0:0]),.QN(n113),.E(p_desc1614_p_O_DFFX1));
  p_O_DFFX1 desc1615(.D(rmndr_i[26:26]),.CLK(clk_i),.Q(s_rmndr_i[26:26]),.E(p_desc1615_p_O_DFFX1));
  p_O_DFFX1 desc1616(.D(rmndr_i[25:25]),.CLK(clk_i),.Q(s_rmndr_i[25:25]),.E(p_desc1616_p_O_DFFX1));
  p_O_DFFX1 desc1617(.D(rmndr_i[24:24]),.CLK(clk_i),.Q(s_rmndr_i[24:24]),.E(p_desc1617_p_O_DFFX1));
  p_O_DFFX1 desc1618(.D(rmndr_i[23:23]),.CLK(clk_i),.Q(s_rmndr_i[23:23]),.E(p_desc1618_p_O_DFFX1));
  p_O_DFFX1 desc1619(.D(rmndr_i[22:22]),.CLK(clk_i),.Q(s_rmndr_i[22:22]),.E(p_desc1619_p_O_DFFX1));
  p_O_DFFX1 desc1620(.D(rmndr_i[21:21]),.CLK(clk_i),.Q(s_rmndr_i[21:21]),.E(p_desc1620_p_O_DFFX1));
  p_O_DFFX1 desc1621(.D(rmndr_i[20:20]),.CLK(clk_i),.Q(s_rmndr_i[20:20]),.E(p_desc1621_p_O_DFFX1));
  p_O_DFFX1 desc1622(.D(rmndr_i[19:19]),.CLK(clk_i),.Q(s_rmndr_i[19:19]),.E(p_desc1622_p_O_DFFX1));
  p_O_DFFX1 desc1623(.D(rmndr_i[18:18]),.CLK(clk_i),.Q(s_rmndr_i[18:18]),.E(p_desc1623_p_O_DFFX1));
  p_O_DFFX1 desc1624(.D(rmndr_i[17:17]),.CLK(clk_i),.Q(s_rmndr_i[17:17]),.E(p_desc1624_p_O_DFFX1));
  p_O_DFFX1 desc1625(.D(rmndr_i[16:16]),.CLK(clk_i),.Q(s_rmndr_i[16:16]),.E(p_desc1625_p_O_DFFX1));
  p_O_DFFX1 desc1626(.D(rmndr_i[15:15]),.CLK(clk_i),.Q(s_rmndr_i[15:15]),.E(p_desc1626_p_O_DFFX1));
  p_O_DFFX1 desc1627(.D(rmndr_i[14:14]),.CLK(clk_i),.Q(s_rmndr_i[14:14]),.E(p_desc1627_p_O_DFFX1));
  p_O_DFFX1 desc1628(.D(rmndr_i[13:13]),.CLK(clk_i),.Q(s_rmndr_i[13:13]),.E(p_desc1628_p_O_DFFX1));
  p_O_DFFX1 desc1629(.D(rmndr_i[12:12]),.CLK(clk_i),.Q(s_rmndr_i[12:12]),.E(p_desc1629_p_O_DFFX1));
  p_O_DFFX1 desc1630(.D(rmndr_i[11:11]),.CLK(clk_i),.Q(s_rmndr_i[11:11]),.E(p_desc1630_p_O_DFFX1));
  p_O_DFFX1 desc1631(.D(rmndr_i[10:10]),.CLK(clk_i),.Q(s_rmndr_i[10:10]),.E(p_desc1631_p_O_DFFX1));
  p_O_DFFX1 desc1632(.D(rmndr_i[9:9]),.CLK(clk_i),.Q(s_rmndr_i[9:9]),.E(p_desc1632_p_O_DFFX1));
  p_O_DFFX1 desc1633(.D(rmndr_i[8:8]),.CLK(clk_i),.Q(s_rmndr_i[8:8]),.E(p_desc1633_p_O_DFFX1));
  p_O_DFFX1 desc1634(.D(rmndr_i[7:7]),.CLK(clk_i),.Q(s_rmndr_i[7:7]),.E(p_desc1634_p_O_DFFX1));
  p_O_DFFX1 desc1635(.D(rmndr_i[6:6]),.CLK(clk_i),.Q(s_rmndr_i[6:6]),.E(p_desc1635_p_O_DFFX1));
  p_O_DFFX1 desc1636(.D(rmndr_i[5:5]),.CLK(clk_i),.Q(s_rmndr_i[5:5]),.E(p_desc1636_p_O_DFFX1));
  p_O_DFFX1 desc1637(.D(rmndr_i[4:4]),.CLK(clk_i),.Q(s_rmndr_i[4:4]),.E(p_desc1637_p_O_DFFX1));
  p_O_DFFX1 desc1638(.D(rmndr_i[3:3]),.CLK(clk_i),.Q(s_rmndr_i[3:3]),.E(p_desc1638_p_O_DFFX1));
  p_O_DFFX1 desc1639(.D(rmndr_i[2:2]),.CLK(clk_i),.Q(s_rmndr_i[2:2]),.E(p_desc1639_p_O_DFFX1));
  p_O_DFFX1 desc1640(.D(rmndr_i[1:1]),.CLK(clk_i),.Q(s_rmndr_i[1:1]),.E(p_desc1640_p_O_DFFX1));
  p_O_DFFX1 desc1641(.D(rmndr_i[0:0]),.CLK(clk_i),.Q(s_rmndr_i[0:0]),.E(p_desc1641_p_O_DFFX1));
  p_O_DFFX1 desc1642(.D(exp_10_i[9:9]),.CLK(clk_i),.Q(s_exp_10_i[9:9]),.E(p_desc1642_p_O_DFFX1));
  p_O_DFFX1 desc1643(.D(exp_10_i[8:8]),.CLK(clk_i),.Q(s_exp_10_i[8:8]),.E(p_desc1643_p_O_DFFX1));
  p_O_DFFX1 desc1644(.D(exp_10_i[7:7]),.CLK(clk_i),.Q(s_exp_10_i[7:7]),.E(p_desc1644_p_O_DFFX1));
  p_O_DFFX1 desc1645(.D(exp_10_i[6:6]),.CLK(clk_i),.Q(s_exp_10_i[6:6]),.E(p_desc1645_p_O_DFFX1));
  p_O_DFFX1 desc1646(.D(exp_10_i[5:5]),.CLK(clk_i),.Q(s_exp_10_i[5:5]),.E(p_desc1646_p_O_DFFX1));
  p_O_DFFX1 desc1647(.D(exp_10_i[4:4]),.CLK(clk_i),.Q(s_exp_10_i[4:4]),.E(p_desc1647_p_O_DFFX1));
  p_O_DFFX1 desc1648(.D(exp_10_i[3:3]),.CLK(clk_i),.Q(s_exp_10_i[3:3]),.E(p_desc1648_p_O_DFFX1));
  p_O_DFFX1 desc1649(.D(exp_10_i[2:2]),.CLK(clk_i),.Q(s_exp_10_i[2:2]),.E(p_desc1649_p_O_DFFX1));
  p_O_DFFX1 desc1650(.D(exp_10_i[1:1]),.CLK(clk_i),.Q(s_exp_10_i[1:1]),.E(p_desc1650_p_O_DFFX1));
  p_O_DFFX1 desc1651(.D(exp_10_i[0:0]),.CLK(clk_i),.Q(s_exp_10_i[0:0]),.E(p_desc1651_p_O_DFFX1));
  p_O_DFFX1 s_sign_i_reg(.D(sign_i),.CLK(clk_i),.Q(s_sign_i),.QN(n117),.E(p_s_sign_i_reg_p_O_DFFX1));
  p_O_DFFX1 desc1652(.D(rmode_i[1:1]),.CLK(clk_i),.Q(\s_rmode_i[1] ),.QN(n118),.E(p_desc1652_p_O_DFFX1));
  p_O_DFFX1 desc1653(.D(rmode_i[0:0]),.CLK(clk_i),.QN(n119),.E(p_desc1653_p_O_DFFX1));
  p_O_DFFX1 desc1654(.D(s_output_o[31:31]),.CLK(clk_i),.Q(output_o[31:31]),.E(p_desc1654_p_O_DFFX1));
  DFFSSRX1 desc1655(.D(n264),.RSTB(s_exp_10b[8:8]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[8:8]));
  DFFSSRX1 desc1656(.D(n264),.RSTB(s_exp_10b[7:7]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[7:7]));
  DFFSSRX1 desc1657(.D(n264),.RSTB(s_exp_10b[6:6]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[6:6]));
  p_O_DFFX1 desc1658(.D(N167),.CLK(clk_i),.Q(s_expo1[5:5]),.E(p_desc1658_p_O_DFFX1));
  p_O_DFFX1 desc1659(.D(N166),.CLK(clk_i),.Q(s_expo1[4:4]),.E(p_desc1659_p_O_DFFX1));
  DFFSSRX1 desc1660(.D(n264),.RSTB(s_exp_10b[3:3]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[3:3]));
  DFFSSRX1 desc1661(.D(n264),.RSTB(s_exp_10b[2:2]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[2:2]));
  DFFSSRX1 desc1662(.D(n264),.RSTB(s_exp_10b[1:1]),.SETB(1'b1),.CLK(clk_i),.Q(s_expo1[1:1]));
  p_O_DFFX1 desc1663(.D(N162),.CLK(clk_i),.Q(s_expo1[0:0]),.E(p_desc1663_p_O_DFFX1));
  p_O_DFFX1 desc1664(.D(N177),.CLK(clk_i),.Q(s_shr1[5:5]),.E(p_desc1664_p_O_DFFX1));
  p_O_DFFX1 desc1665(.D(N176),.CLK(clk_i),.Q(s_shr1[4:4]),.E(p_desc1665_p_O_DFFX1));
  p_O_DFFX1 desc1666(.D(N174),.CLK(clk_i),.Q(s_shr1[2:2]),.QN(n2),.E(p_desc1666_p_O_DFFX1));
  p_O_DFFX1 desc1667(.D(N173),.CLK(clk_i),.Q(s_shr1[1:1]),.QN(n5),.E(p_desc1667_p_O_DFFX1));
  p_O_DFFX1 desc1668(.D(N172),.CLK(clk_i),.Q(s_shr1[0:0]),.QN(n6),.E(p_desc1668_p_O_DFFX1));
  p_O_DFFX1 desc1669(.D(N161),.CLK(clk_i),.Q(\s_shl1[0] ),.E(p_desc1669_p_O_DFFX1));
  p_O_DFFX1 desc1670(.D(N264),.CLK(clk_i),.Q(s_fraco1[26:26]),.E(p_desc1670_p_O_DFFX1));
  p_O_DFFX1 desc1671(.D(N263),.CLK(clk_i),.Q(s_fraco1[25:25]),.E(p_desc1671_p_O_DFFX1));
  p_O_DFFX1 desc1672(.D(N262),.CLK(clk_i),.Q(s_fraco1[24:24]),.E(p_desc1672_p_O_DFFX1));
  p_O_DFFX1 desc1673(.D(N261),.CLK(clk_i),.Q(s_fraco1[23:23]),.E(p_desc1673_p_O_DFFX1));
  p_O_DFFX1 desc1674(.D(N260),.CLK(clk_i),.Q(s_fraco1[22:22]),.E(p_desc1674_p_O_DFFX1));
  p_O_DFFX1 desc1675(.D(N259),.CLK(clk_i),.Q(s_fraco1[21:21]),.E(p_desc1675_p_O_DFFX1));
  p_O_DFFX1 desc1676(.D(N258),.CLK(clk_i),.Q(s_fraco1[20:20]),.E(p_desc1676_p_O_DFFX1));
  p_O_DFFX1 desc1677(.D(N257),.CLK(clk_i),.Q(s_fraco1[19:19]),.E(p_desc1677_p_O_DFFX1));
  p_O_DFFX1 desc1678(.D(N256),.CLK(clk_i),.Q(s_fraco1[18:18]),.E(p_desc1678_p_O_DFFX1));
  p_O_DFFX1 desc1679(.D(N255),.CLK(clk_i),.Q(s_fraco1[17:17]),.E(p_desc1679_p_O_DFFX1));
  p_O_DFFX1 desc1680(.D(N254),.CLK(clk_i),.Q(s_fraco1[16:16]),.E(p_desc1680_p_O_DFFX1));
  p_O_DFFX1 desc1681(.D(N253),.CLK(clk_i),.Q(s_fraco1[15:15]),.E(p_desc1681_p_O_DFFX1));
  p_O_DFFX1 desc1682(.D(N252),.CLK(clk_i),.Q(s_fraco1[14:14]),.E(p_desc1682_p_O_DFFX1));
  p_O_DFFX1 desc1683(.D(N251),.CLK(clk_i),.Q(s_fraco1[13:13]),.E(p_desc1683_p_O_DFFX1));
  p_O_DFFX1 desc1684(.D(N250),.CLK(clk_i),.Q(s_fraco1[12:12]),.E(p_desc1684_p_O_DFFX1));
  p_O_DFFX1 desc1685(.D(N249),.CLK(clk_i),.Q(s_fraco1[11:11]),.E(p_desc1685_p_O_DFFX1));
  p_O_DFFX1 desc1686(.D(N248),.CLK(clk_i),.Q(s_fraco1[10:10]),.E(p_desc1686_p_O_DFFX1));
  p_O_DFFX1 desc1687(.D(N247),.CLK(clk_i),.Q(s_fraco1[9:9]),.E(p_desc1687_p_O_DFFX1));
  p_O_DFFX1 desc1688(.D(N246),.CLK(clk_i),.Q(s_fraco1[8:8]),.E(p_desc1688_p_O_DFFX1));
  p_O_DFFX1 desc1689(.D(N245),.CLK(clk_i),.Q(s_fraco1[7:7]),.E(p_desc1689_p_O_DFFX1));
  p_O_DFFX1 desc1690(.D(N244),.CLK(clk_i),.Q(s_fraco1[6:6]),.E(p_desc1690_p_O_DFFX1));
  p_O_DFFX1 desc1691(.D(N243),.CLK(clk_i),.Q(s_fraco1[5:5]),.E(p_desc1691_p_O_DFFX1));
  p_O_DFFX1 desc1692(.D(N242),.CLK(clk_i),.Q(s_fraco1[4:4]),.E(p_desc1692_p_O_DFFX1));
  p_O_DFFX1 desc1693(.D(N241),.CLK(clk_i),.Q(s_fraco1[3:3]),.QN(n122),.E(p_desc1693_p_O_DFFX1));
  p_O_DFFX1 desc1694(.D(N240),.CLK(clk_i),.Q(s_fraco1[2:2]),.QN(n123),.E(p_desc1694_p_O_DFFX1));
  p_O_DFFX1 desc1695(.D(N239),.CLK(clk_i),.QN(n124),.E(p_desc1695_p_O_DFFX1));
  p_O_DFFX1 desc1696(.D(N238),.CLK(clk_i),.Q(s_fraco1[0:0]),.E(p_desc1696_p_O_DFFX1));
  p_O_DFFX1 desc1697(.D(N1131),.CLK(clk_i),.Q(s_fraco2[22:22]),.E(p_desc1697_p_O_DFFX1));
  p_O_DFFX1 desc1698(.D(N1130),.CLK(clk_i),.Q(s_fraco2[21:21]),.E(p_desc1698_p_O_DFFX1));
  p_O_DFFX1 desc1699(.D(N1129),.CLK(clk_i),.Q(s_fraco2[20:20]),.E(p_desc1699_p_O_DFFX1));
  p_O_DFFX1 desc1700(.D(N1128),.CLK(clk_i),.Q(s_fraco2[19:19]),.E(p_desc1700_p_O_DFFX1));
  p_O_DFFX1 desc1701(.D(N1127),.CLK(clk_i),.Q(s_fraco2[18:18]),.E(p_desc1701_p_O_DFFX1));
  p_O_DFFX1 desc1702(.D(N1126),.CLK(clk_i),.Q(s_fraco2[17:17]),.E(p_desc1702_p_O_DFFX1));
  p_O_DFFX1 desc1703(.D(N1125),.CLK(clk_i),.Q(s_fraco2[16:16]),.E(p_desc1703_p_O_DFFX1));
  p_O_DFFX1 desc1704(.D(N1124),.CLK(clk_i),.Q(s_fraco2[15:15]),.E(p_desc1704_p_O_DFFX1));
  p_O_DFFX1 desc1705(.D(N1123),.CLK(clk_i),.Q(s_fraco2[14:14]),.E(p_desc1705_p_O_DFFX1));
  p_O_DFFX1 desc1706(.D(N1122),.CLK(clk_i),.Q(s_fraco2[13:13]),.E(p_desc1706_p_O_DFFX1));
  p_O_DFFX1 desc1707(.D(N1121),.CLK(clk_i),.Q(s_fraco2[12:12]),.E(p_desc1707_p_O_DFFX1));
  p_O_DFFX1 desc1708(.D(N1120),.CLK(clk_i),.Q(s_fraco2[11:11]),.E(p_desc1708_p_O_DFFX1));
  p_O_DFFX1 desc1709(.D(N1119),.CLK(clk_i),.Q(s_fraco2[10:10]),.E(p_desc1709_p_O_DFFX1));
  p_O_DFFX1 desc1710(.D(N1118),.CLK(clk_i),.Q(s_fraco2[9:9]),.E(p_desc1710_p_O_DFFX1));
  p_O_DFFX1 desc1711(.D(N1117),.CLK(clk_i),.Q(s_fraco2[8:8]),.E(p_desc1711_p_O_DFFX1));
  p_O_DFFX1 desc1712(.D(N1116),.CLK(clk_i),.Q(s_fraco2[7:7]),.E(p_desc1712_p_O_DFFX1));
  p_O_DFFX1 desc1713(.D(N1115),.CLK(clk_i),.Q(s_fraco2[6:6]),.E(p_desc1713_p_O_DFFX1));
  p_O_DFFX1 desc1714(.D(N1114),.CLK(clk_i),.Q(s_fraco2[5:5]),.E(p_desc1714_p_O_DFFX1));
  p_O_DFFX1 desc1715(.D(N1113),.CLK(clk_i),.Q(s_fraco2[4:4]),.E(p_desc1715_p_O_DFFX1));
  p_O_DFFX1 desc1716(.D(N1112),.CLK(clk_i),.Q(s_fraco2[3:3]),.E(p_desc1716_p_O_DFFX1));
  p_O_DFFX1 desc1717(.D(N1111),.CLK(clk_i),.Q(s_fraco2[2:2]),.E(p_desc1717_p_O_DFFX1));
  p_O_DFFX1 desc1718(.D(N1110),.CLK(clk_i),.Q(s_fraco2[1:1]),.E(p_desc1718_p_O_DFFX1));
  p_O_DFFX1 desc1719(.D(N1109),.CLK(clk_i),.Q(s_fraco2[0:0]),.E(p_desc1719_p_O_DFFX1));
  p_O_DFFX1 desc1720(.D(N1108),.CLK(clk_i),.Q(s_expo3[8:8]),.E(p_desc1720_p_O_DFFX1));
  p_O_DFFX1 desc1721(.D(N1107),.CLK(clk_i),.Q(s_expo3[7:7]),.E(p_desc1721_p_O_DFFX1));
  p_O_DFFX1 desc1722(.D(N1106),.CLK(clk_i),.Q(s_expo3[6:6]),.E(p_desc1722_p_O_DFFX1));
  p_O_DFFX1 desc1723(.D(N1105),.CLK(clk_i),.Q(s_expo3[5:5]),.E(p_desc1723_p_O_DFFX1));
  p_O_DFFX1 desc1724(.D(N1104),.CLK(clk_i),.Q(s_expo3[4:4]),.E(p_desc1724_p_O_DFFX1));
  p_O_DFFX1 desc1725(.D(N1103),.CLK(clk_i),.Q(s_expo3[3:3]),.E(p_desc1725_p_O_DFFX1));
  p_O_DFFX1 desc1726(.D(N1102),.CLK(clk_i),.Q(s_expo3[2:2]),.E(p_desc1726_p_O_DFFX1));
  p_O_DFFX1 desc1727(.D(N1101),.CLK(clk_i),.Q(s_expo3[1:1]),.E(p_desc1727_p_O_DFFX1));
  p_O_DFFX1 desc1728(.D(N1100),.CLK(clk_i),.Q(s_expo3[0:0]),.E(p_desc1728_p_O_DFFX1));
  p_O_DFFX1 ine_o_reg(.D(N1386),.CLK(clk_i),.Q(ine_o),.E(p_ine_o_reg_p_O_DFFX1));
  p_O_DFFX1 desc1729(.D(s_output_o[22:22]),.CLK(clk_i),.Q(output_o[22:22]),.E(p_desc1729_p_O_DFFX1));
  DFFSSRX1 desc1730(.D(n247),.RSTB(s_expo3[1:1]),.SETB(n249),.CLK(clk_i),.Q(output_o[24:24]));
  DFFSSRX1 desc1731(.D(n247),.RSTB(s_expo3[2:2]),.SETB(n249),.CLK(clk_i),.Q(output_o[25:25]));
  DFFSSRX1 desc1732(.D(n247),.RSTB(s_expo3[3:3]),.SETB(n249),.CLK(clk_i),.Q(output_o[26:26]));
  DFFSSRX1 desc1733(.D(n247),.RSTB(s_expo3[4:4]),.SETB(n249),.CLK(clk_i),.Q(output_o[27:27]));
  DFFSSRX1 desc1734(.D(n247),.RSTB(s_expo3[5:5]),.SETB(n249),.CLK(clk_i),.Q(output_o[28:28]));
  DFFSSRX1 desc1735(.D(n247),.RSTB(s_expo3[6:6]),.SETB(n249),.CLK(clk_i),.Q(output_o[29:29]));
  DFFSSRX1 desc1736(.D(n247),.RSTB(s_expo3[7:7]),.SETB(n249),.CLK(clk_i),.Q(output_o[30:30]));
  p_O_DFFX1 desc1737(.D(s_output_o[9:9]),.CLK(clk_i),.Q(output_o[9:9]),.E(p_desc1737_p_O_DFFX1));
  p_O_DFFX1 desc1738(.D(s_output_o[8:8]),.CLK(clk_i),.Q(output_o[8:8]),.E(p_desc1738_p_O_DFFX1));
  p_O_DFFX1 desc1739(.D(s_output_o[7:7]),.CLK(clk_i),.Q(output_o[7:7]),.E(p_desc1739_p_O_DFFX1));
  p_O_DFFX1 desc1740(.D(s_output_o[6:6]),.CLK(clk_i),.Q(output_o[6:6]),.E(p_desc1740_p_O_DFFX1));
  p_O_DFFX1 desc1741(.D(s_output_o[5:5]),.CLK(clk_i),.Q(output_o[5:5]),.E(p_desc1741_p_O_DFFX1));
  p_O_DFFX1 desc1742(.D(s_output_o[4:4]),.CLK(clk_i),.Q(output_o[4:4]),.E(p_desc1742_p_O_DFFX1));
  p_O_DFFX1 desc1743(.D(s_output_o[3:3]),.CLK(clk_i),.Q(output_o[3:3]),.E(p_desc1743_p_O_DFFX1));
  p_O_DFFX1 desc1744(.D(s_output_o[2:2]),.CLK(clk_i),.Q(output_o[2:2]),.E(p_desc1744_p_O_DFFX1));
  p_O_DFFX1 desc1745(.D(s_output_o[21:21]),.CLK(clk_i),.Q(output_o[21:21]),.E(p_desc1745_p_O_DFFX1));
  p_O_DFFX1 desc1746(.D(s_output_o[20:20]),.CLK(clk_i),.Q(output_o[20:20]),.E(p_desc1746_p_O_DFFX1));
  p_O_DFFX1 desc1747(.D(s_output_o[1:1]),.CLK(clk_i),.Q(output_o[1:1]),.E(p_desc1747_p_O_DFFX1));
  p_O_DFFX1 desc1748(.D(s_output_o[19:19]),.CLK(clk_i),.Q(output_o[19:19]),.E(p_desc1748_p_O_DFFX1));
  p_O_DFFX1 desc1749(.D(s_output_o[18:18]),.CLK(clk_i),.Q(output_o[18:18]),.E(p_desc1749_p_O_DFFX1));
  p_O_DFFX1 desc1750(.D(s_output_o[17:17]),.CLK(clk_i),.Q(output_o[17:17]),.E(p_desc1750_p_O_DFFX1));
  p_O_DFFX1 desc1751(.D(s_output_o[16:16]),.CLK(clk_i),.Q(output_o[16:16]),.E(p_desc1751_p_O_DFFX1));
  p_O_DFFX1 desc1752(.D(s_output_o[15:15]),.CLK(clk_i),.Q(output_o[15:15]),.E(p_desc1752_p_O_DFFX1));
  p_O_DFFX1 desc1753(.D(s_output_o[14:14]),.CLK(clk_i),.Q(output_o[14:14]),.E(p_desc1753_p_O_DFFX1));
  p_O_DFFX1 desc1754(.D(s_output_o[13:13]),.CLK(clk_i),.Q(output_o[13:13]),.E(p_desc1754_p_O_DFFX1));
  p_O_DFFX1 desc1755(.D(s_output_o[12:12]),.CLK(clk_i),.Q(output_o[12:12]),.E(p_desc1755_p_O_DFFX1));
  p_O_DFFX1 desc1756(.D(s_output_o[11:11]),.CLK(clk_i),.Q(output_o[11:11]),.E(p_desc1756_p_O_DFFX1));
  p_O_DFFX1 desc1757(.D(s_output_o[10:10]),.CLK(clk_i),.Q(output_o[10:10]),.E(p_desc1757_p_O_DFFX1));
  p_O_DFFX1 desc1758(.D(s_output_o[0:0]),.CLK(clk_i),.Q(output_o[0:0]),.E(p_desc1758_p_O_DFFX1));
  DFFSSRX1 desc1759(.D(n247),.RSTB(s_expo3[0:0]),.SETB(n249),.CLK(clk_i),.Q(output_o[23:23]));
  AO22X1 U128(.IN1(n130),.IN2(N364),.IN3(n131),.IN4(n12),.Q(n129));
  NAND3X0 U129(.IN1(n132),.IN2(n133),.IN3(n134),.QN(n128));
  AOI222X1 U130(.IN1(n135),.IN2(N432),.IN3(n136),.IN4(N483),.IN5(n137),.IN6(n138),.QN(n134));
  NAND3X0 U131(.IN1(n139),.IN2(n140),.IN3(n141),.QN(n138));
  OA222X1 U132(.IN1(n66),.IN2(n142),.IN3(n58),.IN4(n143),.IN5(n144),.IN6(n145),.Q(n141));
  AO222X1 U133(.IN1(n148),.IN2(N619),.IN3(s_qutnt_i[21:21]),.IN4(N602),.IN5(n149),.IN6(N636),.Q(n147));
  AO222X1 U134(.IN1(N681),.IN2(n75),.IN3(n150),.IN4(N653),.IN5(n151),.IN6(N670),.Q(n146));
  AOI22X1 U135(.IN1(N500),.IN2(s_qutnt_i[15:15]),.IN3(N517),.IN4(n152),.QN(n140));
  OA22X1 U136(.IN1(n65),.IN2(n153),.IN3(n59),.IN4(n154),.Q(n139));
  AOI22X1 U137(.IN1(N398),.IN2(s_qutnt_i[9:9]),.IN3(N415),.IN4(n155),.QN(n133));
  AOI22X1 U138(.IN1(N449),.IN2(n156),.IN3(N466),.IN4(n157),.QN(n132));
  AO222X1 U140(.IN1(n130),.IN2(N363),.IN3(n131),.IN4(N346),.IN5(n126),.IN6(N380),.Q(n160));
  NAND3X0 U141(.IN1(n161),.IN2(n162),.IN3(n163),.QN(n158));
  AOI222X1 U142(.IN1(n135),.IN2(N431),.IN3(n136),.IN4(N482),.IN5(n137),.IN6(n164),.QN(n163));
  NAND3X0 U143(.IN1(n165),.IN2(n166),.IN3(n167),.QN(n164));
  OA222X1 U144(.IN1(n70),.IN2(n142),.IN3(n67),.IN4(n143),.IN5(n168),.IN6(n145),.Q(n167));
  AO222X1 U145(.IN1(n148),.IN2(N618),.IN3(s_qutnt_i[21:21]),.IN4(N601),.IN5(n149),.IN6(N635),.Q(n170));
  AO222X1 U146(.IN1(N680),.IN2(n75),.IN3(n150),.IN4(N652),.IN5(n151),.IN6(N669),.Q(n169));
  AOI22X1 U147(.IN1(N499),.IN2(s_qutnt_i[15:15]),.IN3(N516),.IN4(n152),.QN(n166));
  OA22X1 U148(.IN1(n69),.IN2(n153),.IN3(n68),.IN4(n154),.Q(n165));
  AOI22X1 U149(.IN1(N397),.IN2(s_qutnt_i[9:9]),.IN3(N414),.IN4(n155),.QN(n162));
  AOI22X1 U150(.IN1(N448),.IN2(n156),.IN3(N465),.IN4(n157),.QN(n161));
  AO222X1 U152(.IN1(n130),.IN2(N362),.IN3(n131),.IN4(N345),.IN5(n126),.IN6(N379),.Q(n172));
  NAND3X0 U153(.IN1(n173),.IN2(n174),.IN3(n175),.QN(n171));
  AOI222X1 U154(.IN1(n135),.IN2(N430),.IN3(n136),.IN4(N481),.IN5(n137),.IN6(n176),.QN(n175));
  NAND3X0 U155(.IN1(n177),.IN2(n178),.IN3(n179),.QN(n176));
  OA222X1 U156(.IN1(n116),.IN2(n142),.IN3(n85),.IN4(n143),.IN5(n180),.IN6(n145),.Q(n179));
  AO222X1 U157(.IN1(n148),.IN2(N617),.IN3(s_qutnt_i[21:21]),.IN4(N600),.IN5(n149),.IN6(N634),.Q(n182));
  AO222X1 U158(.IN1(N679),.IN2(n75),.IN3(n150),.IN4(N651),.IN5(n151),.IN6(N668),.Q(n181));
  AOI22X1 U159(.IN1(N498),.IN2(s_qutnt_i[15:15]),.IN3(N515),.IN4(n152),.QN(n178));
  OA22X1 U160(.IN1(n110),.IN2(n153),.IN3(n92),.IN4(n154),.Q(n177));
  AOI22X1 U161(.IN1(N396),.IN2(s_qutnt_i[9:9]),.IN3(N413),.IN4(n155),.QN(n174));
  AOI22X1 U162(.IN1(N447),.IN2(n156),.IN3(N464),.IN4(n157),.QN(n173));
  AOI222X1 U163(.IN1(N361),.IN2(n130),.IN3(n185),.IN4(n186),.IN5(N344),.IN6(n131),.QN(n184));
  AOI222X1 U164(.IN1(N327),.IN2(n159),.IN3(N378),.IN4(n126),.IN5(n187),.IN6(n127),.QN(n183));
  OR2X1 U165(.IN1(n188),.IN2(n189),.Q(n187));
  AO222X1 U166(.IN1(n137),.IN2(n190),.IN3(n136),.IN4(N480),.IN5(n135),.IN6(N429),.Q(n189));
  NAND3X0 U167(.IN1(n191),.IN2(n192),.IN3(n193),.QN(n190));
  OA222X1 U168(.IN1(n120),.IN2(n142),.IN3(n87),.IN4(n143),.IN5(n194),.IN6(n145),.Q(n193));
  AO222X1 U169(.IN1(n148),.IN2(N616),.IN3(s_qutnt_i[21:21]),.IN4(N599),.IN5(n149),.IN6(N633),.Q(n196));
  AO222X1 U170(.IN1(N678),.IN2(n75),.IN3(n150),.IN4(N650),.IN5(n151),.IN6(N667),.Q(n195));
  AOI22X1 U171(.IN1(N497),.IN2(s_qutnt_i[15:15]),.IN3(N514),.IN4(n152),.QN(n192));
  OA22X1 U172(.IN1(n111),.IN2(n153),.IN3(n102),.IN4(n154),.Q(n191));
  AO221X1 U173(.IN1(n156),.IN2(N446),.IN3(n157),.IN4(N463),.IN5(n197),.Q(n188));
  AO22X1 U174(.IN1(n155),.IN2(N412),.IN3(s_qutnt_i[9:9]),.IN4(N395),.Q(n197));
  NAND4X0 U176(.IN1(n201),.IN2(n202),.IN3(n203),.IN4(n204),.QN(n198));
  AOI222X1 U177(.IN1(N377),.IN2(n126),.IN3(N343),.IN4(n131),.IN5(N360),.IN6(n130),.QN(n204));
  AO21X1 U178(.IN1(n205),.IN2(n206),.IN3(n321),.Q(n202));
  AOI221X1 U179(.IN1(N462),.IN2(n157),.IN3(N445),.IN4(n156),.IN5(n207),.QN(n206));
  AO22X1 U180(.IN1(N394),.IN2(s_qutnt_i[9:9]),.IN3(N411),.IN4(n155),.Q(n207));
  AOI222X1 U181(.IN1(n135),.IN2(N428),.IN3(n136),.IN4(N479),.IN5(n137),.IN6(n208),.QN(n205));
  NAND3X0 U182(.IN1(n209),.IN2(n210),.IN3(n211),.QN(n208));
  OA222X1 U183(.IN1(n121),.IN2(n142),.IN3(n88),.IN4(n143),.IN5(n212),.IN6(n145),.Q(n211));
  AO222X1 U184(.IN1(n148),.IN2(N615),.IN3(s_qutnt_i[21:21]),.IN4(N598),.IN5(n149),.IN6(N632),.Q(n214));
  AO222X1 U185(.IN1(N677),.IN2(n75),.IN3(n150),.IN4(N649),.IN5(n151),.IN6(N666),.Q(n213));
  AOI22X1 U186(.IN1(N496),.IN2(s_qutnt_i[15:15]),.IN3(N513),.IN4(n152),.QN(n210));
  OA22X1 U187(.IN1(n114),.IN2(n153),.IN3(n107),.IN4(n154),.Q(n209));
  AO22X1 U188(.IN1(n328),.IN2(n215),.IN3(n216),.IN4(n113),.Q(s_r_zeros[0:0]));
  NAND4X0 U189(.IN1(n217),.IN2(n218),.IN3(N304),.IN4(n219),.QN(n215));
  AOI222X1 U190(.IN1(N376),.IN2(n126),.IN3(N342),.IN4(n131),.IN5(N359),.IN6(n130),.QN(n219));
  AND2X1 U191(.IN1(n220),.IN2(n221),.Q(n130));
  AO21X1 U192(.IN1(n223),.IN2(n224),.IN3(n321),.Q(n218));
  AOI221X1 U193(.IN1(N461),.IN2(n157),.IN3(N444),.IN4(n156),.IN5(n225),.QN(n224));
  AO22X1 U194(.IN1(N393),.IN2(s_qutnt_i[9:9]),.IN3(N410),.IN4(n155),.Q(n225));
  AND2X1 U195(.IN1(n228),.IN2(n229),.Q(n157));
  AOI222X1 U196(.IN1(n135),.IN2(N427),.IN3(n136),.IN4(N478),.IN5(n137),.IN6(n230),.QN(n223));
  NAND3X0 U197(.IN1(n231),.IN2(n232),.IN3(n233),.QN(n230));
  OA222X1 U198(.IN1(N540),.IN2(n142),.IN3(n89),.IN4(n143),.IN5(n234),.IN6(n145),.Q(n233));
  AO222X1 U199(.IN1(n148),.IN2(N614),.IN3(s_qutnt_i[21:21]),.IN4(N597),.IN5(n149),.IN6(N631),.Q(n236));
  AND2X1 U200(.IN1(n237),.IN2(n238),.Q(n149));
  AO222X1 U201(.IN1(N676),.IN2(n75),.IN3(n150),.IN4(N648),.IN5(n151),.IN6(N665),.Q(n235));
  AND2X1 U202(.IN1(n239),.IN2(n240),.Q(n151));
  NAND3X0 U203(.IN1(n60),.IN2(\sub_1_root_sub_150_2/CI ),.IN3(n239),.QN(n240));
  AOI22X1 U204(.IN1(N495),.IN2(s_qutnt_i[15:15]),.IN3(N512),.IN4(n152),.QN(n232));
  OA22X1 U205(.IN1(N557),.IN2(n153),.IN3(N574),.IN4(n154),.Q(n231));
  OR2X1 U206(.IN1(n243),.IN2(n244),.Q(n153));
  AND2X1 U207(.IN1(n226),.IN2(n227),.Q(n135));
  AND2X1 U208(.IN1(n327),.IN2(n222),.Q(n159));
  AND2X1 U209(.IN1(s_fraco2[9:9]),.IN2(n245),.Q(s_output_o[9:9]));
  AND2X1 U210(.IN1(s_fraco2[8:8]),.IN2(n14),.Q(s_output_o[8:8]));
  AND2X1 U211(.IN1(s_fraco2[7:7]),.IN2(n245),.Q(s_output_o[7:7]));
  AND2X1 U212(.IN1(s_fraco2[6:6]),.IN2(n14),.Q(s_output_o[6:6]));
  AND2X1 U213(.IN1(s_fraco2[5:5]),.IN2(n245),.Q(s_output_o[5:5]));
  AND2X1 U214(.IN1(s_fraco2[4:4]),.IN2(n14),.Q(s_output_o[4:4]));
  AND2X1 U215(.IN1(s_fraco2[3:3]),.IN2(n245),.Q(s_output_o[3:3]));
  AND2X1 U216(.IN1(s_fraco2[2:2]),.IN2(n14),.Q(s_output_o[2:2]));
  NAND3X0 U217(.IN1(n247),.IN2(n249),.IN3(s_fraco2[22:22]),.QN(n248));
  AOI222X1 U218(.IN1(n250),.IN2(n251),.IN3(n252),.IN4(n253),.IN5(n254),.IN6(n255),.QN(n246));
  OR2X1 U219(.IN1(n256),.IN2(n250),.Q(n253));
  AND2X1 U220(.IN1(s_fraco2[21:21]),.IN2(n245),.Q(s_output_o[21:21]));
  AND2X1 U221(.IN1(s_fraco2[20:20]),.IN2(n14),.Q(s_output_o[20:20]));
  AND2X1 U222(.IN1(s_fraco2[1:1]),.IN2(n245),.Q(s_output_o[1:1]));
  AND2X1 U223(.IN1(s_fraco2[19:19]),.IN2(n14),.Q(s_output_o[19:19]));
  AND2X1 U224(.IN1(s_fraco2[18:18]),.IN2(n245),.Q(s_output_o[18:18]));
  AND2X1 U225(.IN1(s_fraco2[17:17]),.IN2(n14),.Q(s_output_o[17:17]));
  AND2X1 U226(.IN1(s_fraco2[16:16]),.IN2(n245),.Q(s_output_o[16:16]));
  AND2X1 U227(.IN1(s_fraco2[15:15]),.IN2(n14),.Q(s_output_o[15:15]));
  AND2X1 U228(.IN1(s_fraco2[14:14]),.IN2(n245),.Q(s_output_o[14:14]));
  AND2X1 U229(.IN1(s_fraco2[13:13]),.IN2(n14),.Q(s_output_o[13:13]));
  AND2X1 U230(.IN1(s_fraco2[12:12]),.IN2(n245),.Q(s_output_o[12:12]));
  AND2X1 U231(.IN1(s_fraco2[11:11]),.IN2(n14),.Q(s_output_o[11:11]));
  AND2X1 U232(.IN1(s_fraco2[10:10]),.IN2(n245),.Q(s_output_o[10:10]));
  AND2X1 U233(.IN1(s_fraco2[0:0]),.IN2(n14),.Q(s_output_o[0:0]));
  NOR3X0 U234(.IN1(n250),.IN2(n252),.IN3(n74),.QN(n249));
  AO22X1 U235(.IN1(N664),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N653),.Q(N670));
  AO22X1 U236(.IN1(N663),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N652),.Q(N669));
  AO22X1 U237(.IN1(N662),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N651),.Q(N668));
  AO22X1 U238(.IN1(N661),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N650),.Q(N667));
  AO22X1 U239(.IN1(N660),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N649),.Q(N666));
  AO22X1 U240(.IN1(N659),.IN2(n60),.IN3(s_qutnt_i[25:25]),.IN4(N648),.Q(N665));
  AO22X1 U241(.IN1(N647),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N636),.Q(N653));
  AO22X1 U242(.IN1(N646),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N635),.Q(N652));
  AO22X1 U243(.IN1(N645),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N634),.Q(N651));
  AO22X1 U244(.IN1(N644),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N633),.Q(N650));
  AO22X1 U245(.IN1(N643),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N632),.Q(N649));
  AO22X1 U246(.IN1(N642),.IN2(n61),.IN3(s_qutnt_i[24:24]),.IN4(N631),.Q(N648));
  AO22X1 U247(.IN1(N630),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N619),.Q(N636));
  AO22X1 U248(.IN1(N629),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N618),.Q(N635));
  AO22X1 U249(.IN1(N628),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N617),.Q(N634));
  AO22X1 U250(.IN1(N627),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N616),.Q(N633));
  AO22X1 U251(.IN1(N626),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N615),.Q(N632));
  AO22X1 U252(.IN1(N625),.IN2(n62),.IN3(s_qutnt_i[23:23]),.IN4(N614),.Q(N631));
  AO22X1 U253(.IN1(N613),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N602),.Q(N619));
  AO22X1 U254(.IN1(N612),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N601),.Q(N618));
  AO22X1 U255(.IN1(N611),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N600),.Q(N617));
  AO22X1 U256(.IN1(N610),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N599),.Q(N616));
  AO22X1 U257(.IN1(N609),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N598),.Q(N615));
  AO22X1 U258(.IN1(N608),.IN2(n63),.IN3(s_qutnt_i[22:22]),.IN4(N597),.Q(N614));
  AO22X1 U259(.IN1(N596),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N585),.Q(N602));
  AO22X1 U260(.IN1(N595),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N584),.Q(N601));
  AO22X1 U261(.IN1(N594),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N583),.Q(N600));
  AO22X1 U262(.IN1(N593),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N582),.Q(N599));
  AO22X1 U263(.IN1(N592),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N581),.Q(N598));
  AO22X1 U264(.IN1(n89),.IN2(n64),.IN3(s_qutnt_i[21:21]),.IN4(N580),.Q(N597));
  AO22X1 U265(.IN1(N579),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N568),.Q(N585));
  AO22X1 U266(.IN1(N578),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N567),.Q(N584));
  AO22X1 U267(.IN1(N577),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N566),.Q(N583));
  AO22X1 U268(.IN1(N576),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N565),.Q(N582));
  AO22X1 U269(.IN1(N575),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N564),.Q(N581));
  AO22X1 U270(.IN1(N574),.IN2(n71),.IN3(s_qutnt_i[20:20]),.IN4(N563),.Q(N580));
  AO22X1 U271(.IN1(N562),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N551),.Q(N568));
  AO22X1 U272(.IN1(N561),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N550),.Q(N567));
  AO22X1 U273(.IN1(N560),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N549),.Q(N566));
  AO22X1 U274(.IN1(N559),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N548),.Q(N565));
  AO22X1 U275(.IN1(N558),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N547),.Q(N564));
  AO22X1 U276(.IN1(N557),.IN2(n79),.IN3(s_qutnt_i[19:19]),.IN4(N546),.Q(N563));
  AO22X1 U277(.IN1(N545),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N534),.Q(N551));
  AO22X1 U278(.IN1(N544),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N533),.Q(N550));
  AO22X1 U279(.IN1(N543),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N532),.Q(N549));
  AO22X1 U280(.IN1(N542),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N531),.Q(N548));
  AO22X1 U281(.IN1(N541),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N530),.Q(N547));
  AO22X1 U282(.IN1(N540),.IN2(n86),.IN3(s_qutnt_i[18:18]),.IN4(N529),.Q(N546));
  AO22X1 U283(.IN1(N528),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N517),.Q(N534));
  AO22X1 U284(.IN1(N527),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N516),.Q(N533));
  AO22X1 U285(.IN1(N526),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N515),.Q(N532));
  AO22X1 U286(.IN1(N525),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N514),.Q(N531));
  AO22X1 U287(.IN1(N524),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N513),.Q(N530));
  AO22X1 U288(.IN1(N523),.IN2(n93),.IN3(s_qutnt_i[17:17]),.IN4(N512),.Q(N529));
  AO22X1 U289(.IN1(N511),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N500),.Q(N517));
  AO22X1 U290(.IN1(N510),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N499),.Q(N516));
  AO22X1 U291(.IN1(N509),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N498),.Q(N515));
  AO22X1 U292(.IN1(N508),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N497),.Q(N514));
  AO22X1 U293(.IN1(N507),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N496),.Q(N513));
  AO22X1 U294(.IN1(N506),.IN2(n94),.IN3(s_qutnt_i[16:16]),.IN4(N495),.Q(N512));
  AO22X1 U295(.IN1(N494),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N483),.Q(N500));
  AO22X1 U296(.IN1(N493),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N482),.Q(N499));
  AO22X1 U297(.IN1(N492),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N481),.Q(N498));
  AO22X1 U298(.IN1(N491),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N480),.Q(N497));
  AO22X1 U299(.IN1(N490),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N479),.Q(N496));
  AO22X1 U300(.IN1(N489),.IN2(n95),.IN3(s_qutnt_i[15:15]),.IN4(N478),.Q(N495));
  AO22X1 U301(.IN1(N477),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N466),.Q(N483));
  AO22X1 U302(.IN1(N476),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N465),.Q(N482));
  AO22X1 U303(.IN1(N475),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N464),.Q(N481));
  AO22X1 U304(.IN1(N474),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N463),.Q(N480));
  AO22X1 U305(.IN1(N473),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N462),.Q(N479));
  AO22X1 U306(.IN1(N472),.IN2(n96),.IN3(s_qutnt_i[14:14]),.IN4(N461),.Q(N478));
  AO22X1 U307(.IN1(N460),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N449),.Q(N466));
  AO22X1 U308(.IN1(N459),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N448),.Q(N465));
  AO22X1 U309(.IN1(N458),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N447),.Q(N464));
  AO22X1 U310(.IN1(N457),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N446),.Q(N463));
  AO22X1 U311(.IN1(N456),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N445),.Q(N462));
  AO22X1 U312(.IN1(N455),.IN2(n97),.IN3(s_qutnt_i[13:13]),.IN4(N444),.Q(N461));
  AO22X1 U313(.IN1(N443),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N432),.Q(N449));
  AO22X1 U314(.IN1(N442),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N431),.Q(N448));
  AO22X1 U315(.IN1(N441),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N430),.Q(N447));
  AO22X1 U316(.IN1(N440),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N429),.Q(N446));
  AO22X1 U317(.IN1(N439),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N428),.Q(N445));
  AO22X1 U318(.IN1(N438),.IN2(n98),.IN3(s_qutnt_i[12:12]),.IN4(N427),.Q(N444));
  AO22X1 U319(.IN1(N426),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N415),.Q(N432));
  AO22X1 U320(.IN1(N425),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N414),.Q(N431));
  AO22X1 U321(.IN1(N424),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N413),.Q(N430));
  AO22X1 U322(.IN1(N423),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N412),.Q(N429));
  AO22X1 U323(.IN1(N422),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N411),.Q(N428));
  AO22X1 U324(.IN1(N421),.IN2(n99),.IN3(s_qutnt_i[11:11]),.IN4(N410),.Q(N427));
  AO22X1 U325(.IN1(N409),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N398),.Q(N415));
  AO22X1 U326(.IN1(N408),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N397),.Q(N414));
  AO22X1 U327(.IN1(N407),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N396),.Q(N413));
  AO22X1 U328(.IN1(N406),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N395),.Q(N412));
  AO22X1 U329(.IN1(N405),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N394),.Q(N411));
  AO22X1 U330(.IN1(N404),.IN2(n100),.IN3(s_qutnt_i[10:10]),.IN4(N393),.Q(N410));
  AO22X1 U331(.IN1(N392),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N381),.Q(N398));
  AO22X1 U332(.IN1(N391),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N380),.Q(N397));
  AO22X1 U333(.IN1(N390),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N379),.Q(N396));
  AO22X1 U334(.IN1(N389),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N378),.Q(N395));
  AO22X1 U335(.IN1(N388),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N377),.Q(N394));
  AO22X1 U336(.IN1(N387),.IN2(n101),.IN3(s_qutnt_i[9:9]),.IN4(N376),.Q(N393));
  AO22X1 U337(.IN1(N375),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N364),.Q(N381));
  AO22X1 U338(.IN1(N374),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N363),.Q(N380));
  AO22X1 U339(.IN1(N373),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N362),.Q(N379));
  AO22X1 U340(.IN1(N372),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N361),.Q(N378));
  AO22X1 U341(.IN1(N371),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N360),.Q(N377));
  AO22X1 U342(.IN1(N370),.IN2(n103),.IN3(s_qutnt_i[8:8]),.IN4(N359),.Q(N376));
  AO22X1 U343(.IN1(N358),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(n12),.Q(N364));
  AO22X1 U344(.IN1(N357),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(N346),.Q(N363));
  AO22X1 U345(.IN1(N356),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(N345),.Q(N362));
  AO22X1 U346(.IN1(N355),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(N344),.Q(N361));
  AO22X1 U347(.IN1(N354),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(N343),.Q(N360));
  AO22X1 U348(.IN1(N353),.IN2(n104),.IN3(s_qutnt_i[7:7]),.IN4(N342),.Q(N359));
  AO22X1 U350(.IN1(N340),.IN2(n105),.IN3(s_qutnt_i[6:6]),.IN4(N329),.Q(N346));
  AO22X1 U351(.IN1(N339),.IN2(n105),.IN3(s_qutnt_i[6:6]),.IN4(N328),.Q(N345));
  AO22X1 U352(.IN1(N338),.IN2(n105),.IN3(s_qutnt_i[6:6]),.IN4(N327),.Q(N344));
  AO22X1 U353(.IN1(N337),.IN2(n105),.IN3(s_qutnt_i[6:6]),.IN4(N326),.Q(N343));
  AO22X1 U354(.IN1(N336),.IN2(n105),.IN3(s_qutnt_i[6:6]),.IN4(N325),.Q(N342));
  AO22X1 U357(.IN1(N322),.IN2(n106),.IN3(N312),.IN4(s_qutnt_i[5:5]),.Q(N328));
  AO22X1 U358(.IN1(N321),.IN2(n106),.IN3(s_qutnt_i[5:5]),.IN4(N311),.Q(N327));
  AO22X1 U359(.IN1(N320),.IN2(n106),.IN3(s_qutnt_i[5:5]),.IN4(N310),.Q(N326));
  AO22X1 U360(.IN1(N319),.IN2(n106),.IN3(s_qutnt_i[5:5]),.IN4(N309),.Q(N325));
  AND2X1 U362(.IN1(N307),.IN2(n108),.Q(N312));
  AO22X1 U363(.IN1(N306),.IN2(n108),.IN3(s_qutnt_i[4:4]),.IN4(N297),.Q(N311));
  AO22X1 U364(.IN1(N305),.IN2(n108),.IN3(s_qutnt_i[4:4]),.IN4(\add_105_I5_L14036_C191/A[1] ),.Q(N310));
  AO22X1 U365(.IN1(N304),.IN2(n108),.IN3(s_qutnt_i[4:4]),.IN4(N295),.Q(N309));
  AND2X1 U367(.IN1(n258),.IN2(n259),.Q(N297));
  XNOR2X1 U368(.IN1(n258),.IN2(n259),.Q(n203));
  AO21X1 U369(.IN1(n216),.IN2(n112),.IN3(n199),.Q(n259));
  XOR2X1 U370(.IN1(n260),.IN2(s_qutnt_i[3:3]),.Q(N295));
  XNOR2X1 U371(.IN1(n112),.IN2(n216),.Q(n260));
  XNOR2X1 U372(.IN1(n113),.IN2(s_qutnt_i[1:1]),.Q(n216));
  AO22X1 U373(.IN1(N210),.IN2(n23),.IN3(N237),.IN4(n22),.Q(N264));
  AO22X1 U374(.IN1(N209),.IN2(n23),.IN3(N236),.IN4(n22),.Q(N263));
  AO22X1 U375(.IN1(N208),.IN2(n23),.IN3(N235),.IN4(n261),.Q(N262));
  AO22X1 U376(.IN1(N207),.IN2(n23),.IN3(N234),.IN4(n261),.Q(N261));
  AO22X1 U377(.IN1(N206),.IN2(n23),.IN3(N233),.IN4(n261),.Q(N260));
  AO22X1 U378(.IN1(N205),.IN2(n23),.IN3(N232),.IN4(n261),.Q(N259));
  AO22X1 U379(.IN1(N204),.IN2(n23),.IN3(N231),.IN4(n261),.Q(N258));
  AO22X1 U380(.IN1(N203),.IN2(n23),.IN3(N230),.IN4(n261),.Q(N257));
  AO22X1 U381(.IN1(N202),.IN2(n23),.IN3(N229),.IN4(n261),.Q(N256));
  AO22X1 U382(.IN1(N201),.IN2(n23),.IN3(N228),.IN4(n261),.Q(N255));
  AO22X1 U383(.IN1(N200),.IN2(n23),.IN3(N227),.IN4(n261),.Q(N254));
  AO22X1 U384(.IN1(N199),.IN2(n23),.IN3(N226),.IN4(n261),.Q(N253));
  AO22X1 U385(.IN1(N198),.IN2(n23),.IN3(N225),.IN4(n261),.Q(N252));
  AO22X1 U386(.IN1(N197),.IN2(n23),.IN3(N224),.IN4(n261),.Q(N251));
  AO22X1 U387(.IN1(N196),.IN2(n23),.IN3(N223),.IN4(n261),.Q(N250));
  AO22X1 U388(.IN1(N195),.IN2(n23),.IN3(N222),.IN4(n22),.Q(N249));
  AO22X1 U389(.IN1(N194),.IN2(n23),.IN3(N221),.IN4(n22),.Q(N248));
  AO22X1 U390(.IN1(N193),.IN2(n23),.IN3(N220),.IN4(n22),.Q(N247));
  AO22X1 U391(.IN1(N192),.IN2(n24),.IN3(N219),.IN4(n22),.Q(N246));
  AO22X1 U392(.IN1(N191),.IN2(n24),.IN3(N218),.IN4(n22),.Q(N245));
  AO22X1 U393(.IN1(N190),.IN2(n24),.IN3(N217),.IN4(n22),.Q(N244));
  AO22X1 U394(.IN1(N189),.IN2(n24),.IN3(N216),.IN4(n22),.Q(N243));
  AO22X1 U395(.IN1(N188),.IN2(n24),.IN3(N215),.IN4(n22),.Q(N242));
  AO22X1 U396(.IN1(N187),.IN2(n24),.IN3(N214),.IN4(n22),.Q(N241));
  AO22X1 U397(.IN1(N186),.IN2(n24),.IN3(N213),.IN4(n22),.Q(N240));
  AO22X1 U398(.IN1(N185),.IN2(n24),.IN3(N212),.IN4(n22),.Q(N239));
  AO22X1 U399(.IN1(N184),.IN2(n23),.IN3(N211),.IN4(n22),.Q(N238));
  NOR4X0 U400(.IN1(s_shr1[2:2]),.IN2(s_shr1[1:1]),.IN3(s_shr1[0:0]),.IN4(n262),.QN(n261));
  OR3X1 U401(.IN1(n29),.IN2(n27),.IN3(s_shr1[3:3]),.Q(n262));
  AO21X1 U402(.IN1(N150),.IN2(n52),.IN3(n263),.Q(N177));
  AO21X1 U403(.IN1(N149),.IN2(n52),.IN3(n263),.Q(N176));
  AO21X1 U404(.IN1(N148),.IN2(n52),.IN3(n263),.Q(N175));
  AO21X1 U405(.IN1(N147),.IN2(n52),.IN3(n263),.Q(N174));
  AO21X1 U406(.IN1(N146),.IN2(n52),.IN3(n263),.Q(N173));
  AO21X1 U407(.IN1(N145),.IN2(n52),.IN3(n263),.Q(N172));
  AND2X1 U408(.IN1(N151),.IN2(n52),.Q(n263));
  AND2X1 U409(.IN1(n264),.IN2(s_exp_10b[5:5]),.Q(N167));
  AND2X1 U410(.IN1(n264),.IN2(s_exp_10b[4:4]),.Q(N166));
  AND3X1 U411(.IN1(n264),.IN2(\sub_1_root_sub_150_2/CI ),.IN3(n53),.Q(N161));
  NOR4X0 U412(.IN1(n266),.IN2(n267),.IN3(s_exp_10b[5:5]),.IN4(s_exp_10b[4:4]),.QN(n265));
  NAND3X0 U413(.IN1(n54),.IN2(n53),.IN3(n55),.QN(n267));
  NAND4X0 U414(.IN1(n1),.IN2(n31),.IN3(n57),.IN4(n56),.QN(n266));
  NOR4X0 U415(.IN1(s_opa_i[27:27]),.IN2(s_opa_i[26:26]),.IN3(n269),.IN4(n270),.QN(n254));
  OR4X1 U416(.IN1(s_opa_i[23:23]),.IN2(n256),.IN3(s_opa_i[25:25]),.IN4(s_opa_i[24:24]),.Q(n270));
  NAND4X0 U417(.IN1(n271),.IN2(n272),.IN3(n273),.IN4(n274),.QN(n256));
  NOR4X0 U418(.IN1(n275),.IN2(s_opa_i[4:4]),.IN3(s_opa_i[6:6]),.IN4(s_opa_i[5:5]),.QN(n274));
  OR3X1 U419(.IN1(s_opa_i[9:9]),.IN2(s_opa_i[8:8]),.IN3(s_opa_i[7:7]),.Q(n275));
  NOR4X0 U420(.IN1(n276),.IN2(s_opa_i[1:1]),.IN3(s_opa_i[21:21]),.IN4(s_opa_i[20:20]),.QN(n273));
  OR3X1 U421(.IN1(s_opa_i[3:3]),.IN2(s_opa_i[2:2]),.IN3(s_opa_i[22:22]),.Q(n276));
  NOR4X0 U422(.IN1(n277),.IN2(s_opa_i[14:14]),.IN3(s_opa_i[16:16]),.IN4(s_opa_i[15:15]),.QN(n272));
  OR3X1 U423(.IN1(s_opa_i[19:19]),.IN2(s_opa_i[18:18]),.IN3(s_opa_i[17:17]),.Q(n277));
  NOR4X0 U424(.IN1(n278),.IN2(s_opa_i[11:11]),.IN3(s_opa_i[13:13]),.IN4(s_opa_i[12:12]),.QN(n271));
  OR2X1 U425(.IN1(s_opa_i[10:10]),.IN2(s_opa_i[0:0]),.Q(n278));
  OR3X1 U426(.IN1(s_opa_i[30:30]),.IN2(s_opa_i[29:29]),.IN3(s_opa_i[28:28]),.Q(n269));
  NOR3X0 U427(.IN1(n279),.IN2(N1025),.IN3(n280),.QN(n268));
  NOR3X0 U428(.IN1(n257),.IN2(n252),.IN3(n250),.QN(n280));
  NAND4X0 U429(.IN1(s_expb[7:7]),.IN2(s_expb[6:6]),.IN3(s_expb[5:5]),.IN4(s_expb[4:4]),.QN(n282));
  NAND4X0 U430(.IN1(s_expb[3:3]),.IN2(s_expb[2:2]),.IN3(s_expb[1:1]),.IN4(s_expb[0:0]),.QN(n281));
  NAND4X0 U431(.IN1(s_expa[7:7]),.IN2(s_expa[6:6]),.IN3(s_expa[5:5]),.IN4(s_expa[4:4]),.QN(n284));
  NAND4X0 U432(.IN1(s_expa[3:3]),.IN2(s_expa[2:2]),.IN3(s_expa[1:1]),.IN4(s_expa[0:0]),.QN(n283));
  NOR3X0 U433(.IN1(s_expo3[8:8]),.IN2(n255),.IN3(n285),.QN(n257));
  NAND4X0 U434(.IN1(s_expo3[7:7]),.IN2(s_expo3[6:6]),.IN3(s_expo3[5:5]),.IN4(s_expo3[4:4]),.QN(n287));
  NAND4X0 U435(.IN1(s_expo3[3:3]),.IN2(s_expo3[2:2]),.IN3(s_expo3[1:1]),.IN4(s_expo3[0:0]),.QN(n286));
  NOR4X0 U436(.IN1(s_opb_i[27:27]),.IN2(s_opb_i[26:26]),.IN3(n288),.IN4(n289),.QN(n255));
  OR4X1 U437(.IN1(s_opb_i[23:23]),.IN2(n251),.IN3(s_opb_i[25:25]),.IN4(s_opb_i[24:24]),.Q(n289));
  NAND4X0 U438(.IN1(n290),.IN2(n291),.IN3(n292),.IN4(n293),.QN(n251));
  NOR4X0 U439(.IN1(n294),.IN2(s_opb_i[4:4]),.IN3(s_opb_i[6:6]),.IN4(s_opb_i[5:5]),.QN(n293));
  OR3X1 U440(.IN1(s_opb_i[9:9]),.IN2(s_opb_i[8:8]),.IN3(s_opb_i[7:7]),.Q(n294));
  NOR4X0 U441(.IN1(n295),.IN2(s_opb_i[1:1]),.IN3(s_opb_i[21:21]),.IN4(s_opb_i[20:20]),.QN(n292));
  OR3X1 U442(.IN1(s_opb_i[3:3]),.IN2(s_opb_i[2:2]),.IN3(s_opb_i[22:22]),.Q(n295));
  NOR4X0 U443(.IN1(n296),.IN2(s_opb_i[14:14]),.IN3(s_opb_i[16:16]),.IN4(s_opb_i[15:15]),.QN(n291));
  OR3X1 U444(.IN1(s_opb_i[19:19]),.IN2(s_opb_i[18:18]),.IN3(s_opb_i[17:17]),.Q(n296));
  NOR4X0 U445(.IN1(n297),.IN2(s_opb_i[11:11]),.IN3(s_opb_i[13:13]),.IN4(s_opb_i[12:12]),.QN(n290));
  OR2X1 U446(.IN1(s_opb_i[10:10]),.IN2(s_opb_i[0:0]),.Q(n297));
  OR3X1 U447(.IN1(s_opb_i[30:30]),.IN2(s_opb_i[29:29]),.IN3(s_opb_i[28:28]),.Q(n288));
  AO222X1 U448(.IN1(N1087),.IN2(n298),.IN3(s_fraco1[25:25]),.IN4(n21),.IN5(N1088),.IN6(n15),.Q(N1131));
  AO222X1 U449(.IN1(N1086),.IN2(n298),.IN3(s_fraco1[24:24]),.IN4(n21),.IN5(n15),.IN6(N1087),.Q(N1130));
  AO222X1 U450(.IN1(N1085),.IN2(n298),.IN3(s_fraco1[23:23]),.IN4(n21),.IN5(N1086),.IN6(n15),.Q(N1129));
  AO222X1 U451(.IN1(N1084),.IN2(n298),.IN3(s_fraco1[22:22]),.IN4(n21),.IN5(N1085),.IN6(n15),.Q(N1128));
  AO222X1 U452(.IN1(N1083),.IN2(n298),.IN3(s_fraco1[21:21]),.IN4(n21),.IN5(N1084),.IN6(n15),.Q(N1127));
  AO222X1 U453(.IN1(N1082),.IN2(n298),.IN3(s_fraco1[20:20]),.IN4(n21),.IN5(N1083),.IN6(n15),.Q(N1126));
  AO222X1 U454(.IN1(N1081),.IN2(n298),.IN3(s_fraco1[19:19]),.IN4(n21),.IN5(N1082),.IN6(n15),.Q(N1125));
  AO222X1 U455(.IN1(N1080),.IN2(n298),.IN3(s_fraco1[18:18]),.IN4(n21),.IN5(N1081),.IN6(n15),.Q(N1124));
  AO222X1 U456(.IN1(N1079),.IN2(n298),.IN3(s_fraco1[17:17]),.IN4(n21),.IN5(N1080),.IN6(n15),.Q(N1123));
  AO222X1 U457(.IN1(N1078),.IN2(n298),.IN3(s_fraco1[16:16]),.IN4(n21),.IN5(N1079),.IN6(n15),.Q(N1122));
  AO222X1 U458(.IN1(N1077),.IN2(n298),.IN3(s_fraco1[15:15]),.IN4(n21),.IN5(N1078),.IN6(n15),.Q(N1121));
  AO222X1 U459(.IN1(N1076),.IN2(n298),.IN3(s_fraco1[14:14]),.IN4(n21),.IN5(N1077),.IN6(n15),.Q(N1120));
  AO222X1 U460(.IN1(N1075),.IN2(n298),.IN3(s_fraco1[13:13]),.IN4(n21),.IN5(N1076),.IN6(n15),.Q(N1119));
  AO222X1 U461(.IN1(N1074),.IN2(n298),.IN3(s_fraco1[12:12]),.IN4(n21),.IN5(N1075),.IN6(n15),.Q(N1118));
  AO222X1 U462(.IN1(N1073),.IN2(n298),.IN3(s_fraco1[11:11]),.IN4(n21),.IN5(N1074),.IN6(n15),.Q(N1117));
  AO222X1 U463(.IN1(N1072),.IN2(n298),.IN3(s_fraco1[10:10]),.IN4(n21),.IN5(N1073),.IN6(n15),.Q(N1116));
  AO222X1 U464(.IN1(N1071),.IN2(n298),.IN3(s_fraco1[9:9]),.IN4(n21),.IN5(N1072),.IN6(n15),.Q(N1115));
  AO222X1 U465(.IN1(N1070),.IN2(n298),.IN3(s_fraco1[8:8]),.IN4(n21),.IN5(N1071),.IN6(n16),.Q(N1114));
  AO222X1 U466(.IN1(N1069),.IN2(n298),.IN3(s_fraco1[7:7]),.IN4(n21),.IN5(N1070),.IN6(n16),.Q(N1113));
  AO222X1 U467(.IN1(N1068),.IN2(n298),.IN3(s_fraco1[6:6]),.IN4(n21),.IN5(N1069),.IN6(n16),.Q(N1112));
  AO222X1 U468(.IN1(N1067),.IN2(n298),.IN3(s_fraco1[5:5]),.IN4(n21),.IN5(N1068),.IN6(n16),.Q(N1111));
  AO222X1 U469(.IN1(N1066),.IN2(n298),.IN3(s_fraco1[4:4]),.IN4(n21),.IN5(N1067),.IN6(n16),.Q(N1110));
  AO222X1 U470(.IN1(N1065),.IN2(n298),.IN3(s_fraco1[3:3]),.IN4(n21),.IN5(N1066),.IN6(n16),.Q(N1109));
  AO22X1 U471(.IN1(N1099),.IN2(n16),.IN3(s_expo2[8:8]),.IN4(n300),.Q(N1108));
  AO22X1 U472(.IN1(N1098),.IN2(n16),.IN3(s_expo2[7:7]),.IN4(n300),.Q(N1107));
  AO22X1 U473(.IN1(N1097),.IN2(n16),.IN3(s_expo2[6:6]),.IN4(n300),.Q(N1106));
  AO22X1 U474(.IN1(N1096),.IN2(n16),.IN3(s_expo2[5:5]),.IN4(n300),.Q(N1105));
  AO22X1 U475(.IN1(N1095),.IN2(n16),.IN3(s_expo2[4:4]),.IN4(n300),.Q(N1104));
  AO22X1 U476(.IN1(N1094),.IN2(n16),.IN3(s_expo2[3:3]),.IN4(n300),.Q(N1103));
  AO22X1 U477(.IN1(N1093),.IN2(n16),.IN3(s_expo2[2:2]),.IN4(n300),.Q(N1102));
  AO22X1 U478(.IN1(N1092),.IN2(n16),.IN3(s_expo2[1:1]),.IN4(n300),.Q(N1101));
  AO22X1 U479(.IN1(N1091),.IN2(n16),.IN3(s_expo2[0:0]),.IN4(n300),.Q(N1100));
  NAND4X0 U480(.IN1(s_fraco1[2:2]),.IN2(n303),.IN3(n119),.IN4(n118),.QN(n302));
  NAND3X0 U481(.IN1(n124),.IN2(n122),.IN3(n304),.QN(n303));
  NAND3X0 U482(.IN1(\s_rmode_i[1] ),.IN2(n305),.IN3(s_sign_i),.QN(n306));
  NAND3X0 U483(.IN1(n124),.IN2(n123),.IN3(n304),.QN(n279));
  AND4X1 U484(.IN1(n307),.IN2(n308),.IN3(n309),.IN4(n310),.Q(n304));
  NOR4X0 U485(.IN1(n311),.IN2(s_rmndr_i[3:3]),.IN3(s_rmndr_i[5:5]),.IN4(s_rmndr_i[4:4]),.QN(n310));
  OR4X1 U486(.IN1(s_rmndr_i[7:7]),.IN2(s_rmndr_i[6:6]),.IN3(s_rmndr_i[9:9]),.IN4(s_rmndr_i[8:8]),.Q(n311));
  NOR4X0 U487(.IN1(n312),.IN2(s_rmndr_i[21:21]),.IN3(s_rmndr_i[23:23]),.IN4(s_rmndr_i[22:22]),.QN(n309));
  OR4X1 U488(.IN1(s_rmndr_i[25:25]),.IN2(s_rmndr_i[24:24]),.IN3(s_rmndr_i[2:2]),.IN4(s_rmndr_i[26:26]),.Q(n312));
  NOR4X0 U489(.IN1(n313),.IN2(s_rmndr_i[15:15]),.IN3(s_rmndr_i[17:17]),.IN4(s_rmndr_i[16:16]),.QN(n308));
  OR4X1 U490(.IN1(s_rmndr_i[19:19]),.IN2(s_rmndr_i[18:18]),.IN3(s_rmndr_i[20:20]),.IN4(s_rmndr_i[1:1]),.Q(n313));
  NOR4X0 U491(.IN1(n314),.IN2(s_fraco1[0:0]),.IN3(s_rmndr_i[10:10]),.IN4(s_rmndr_i[0:0]),.QN(n307));
  OR4X1 U492(.IN1(s_rmndr_i[12:12]),.IN2(s_rmndr_i[11:11]),.IN3(s_rmndr_i[14:14]),.IN4(s_rmndr_i[13:13]),.Q(n314));
  post_norm_div_DW01_inc_0_inj add_216(.A(s_expo2),.SUM({N1099,N1098,N1097,N1096,N1095,N1094,N1093,N1092,N1091}));
  post_norm_div_DW01_inc_1_inj add_209(.A({1'b0,s_fraco1[26:3]}),.SUM({N1089,N1088,N1087,N1086,N1085,N1084,N1083,N1082,N1081,N1080,N1079,N1078,N1077,N1076,N1075,N1074,N1073,N1072,N1071,N1070,N1069,N1068,N1067,N1066,N1065}));
  HADDX1 desc1760(.A0(N666),.B0(N665),.C1(\add_105_I27_L14036_C191/carry[2] ),.SO(N677));
  HADDX1 desc1761(.A0(N667),.B0(\add_105_I27_L14036_C191/carry[2] ),.C1(\add_105_I27_L14036_C191/carry[3] ),.SO(N678));
  HADDX1 desc1762(.A0(N668),.B0(\add_105_I27_L14036_C191/carry[3] ),.C1(\add_105_I27_L14036_C191/carry[4] ),.SO(N679));
  HADDX1 desc1763(.A0(N669),.B0(\add_105_I27_L14036_C191/carry[4] ),.C1(\add_105_I27_L14036_C191/carry[5] ),.SO(N680));
  HADDX1 desc1764(.A0(N649),.B0(N648),.C1(\add_105_I26_L14036_C191/carry[2] ),.SO(N660));
  HADDX1 desc1765(.A0(N650),.B0(\add_105_I26_L14036_C191/carry[2] ),.C1(\add_105_I26_L14036_C191/carry[3] ),.SO(N661));
  HADDX1 desc1766(.A0(N651),.B0(\add_105_I26_L14036_C191/carry[3] ),.C1(\add_105_I26_L14036_C191/carry[4] ),.SO(N662));
  HADDX1 desc1767(.A0(N652),.B0(\add_105_I26_L14036_C191/carry[4] ),.C1(\add_105_I26_L14036_C191/carry[5] ),.SO(N663));
  HADDX1 desc1768(.A0(N632),.B0(N631),.C1(\add_105_I25_L14036_C191/carry[2] ),.SO(N643));
  HADDX1 desc1769(.A0(N633),.B0(\add_105_I25_L14036_C191/carry[2] ),.C1(\add_105_I25_L14036_C191/carry[3] ),.SO(N644));
  HADDX1 desc1770(.A0(N634),.B0(\add_105_I25_L14036_C191/carry[3] ),.C1(\add_105_I25_L14036_C191/carry[4] ),.SO(N645));
  HADDX1 desc1771(.A0(N635),.B0(\add_105_I25_L14036_C191/carry[4] ),.C1(\add_105_I25_L14036_C191/carry[5] ),.SO(N646));
  HADDX1 desc1772(.A0(N615),.B0(N614),.C1(\add_105_I24_L14036_C191/carry[2] ),.SO(N626));
  HADDX1 desc1773(.A0(N616),.B0(\add_105_I24_L14036_C191/carry[2] ),.C1(\add_105_I24_L14036_C191/carry[3] ),.SO(N627));
  HADDX1 desc1774(.A0(N617),.B0(\add_105_I24_L14036_C191/carry[3] ),.C1(\add_105_I24_L14036_C191/carry[4] ),.SO(N628));
  HADDX1 desc1775(.A0(N618),.B0(\add_105_I24_L14036_C191/carry[4] ),.C1(\add_105_I24_L14036_C191/carry[5] ),.SO(N629));
  HADDX1 desc1776(.A0(N598),.B0(N597),.C1(\add_105_I23_L14036_C191/carry[2] ),.SO(N609));
  HADDX1 desc1777(.A0(N599),.B0(\add_105_I23_L14036_C191/carry[2] ),.C1(\add_105_I23_L14036_C191/carry[3] ),.SO(N610));
  HADDX1 desc1778(.A0(N600),.B0(\add_105_I23_L14036_C191/carry[3] ),.C1(\add_105_I23_L14036_C191/carry[4] ),.SO(N611));
  HADDX1 desc1779(.A0(N601),.B0(\add_105_I23_L14036_C191/carry[4] ),.C1(\add_105_I23_L14036_C191/carry[5] ),.SO(N612));
  HADDX1 desc1780(.A0(N581),.B0(N580),.C1(\add_105_I22_L14036_C191/carry[2] ),.SO(N592));
  HADDX1 desc1781(.A0(N582),.B0(\add_105_I22_L14036_C191/carry[2] ),.C1(\add_105_I22_L14036_C191/carry[3] ),.SO(N593));
  HADDX1 desc1782(.A0(N583),.B0(\add_105_I22_L14036_C191/carry[3] ),.C1(\add_105_I22_L14036_C191/carry[4] ),.SO(N594));
  HADDX1 desc1783(.A0(N584),.B0(\add_105_I22_L14036_C191/carry[4] ),.C1(\add_105_I22_L14036_C191/carry[5] ),.SO(N595));
  HADDX1 desc1784(.A0(N564),.B0(N563),.C1(\add_105_I21_L14036_C191/carry[2] ),.SO(N575));
  HADDX1 desc1785(.A0(N565),.B0(\add_105_I21_L14036_C191/carry[2] ),.C1(\add_105_I21_L14036_C191/carry[3] ),.SO(N576));
  HADDX1 desc1786(.A0(N566),.B0(\add_105_I21_L14036_C191/carry[3] ),.C1(\add_105_I21_L14036_C191/carry[4] ),.SO(N577));
  HADDX1 desc1787(.A0(N567),.B0(\add_105_I21_L14036_C191/carry[4] ),.C1(\add_105_I21_L14036_C191/carry[5] ),.SO(N578));
  HADDX1 desc1788(.A0(N547),.B0(N546),.C1(\add_105_I20_L14036_C191/carry[2] ),.SO(N558));
  HADDX1 desc1789(.A0(N548),.B0(\add_105_I20_L14036_C191/carry[2] ),.C1(\add_105_I20_L14036_C191/carry[3] ),.SO(N559));
  HADDX1 desc1790(.A0(N549),.B0(\add_105_I20_L14036_C191/carry[3] ),.C1(\add_105_I20_L14036_C191/carry[4] ),.SO(N560));
  HADDX1 desc1791(.A0(N550),.B0(\add_105_I20_L14036_C191/carry[4] ),.C1(\add_105_I20_L14036_C191/carry[5] ),.SO(N561));
  HADDX1 desc1792(.A0(N530),.B0(N529),.C1(\add_105_I19_L14036_C191/carry[2] ),.SO(N541));
  HADDX1 desc1793(.A0(N531),.B0(\add_105_I19_L14036_C191/carry[2] ),.C1(\add_105_I19_L14036_C191/carry[3] ),.SO(N542));
  HADDX1 desc1794(.A0(N532),.B0(\add_105_I19_L14036_C191/carry[3] ),.C1(\add_105_I19_L14036_C191/carry[4] ),.SO(N543));
  HADDX1 desc1795(.A0(N533),.B0(\add_105_I19_L14036_C191/carry[4] ),.C1(\add_105_I19_L14036_C191/carry[5] ),.SO(N544));
  HADDX1 desc1796(.A0(N513),.B0(N512),.C1(\add_105_I18_L14036_C191/carry[2] ),.SO(N524));
  HADDX1 desc1797(.A0(N514),.B0(\add_105_I18_L14036_C191/carry[2] ),.C1(\add_105_I18_L14036_C191/carry[3] ),.SO(N525));
  HADDX1 desc1798(.A0(N515),.B0(\add_105_I18_L14036_C191/carry[3] ),.C1(\add_105_I18_L14036_C191/carry[4] ),.SO(N526));
  HADDX1 desc1799(.A0(N516),.B0(\add_105_I18_L14036_C191/carry[4] ),.C1(\add_105_I18_L14036_C191/carry[5] ),.SO(N527));
  HADDX1 desc1800(.A0(N496),.B0(N495),.C1(\add_105_I17_L14036_C191/carry[2] ),.SO(N507));
  HADDX1 desc1801(.A0(N497),.B0(\add_105_I17_L14036_C191/carry[2] ),.C1(\add_105_I17_L14036_C191/carry[3] ),.SO(N508));
  HADDX1 desc1802(.A0(N498),.B0(\add_105_I17_L14036_C191/carry[3] ),.C1(\add_105_I17_L14036_C191/carry[4] ),.SO(N509));
  HADDX1 desc1803(.A0(N499),.B0(\add_105_I17_L14036_C191/carry[4] ),.C1(\add_105_I17_L14036_C191/carry[5] ),.SO(N510));
  HADDX1 desc1804(.A0(N479),.B0(N478),.C1(\add_105_I16_L14036_C191/carry[2] ),.SO(N490));
  HADDX1 desc1805(.A0(N480),.B0(\add_105_I16_L14036_C191/carry[2] ),.C1(\add_105_I16_L14036_C191/carry[3] ),.SO(N491));
  HADDX1 desc1806(.A0(N481),.B0(\add_105_I16_L14036_C191/carry[3] ),.C1(\add_105_I16_L14036_C191/carry[4] ),.SO(N492));
  HADDX1 desc1807(.A0(N482),.B0(\add_105_I16_L14036_C191/carry[4] ),.C1(\add_105_I16_L14036_C191/carry[5] ),.SO(N493));
  HADDX1 desc1808(.A0(N462),.B0(N461),.C1(\add_105_I15_L14036_C191/carry[2] ),.SO(N473));
  HADDX1 desc1809(.A0(N463),.B0(\add_105_I15_L14036_C191/carry[2] ),.C1(\add_105_I15_L14036_C191/carry[3] ),.SO(N474));
  HADDX1 desc1810(.A0(N464),.B0(\add_105_I15_L14036_C191/carry[3] ),.C1(\add_105_I15_L14036_C191/carry[4] ),.SO(N475));
  HADDX1 desc1811(.A0(N465),.B0(\add_105_I15_L14036_C191/carry[4] ),.C1(\add_105_I15_L14036_C191/carry[5] ),.SO(N476));
  HADDX1 desc1812(.A0(N445),.B0(N444),.C1(\add_105_I14_L14036_C191/carry[2] ),.SO(N456));
  HADDX1 desc1813(.A0(N446),.B0(\add_105_I14_L14036_C191/carry[2] ),.C1(\add_105_I14_L14036_C191/carry[3] ),.SO(N457));
  HADDX1 desc1814(.A0(N447),.B0(\add_105_I14_L14036_C191/carry[3] ),.C1(\add_105_I14_L14036_C191/carry[4] ),.SO(N458));
  HADDX1 desc1815(.A0(N448),.B0(\add_105_I14_L14036_C191/carry[4] ),.C1(\add_105_I14_L14036_C191/carry[5] ),.SO(N459));
  HADDX1 desc1816(.A0(N428),.B0(N427),.C1(\add_105_I13_L14036_C191/carry[2] ),.SO(N439));
  HADDX1 desc1817(.A0(N429),.B0(\add_105_I13_L14036_C191/carry[2] ),.C1(\add_105_I13_L14036_C191/carry[3] ),.SO(N440));
  HADDX1 desc1818(.A0(N430),.B0(\add_105_I13_L14036_C191/carry[3] ),.C1(\add_105_I13_L14036_C191/carry[4] ),.SO(N441));
  HADDX1 desc1819(.A0(N431),.B0(\add_105_I13_L14036_C191/carry[4] ),.C1(\add_105_I13_L14036_C191/carry[5] ),.SO(N442));
  HADDX1 desc1820(.A0(N411),.B0(N410),.C1(\add_105_I12_L14036_C191/carry[2] ),.SO(N422));
  HADDX1 desc1821(.A0(N412),.B0(\add_105_I12_L14036_C191/carry[2] ),.C1(\add_105_I12_L14036_C191/carry[3] ),.SO(N423));
  HADDX1 desc1822(.A0(N413),.B0(\add_105_I12_L14036_C191/carry[3] ),.C1(\add_105_I12_L14036_C191/carry[4] ),.SO(N424));
  HADDX1 desc1823(.A0(N414),.B0(\add_105_I12_L14036_C191/carry[4] ),.C1(\add_105_I12_L14036_C191/carry[5] ),.SO(N425));
  HADDX1 desc1824(.A0(N394),.B0(N393),.C1(\add_105_I11_L14036_C191/carry[2] ),.SO(N405));
  HADDX1 desc1825(.A0(N395),.B0(\add_105_I11_L14036_C191/carry[2] ),.C1(\add_105_I11_L14036_C191/carry[3] ),.SO(N406));
  HADDX1 desc1826(.A0(N396),.B0(\add_105_I11_L14036_C191/carry[3] ),.C1(\add_105_I11_L14036_C191/carry[4] ),.SO(N407));
  HADDX1 desc1827(.A0(N397),.B0(\add_105_I11_L14036_C191/carry[4] ),.C1(\add_105_I11_L14036_C191/carry[5] ),.SO(N408));
  HADDX1 desc1828(.A0(N377),.B0(N376),.C1(\add_105_I10_L14036_C191/carry[2] ),.SO(N388));
  HADDX1 desc1829(.A0(N378),.B0(\add_105_I10_L14036_C191/carry[2] ),.C1(\add_105_I10_L14036_C191/carry[3] ),.SO(N389));
  HADDX1 desc1830(.A0(N379),.B0(\add_105_I10_L14036_C191/carry[3] ),.C1(\add_105_I10_L14036_C191/carry[4] ),.SO(N390));
  HADDX1 desc1831(.A0(N380),.B0(\add_105_I10_L14036_C191/carry[4] ),.C1(\add_105_I10_L14036_C191/carry[5] ),.SO(N391));
  HADDX1 desc1832(.A0(N360),.B0(N359),.C1(\add_105_I9_L14036_C191/carry[2] ),.SO(N371));
  HADDX1 desc1833(.A0(N361),.B0(\add_105_I9_L14036_C191/carry[2] ),.C1(\add_105_I9_L14036_C191/carry[3] ),.SO(N372));
  HADDX1 desc1834(.A0(N362),.B0(\add_105_I9_L14036_C191/carry[3] ),.C1(\add_105_I9_L14036_C191/carry[4] ),.SO(N373));
  HADDX1 desc1835(.A0(N363),.B0(\add_105_I9_L14036_C191/carry[4] ),.C1(\add_105_I9_L14036_C191/carry[5] ),.SO(N374));
  HADDX1 desc1836(.A0(N343),.B0(N342),.C1(\add_105_I8_L14036_C191/carry[2] ),.SO(N354));
  HADDX1 desc1837(.A0(N344),.B0(\add_105_I8_L14036_C191/carry[2] ),.C1(\add_105_I8_L14036_C191/carry[3] ),.SO(N355));
  HADDX1 desc1838(.A0(N345),.B0(\add_105_I8_L14036_C191/carry[3] ),.C1(\add_105_I8_L14036_C191/carry[4] ),.SO(N356));
  HADDX1 desc1839(.A0(N346),.B0(\add_105_I8_L14036_C191/carry[4] ),.C1(\add_105_I8_L14036_C191/carry[5] ),.SO(N357));
  HADDX1 desc1840(.A0(N326),.B0(N325),.C1(\add_105_I7_L14036_C191/carry[2] ),.SO(N337));
  HADDX1 desc1841(.A0(N327),.B0(\add_105_I7_L14036_C191/carry[2] ),.C1(\add_105_I7_L14036_C191/carry[3] ),.SO(N338));
  HADDX1 desc1842(.A0(N328),.B0(\add_105_I7_L14036_C191/carry[3] ),.C1(\add_105_I7_L14036_C191/carry[4] ),.SO(N339));
  HADDX1 desc1843(.A0(N329),.B0(\add_105_I7_L14036_C191/carry[4] ),.C1(N341),.SO(N340));
  HADDX1 desc1844(.A0(N310),.B0(N309),.C1(\add_105_I6_L14036_C191/carry[2] ),.SO(N320));
  HADDX1 desc1845(.A0(N311),.B0(\add_105_I6_L14036_C191/carry[2] ),.C1(\add_105_I6_L14036_C191/carry[3] ),.SO(N321));
  HADDX1 desc1846(.A0(N312),.B0(\add_105_I6_L14036_C191/carry[3] ),.C1(N323),.SO(N322));
  HADDX1 desc1847(.A0(\add_105_I5_L14036_C191/A[1] ),.B0(N295),.C1(\add_105_I5_L14036_C191/carry[2] ),.SO(N305));
  HADDX1 desc1848(.A0(N297),.B0(\add_105_I5_L14036_C191/carry[2] ),.C1(N307),.SO(N306));
  p_O_DFFX1 desc1849(.D(N175),.CLK(clk_i),.Q(s_shr1[3:3]),.QN(n3),.E(p_desc1849_p_O_DFFX1));
  p_O_DFFX1 desc1850(.D(qutnt_i[25:25]),.CLK(clk_i),.Q(s_qutnt_i[25:25]),.QN(n60),.E(p_desc1850_p_O_DFFX1));
  p_O_DFFX1 desc1851(.D(qutnt_i[23:23]),.CLK(clk_i),.Q(s_qutnt_i[23:23]),.QN(n62),.E(p_desc1851_p_O_DFFX1));
  p_O_DFFX1 desc1852(.D(qutnt_i[24:24]),.CLK(clk_i),.Q(s_qutnt_i[24:24]),.QN(n61),.E(p_desc1852_p_O_DFFX1));
  p_O_DFFX1 desc1853(.D(qutnt_i[22:22]),.CLK(clk_i),.Q(s_qutnt_i[22:22]),.QN(n63),.E(p_desc1853_p_O_DFFX1));
  p_O_DFFX1 desc1854(.D(qutnt_i[21:21]),.CLK(clk_i),.Q(s_qutnt_i[21:21]),.QN(n64),.E(p_desc1854_p_O_DFFX1));
  p_O_DFFX1 desc1855(.D(qutnt_i[20:20]),.CLK(clk_i),.Q(s_qutnt_i[20:20]),.QN(n71),.E(p_desc1855_p_O_DFFX1));
  p_O_DFFX1 desc1856(.D(qutnt_i[19:19]),.CLK(clk_i),.Q(s_qutnt_i[19:19]),.QN(n79),.E(p_desc1856_p_O_DFFX1));
  p_O_DFFX1 desc1857(.D(qutnt_i[18:18]),.CLK(clk_i),.Q(s_qutnt_i[18:18]),.QN(n86),.E(p_desc1857_p_O_DFFX1));
  p_O_DFFX1 desc1858(.D(qutnt_i[17:17]),.CLK(clk_i),.Q(s_qutnt_i[17:17]),.QN(n93),.E(p_desc1858_p_O_DFFX1));
  p_O_DFFX1 desc1859(.D(qutnt_i[16:16]),.CLK(clk_i),.Q(s_qutnt_i[16:16]),.QN(n94),.E(p_desc1859_p_O_DFFX1));
  p_O_DFFX1 desc1860(.D(qutnt_i[14:14]),.CLK(clk_i),.Q(s_qutnt_i[14:14]),.QN(n96),.E(p_desc1860_p_O_DFFX1));
  p_O_DFFX1 desc1861(.D(qutnt_i[15:15]),.CLK(clk_i),.Q(s_qutnt_i[15:15]),.QN(n95),.E(p_desc1861_p_O_DFFX1));
  p_O_DFFX1 desc1862(.D(qutnt_i[11:11]),.CLK(clk_i),.Q(s_qutnt_i[11:11]),.QN(n99),.E(p_desc1862_p_O_DFFX1));
  p_O_DFFX1 desc1863(.D(qutnt_i[13:13]),.CLK(clk_i),.Q(s_qutnt_i[13:13]),.QN(n97),.E(p_desc1863_p_O_DFFX1));
  p_O_DFFX1 desc1864(.D(qutnt_i[12:12]),.CLK(clk_i),.Q(s_qutnt_i[12:12]),.QN(n98),.E(p_desc1864_p_O_DFFX1));
  p_O_DFFX1 desc1865(.D(qutnt_i[7:7]),.CLK(clk_i),.Q(s_qutnt_i[7:7]),.QN(n104),.E(p_desc1865_p_O_DFFX1));
  p_O_DFFX1 desc1866(.D(qutnt_i[10:10]),.CLK(clk_i),.Q(s_qutnt_i[10:10]),.QN(n100),.E(p_desc1866_p_O_DFFX1));
  p_O_DFFX1 desc1867(.D(qutnt_i[8:8]),.CLK(clk_i),.Q(s_qutnt_i[8:8]),.QN(n103),.E(p_desc1867_p_O_DFFX1));
  p_O_DFFX1 desc1868(.D(qutnt_i[9:9]),.CLK(clk_i),.Q(s_qutnt_i[9:9]),.QN(n101),.E(p_desc1868_p_O_DFFX1));
  p_O_DFFX1 desc1869(.D(qutnt_i[6:6]),.CLK(clk_i),.Q(s_qutnt_i[6:6]),.QN(n105),.E(p_desc1869_p_O_DFFX1));
  OA21X1 U3(.IN1(s_sign_i),.IN2(n305),.IN3(n306),.Q(n301));
  XOR2X1 U4(.IN1(s_qutnt_i[26:26]),.IN2(s_exp_10_i[0:0]),.Q(n1));
  NAND2X1 U5(.IN1(n159),.IN2(N326),.QN(n201));
  NBUFFX2 U6(.INP(\add_194/B[0] ),.Z(n15));
  NBUFFX2 U7(.INP(\add_194/B[0] ),.Z(n16));
  NOR2X0 U14(.IN1(n72),.IN2(n73),.QN(n14));
  NOR2X0 U15(.IN1(n72),.IN2(n73),.QN(n245));
  INVX0 U16(.INP(n203),.ZN(\add_105_I5_L14036_C191/A[1] ));
  NOR2X0 U17(.IN1(n21),.IN2(n15),.QN(n298));
  INVX0 U18(.INP(n300),.ZN(\add_194/B[0] ));
  INVX0 U19(.INP(n249),.ZN(n73));
  INVX0 U20(.INP(n247),.ZN(n72));
  INVX0 U21(.INP(n377),.ZN(n77));
  NOR2X0 U22(.IN1(n268),.IN2(n72),.QN(N1386));
  INVX0 U23(.INP(N532),.ZN(n116));
  INVX0 U24(.INP(N583),.ZN(n85));
  NOR2X0 U25(.IN1(n181),.IN2(n182),.QN(n180));
  INVX0 U26(.INP(N531),.ZN(n120));
  INVX0 U27(.INP(N582),.ZN(n87));
  NOR2X0 U28(.IN1(n195),.IN2(n196),.QN(n194));
  INVX0 U29(.INP(N534),.ZN(n66));
  INVX0 U30(.INP(N585),.ZN(n58));
  NOR2X0 U31(.IN1(n146),.IN2(n147),.QN(n144));
  INVX0 U32(.INP(N533),.ZN(n70));
  INVX0 U33(.INP(N584),.ZN(n67));
  NOR2X0 U34(.IN1(n169),.IN2(n170),.QN(n168));
  AOI221X1 U35(.IN1(n126),.IN2(N381),.IN3(n127),.IN4(n128),.IN5(n129),.QN(n7));
  NAND2X1 U36(.IN1(n183),.IN2(n184),.QN(s_r_zeros[2:2]));
  AOI221X1 U37(.IN1(n127),.IN2(n171),.IN3(n159),.IN4(N328),.IN5(n172),.QN(n8));
  AOI221X1 U39(.IN1(n127),.IN2(n158),.IN3(n159),.IN4(N329),.IN5(n160),.QN(n9));
  AOI22X1 U40(.IN1(n328),.IN2(n198),.IN3(n199),.IN4(n200),.QN(n10));
  INVX0 U41(.INP(N547),.ZN(n114));
  INVX0 U42(.INP(N549),.ZN(n110));
  INVX0 U43(.INP(N548),.ZN(n111));
  INVX0 U44(.INP(N550),.ZN(n69));
  INVX0 U45(.INP(N551),.ZN(n65));
  INVX0 U46(.INP(N564),.ZN(n107));
  INVX0 U47(.INP(N566),.ZN(n92));
  INVX0 U48(.INP(N565),.ZN(n102));
  INVX0 U49(.INP(N567),.ZN(n68));
  INVX0 U50(.INP(N568),.ZN(n59));
  INVX0 U51(.INP(N581),.ZN(n88));
  INVX0 U52(.INP(N580),.ZN(n89));
  INVX0 U53(.INP(N530),.ZN(n121));
  NAND2X1 U54(.IN1(N1089),.IN2(n13),.QN(n300));
  INVX0 U55(.INP(N1021),.ZN(n51));
  NOR2X0 U56(.IN1(n238),.IN2(n239),.QN(n150));
  NOR2X0 U57(.IN1(n229),.IN2(n137),.QN(n136));
  NOR2X0 U58(.IN1(n221),.IN2(n127),.QN(n126));
  INVX0 U59(.INP(n240),.ZN(n75));
  INVX0 U60(.INP(n241),.ZN(n91));
  NAND2X1 U61(.IN1(n91),.IN2(n145),.QN(n143));
  INVX0 U62(.INP(n127),.ZN(n321));
  INVX0 U63(.INP(n185),.ZN(n327));
  INVX0 U64(.INP(n13),.ZN(n21));
  INVX0 U65(.INP(n264),.ZN(n52));
  NOR2X0 U66(.IN1(n222),.IN2(n220),.QN(n131));
  XOR2X1 U67(.IN1(s_exp_10b[6:6]),.IN2(n11),.Q(N151));
  NAND2X1 U68(.IN1(\sub_1_root_sub_150_2/carry[5] ),.IN2(n33),.QN(n11));
  NOR2X0 U69(.IN1(n227),.IN2(n228),.QN(n156));
  INVX0 U70(.INP(s_exp_10b[6:6]),.ZN(n55));
  INVX0 U71(.INP(s_exp_10b[7:7]),.ZN(n54));
  NAND2X1 U72(.IN1(n242),.IN2(n243),.QN(n142));
  NAND2X1 U73(.IN1(n244),.IN2(n241),.QN(n154));
  NAND2X1 U74(.IN1(n159),.IN2(N325),.QN(n217));
  NAND2X1 U75(.IN1(n264),.IN2(n1),.QN(N162));
  INVX0 U76(.INP(n279),.ZN(n329));
  INVX0 U77(.INP(s_exp_10b[8:8]),.ZN(n53));
  INVX0 U78(.INP(n261),.ZN(n24));
  INVX0 U79(.INP(n261),.ZN(n23));
  NBUFFX2 U80(.INP(n6),.Z(n20));
  NOR2X0 U81(.IN1(n255),.IN2(n254),.QN(n247));
  NBUFFX2 U82(.INP(n5),.Z(n18));
  NAND2X1 U83(.IN1(n368),.IN2(n2),.QN(n388));
  NAND2X1 U84(.IN1(n377),.IN2(n3),.QN(n409));
  NAND2X1 U85(.IN1(n390),.IN2(n3),.QN(n446));
  NAND2X1 U86(.IN1(n375),.IN2(n3),.QN(n391));
  INVX0 U87(.INP(s_exp_10b[2:2]),.ZN(n57));
  INVX0 U88(.INP(s_exp_10b[3:3]),.ZN(n56));
  NAND2X1 U89(.IN1(n352),.IN2(n17),.QN(n374));
  INVX0 U90(.INP(n390),.ZN(n78));
  INVX0 U91(.INP(n375),.ZN(n76));
  INVX0 U92(.INP(n369),.ZN(n115));
  INVX0 U93(.INP(n381),.ZN(n318));
  INVX0 U94(.INP(n371),.ZN(n83));
  INVX0 U95(.INP(n257),.ZN(n74));
  INVX0 U96(.INP(n392),.ZN(n324));
  INVX0 U97(.INP(n359),.ZN(n316));
  INVX0 U98(.INP(n402),.ZN(n320));
  INVX0 U99(.INP(n396),.ZN(n326));
  INVX0 U100(.INP(n406),.ZN(n325));
  INVX0 U101(.INP(n412),.ZN(n323));
  INVX0 U102(.INP(n419),.ZN(n319));
  INVX0 U103(.INP(s_exp_10b[1:1]),.ZN(n31));
  INVX0 U104(.INP(s_exp_10b[4:4]),.ZN(n32));
  INVX0 U105(.INP(s_exp_10b[5:5]),.ZN(n33));
  INVX0 U106(.INP(n361),.ZN(n299));
  INVX0 U107(.INP(n355),.ZN(n81));
  INVX0 U108(.INP(n358),.ZN(n90));
  INVX0 U109(.INP(n200),.ZN(n328));
  INVX0 U110(.INP(N309),.ZN(N319));
  INVX0 U111(.INP(N342),.ZN(N353));
  INVX0 U112(.INP(N393),.ZN(N404));
  INVX0 U113(.INP(N359),.ZN(N370));
  INVX0 U114(.INP(N376),.ZN(N387));
  INVX0 U115(.INP(N444),.ZN(N455));
  INVX0 U116(.INP(N427),.ZN(N438));
  INVX0 U117(.INP(N410),.ZN(N421));
  NOR2X0 U118(.IN1(s_qutnt_i[0:0]),.IN2(s_qutnt_i[1:1]),.QN(n199));
  NOR2X0 U119(.IN1(n213),.IN2(n214),.QN(n212));
  INVX0 U120(.INP(N295),.ZN(N304));
  NOR2X0 U121(.IN1(n260),.IN2(s_qutnt_i[3:3]),.QN(n258));
  AND2X1 U122(.IN1(N341),.IN2(n105),.Q(n12));
  INVX0 U123(.INP(N325),.ZN(N336));
  INVX0 U124(.INP(N512),.ZN(N523));
  INVX0 U125(.INP(N529),.ZN(N540));
  INVX0 U126(.INP(N546),.ZN(N557));
  INVX0 U127(.INP(N563),.ZN(N574));
  INVX0 U139(.INP(N631),.ZN(N642));
  INVX0 U151(.INP(N614),.ZN(N625));
  INVX0 U175(.INP(N495),.ZN(N506));
  INVX0 U349(.INP(N597),.ZN(N608));
  INVX0 U355(.INP(N478),.ZN(N489));
  INVX0 U356(.INP(N648),.ZN(N659));
  INVX0 U361(.INP(N461),.ZN(N472));
  NOR2X0 U366(.IN1(n235),.IN2(n236),.QN(n234));
  INVX0 U493(.INP(N665),.ZN(N676));
  NOR2X0 U494(.IN1(s_qutnt_i[15:15]),.IN2(s_qutnt_i[16:16]),.QN(n242));
  NOR2X0 U495(.IN1(n229),.IN2(s_qutnt_i[14:14]),.QN(n137));
  NOR2X0 U496(.IN1(n221),.IN2(s_qutnt_i[8:8]),.QN(n127));
  NOR2X0 U497(.IN1(s_qutnt_i[21:21]),.IN2(s_qutnt_i[22:22]),.QN(n237));
  NOR2X0 U498(.IN1(n243),.IN2(s_qutnt_i[18:18]),.QN(n244));
  NOR2X0 U499(.IN1(s_qutnt_i[10:10]),.IN2(s_qutnt_i[9:9]),.QN(n226));
  NOR2X0 U500(.IN1(n227),.IN2(s_qutnt_i[12:12]),.QN(n228));
  NOR2X0 U501(.IN1(n222),.IN2(s_qutnt_i[6:6]),.QN(n220));
  NAND2X1 U502(.IN1(n91),.IN2(n71),.QN(n145));
  NAND2X1 U503(.IN1(n242),.IN2(n93),.QN(n243));
  NAND2X1 U504(.IN1(n327),.IN2(n106),.QN(n222));
  NAND2X1 U505(.IN1(n237),.IN2(n62),.QN(n238));
  NAND2X1 U506(.IN1(n226),.IN2(n99),.QN(n227));
  NAND2X1 U507(.IN1(n228),.IN2(n97),.QN(n229));
  NAND2X1 U508(.IN1(n220),.IN2(n104),.QN(n221));
  NOR2X0 U509(.IN1(n238),.IN2(s_qutnt_i[24:24]),.QN(n239));
  NOR2X0 U510(.IN1(n200),.IN2(s_qutnt_i[3:3]),.QN(n186));
  NAND2X1 U511(.IN1(n199),.IN2(n112),.QN(n200));
  NAND2X1 U512(.IN1(n244),.IN2(n79),.QN(n241));
  NAND2X1 U513(.IN1(n186),.IN2(n108),.QN(n185));
  NOR2X0 U514(.IN1(n265),.IN2(s_exp_10b[9:9]),.QN(n264));
  OAI21X1 U515(.IN1(n329),.IN2(n301),.IN3(n302),.QN(n13));
  NOR2X0 U516(.IN1(n237),.IN2(s_qutnt_i[21:21]),.QN(n148));
  NOR2X0 U517(.IN1(n226),.IN2(s_qutnt_i[9:9]),.QN(n155));
  NOR2X0 U518(.IN1(n242),.IN2(s_qutnt_i[15:15]),.QN(n152));
  NAND2X1 U519(.IN1(\s_rmode_i[1] ),.IN2(n119),.QN(n305));
  NBUFFX2 U520(.INP(s_shr1[5:5]),.Z(n29));
  NOR2X0 U521(.IN1(n286),.IN2(n287),.QN(n285));
  NOR2X0 U522(.IN1(n374),.IN2(s_shr1[2:2]),.QN(n390));
  NOR2X0 U523(.IN1(n364),.IN2(s_shr1[2:2]),.QN(n375));
  NOR2X0 U524(.IN1(n281),.IN2(n282),.QN(n250));
  NOR2X0 U525(.IN1(n283),.IN2(n284),.QN(n252));
  NAND2X1 U526(.IN1(s_qutnt_i[26:26]),.IN2(n19),.QN(n343));
  NOR2X0 U527(.IN1(n29),.IN2(n425),.QN(N189));
  INVX0 U528(.INP(n332),.ZN(n322));
  NAND2X1 U529(.IN1(n246),.IN2(n248),.QN(s_output_o[22:22]));
  NOR2X0 U530(.IN1(n29),.IN2(n401),.QN(N186));
  NOR2X0 U531(.IN1(n29),.IN2(n411),.QN(N187));
  NOR2X0 U532(.IN1(n29),.IN2(n418),.QN(N188));
  NOR2X0 U533(.IN1(n29),.IN2(n432),.QN(N190));
  NOR2X0 U534(.IN1(n29),.IN2(n438),.QN(N191));
  NOR2X0 U535(.IN1(n29),.IN2(n443),.QN(N192));
  NOR2X0 U536(.IN1(n29),.IN2(n448),.QN(N193));
  NOR2X0 U537(.IN1(n29),.IN2(n345),.QN(N194));
  NOR2X0 U538(.IN1(n29),.IN2(n384),.QN(N185));
  NOR2X0 U539(.IN1(n25),.IN2(n113),.QN(N211));
  NOR2X0 U540(.IN1(n341),.IN2(n29),.QN(N184));
  NAND2X1 U541(.IN1(n246),.IN2(n117),.QN(s_output_o[31:31]));
  INVX0 U542(.INP(n337),.ZN(n84));
  INVX0 U543(.INP(n334),.ZN(n317));
  INVX0 U544(.INP(n338),.ZN(n109));
  INVX0 U545(.INP(n336),.ZN(n82));
  INVX0 U546(.INP(n335),.ZN(n80));
  INVX0 U547(.INP(n339),.ZN(n125));
  INVX0 U548(.INP(n333),.ZN(n315));
  NBUFFX2 U549(.INP(s_shr1[4:4]),.Z(n28));
  NBUFFX2 U550(.INP(s_shr1[5:5]),.Z(n30));
  NBUFFX2 U551(.INP(\s_shl1[0] ),.Z(n26));
  NBUFFX4 U552(.INP(n5),.Z(n17));
  NBUFFX4 U553(.INP(n6),.Z(n19));
  NBUFFX4 U554(.INP(\s_shl1[0] ),.Z(n25));
  NBUFFX4 U555(.INP(s_shr1[4:4]),.Z(n27));
  INVX0 U556(.INP(n24),.ZN(n22));
  XOR2X1 U557(.IN1(n29),.IN2(\add_194/carry[5] ),.Q(N1024));
  AND2X1 U558(.IN1(\add_194/carry[4] ),.IN2(s_shr1[4:4]),.Q(\add_194/carry[5] ));
  XOR2X1 U559(.IN1(n27),.IN2(\add_194/carry[4] ),.Q(N1023));
  AND2X1 U560(.IN1(\add_194/carry[3] ),.IN2(s_shr1[3:3]),.Q(\add_194/carry[4] ));
  XOR2X1 U561(.IN1(s_shr1[3:3]),.IN2(\add_194/carry[3] ),.Q(N1022));
  AND2X1 U562(.IN1(\add_194/carry[2] ),.IN2(s_shr1[2:2]),.Q(\add_194/carry[3] ));
  XOR2X1 U563(.IN1(s_shr1[2:2]),.IN2(\add_194/carry[2] ),.Q(N1021));
  AND2X1 U564(.IN1(\add_194/carry[1] ),.IN2(s_shr1[1:1]),.Q(\add_194/carry[2] ));
  XOR2X1 U565(.IN1(s_shr1[1:1]),.IN2(\add_194/carry[1] ),.Q(N1020));
  AND2X1 U566(.IN1(n16),.IN2(s_shr1[0:0]),.Q(\add_194/carry[1] ));
  XOR2X1 U567(.IN1(s_shr1[0:0]),.IN2(n15),.Q(N1019));
  XNOR2X1 U568(.IN1(s_expo1[8:8]),.IN2(\sub_188_aco/carry[8] ),.Q(s_expo2[8:8]));
  OR2X1 U569(.IN1(s_expo1[7:7]),.IN2(\sub_188_aco/carry[7] ),.Q(\sub_188_aco/carry[8] ));
  XNOR2X1 U570(.IN1(\sub_188_aco/carry[7] ),.IN2(s_expo1[7:7]),.Q(s_expo2[7:7]));
  OR2X1 U571(.IN1(s_expo1[6:6]),.IN2(\sub_188_aco/carry[6] ),.Q(\sub_188_aco/carry[7] ));
  XNOR2X1 U572(.IN1(\sub_188_aco/carry[6] ),.IN2(s_expo1[6:6]),.Q(s_expo2[6:6]));
  OR2X1 U573(.IN1(s_expo1[5:5]),.IN2(\sub_188_aco/carry[5] ),.Q(\sub_188_aco/carry[6] ));
  XNOR2X1 U574(.IN1(\sub_188_aco/carry[5] ),.IN2(s_expo1[5:5]),.Q(s_expo2[5:5]));
  OR2X1 U575(.IN1(s_expo1[4:4]),.IN2(\sub_188_aco/carry[4] ),.Q(\sub_188_aco/carry[5] ));
  XNOR2X1 U576(.IN1(\sub_188_aco/carry[4] ),.IN2(s_expo1[4:4]),.Q(s_expo2[4:4]));
  OR2X1 U577(.IN1(s_expo1[3:3]),.IN2(\sub_188_aco/carry[3] ),.Q(\sub_188_aco/carry[4] ));
  XNOR2X1 U578(.IN1(\sub_188_aco/carry[3] ),.IN2(s_expo1[3:3]),.Q(s_expo2[3:3]));
  OR2X1 U579(.IN1(s_expo1[2:2]),.IN2(\sub_188_aco/carry[2] ),.Q(\sub_188_aco/carry[3] ));
  XNOR2X1 U580(.IN1(\sub_188_aco/carry[2] ),.IN2(s_expo1[2:2]),.Q(s_expo2[2:2]));
  OR2X1 U581(.IN1(s_expo1[1:1]),.IN2(\sub_188_aco/carry[1] ),.Q(\sub_188_aco/carry[2] ));
  XNOR2X1 U582(.IN1(\sub_188_aco/carry[1] ),.IN2(s_expo1[1:1]),.Q(s_expo2[1:1]));
  OR2X1 U583(.IN1(s_expo1[0:0]),.IN2(s_fraco1[26:26]),.Q(\sub_188_aco/carry[1] ));
  XNOR2X1 U584(.IN1(s_fraco1[26:26]),.IN2(s_expo1[0:0]),.Q(s_expo2[0:0]));
  XOR2X1 U585(.IN1(n33),.IN2(\sub_1_root_sub_150_2/carry[5] ),.Q(N150));
  AND2X1 U586(.IN1(\sub_1_root_sub_150_2/carry[4] ),.IN2(n32),.Q(\sub_1_root_sub_150_2/carry[5] ));
  XOR2X1 U587(.IN1(n32),.IN2(\sub_1_root_sub_150_2/carry[4] ),.Q(N149));
  AND2X1 U588(.IN1(\sub_1_root_sub_150_2/carry[3] ),.IN2(n56),.Q(\sub_1_root_sub_150_2/carry[4] ));
  XOR2X1 U589(.IN1(n56),.IN2(\sub_1_root_sub_150_2/carry[3] ),.Q(N148));
  AND2X1 U590(.IN1(\sub_1_root_sub_150_2/carry[2] ),.IN2(n57),.Q(\sub_1_root_sub_150_2/carry[3] ));
  XOR2X1 U591(.IN1(n57),.IN2(\sub_1_root_sub_150_2/carry[2] ),.Q(N147));
  AND2X1 U592(.IN1(\sub_1_root_sub_150_2/carry[1] ),.IN2(n31),.Q(\sub_1_root_sub_150_2/carry[2] ));
  XOR2X1 U593(.IN1(n31),.IN2(\sub_1_root_sub_150_2/carry[1] ),.Q(N146));
  OR2X1 U594(.IN1(n1),.IN2(s_qutnt_i[26:26]),.Q(\sub_1_root_sub_150_2/carry[1] ));
  XNOR2X1 U595(.IN1(s_qutnt_i[26:26]),.IN2(n1),.Q(N145));
  XNOR2X1 U596(.IN1(s_exp_10_i[9:9]),.IN2(\sub_141/carry[9] ),.Q(s_exp_10b[9:9]));
  OR2X1 U597(.IN1(s_exp_10_i[8:8]),.IN2(\sub_141/carry[8] ),.Q(\sub_141/carry[9] ));
  XNOR2X1 U598(.IN1(\sub_141/carry[8] ),.IN2(s_exp_10_i[8:8]),.Q(s_exp_10b[8:8]));
  OR2X1 U599(.IN1(s_exp_10_i[7:7]),.IN2(\sub_141/carry[7] ),.Q(\sub_141/carry[8] ));
  XNOR2X1 U600(.IN1(\sub_141/carry[7] ),.IN2(s_exp_10_i[7:7]),.Q(s_exp_10b[7:7]));
  OR2X1 U601(.IN1(s_exp_10_i[6:6]),.IN2(\sub_141/carry[6] ),.Q(\sub_141/carry[7] ));
  XNOR2X1 U602(.IN1(\sub_141/carry[6] ),.IN2(s_exp_10_i[6:6]),.Q(s_exp_10b[6:6]));
  OR2X1 U603(.IN1(s_exp_10_i[5:5]),.IN2(\sub_141/carry[5] ),.Q(\sub_141/carry[6] ));
  XNOR2X1 U604(.IN1(\sub_141/carry[5] ),.IN2(s_exp_10_i[5:5]),.Q(s_exp_10b[5:5]));
  OR2X1 U605(.IN1(s_exp_10_i[4:4]),.IN2(\sub_141/carry[4] ),.Q(\sub_141/carry[5] ));
  XNOR2X1 U606(.IN1(\sub_141/carry[4] ),.IN2(s_exp_10_i[4:4]),.Q(s_exp_10b[4:4]));
  OR2X1 U607(.IN1(s_exp_10_i[3:3]),.IN2(\sub_141/carry[3] ),.Q(\sub_141/carry[4] ));
  XNOR2X1 U608(.IN1(\sub_141/carry[3] ),.IN2(s_exp_10_i[3:3]),.Q(s_exp_10b[3:3]));
  OR2X1 U609(.IN1(s_exp_10_i[2:2]),.IN2(\sub_141/carry[2] ),.Q(\sub_141/carry[3] ));
  XNOR2X1 U610(.IN1(\sub_141/carry[2] ),.IN2(s_exp_10_i[2:2]),.Q(s_exp_10b[2:2]));
  OR2X1 U611(.IN1(s_exp_10_i[1:1]),.IN2(\sub_141/carry[1] ),.Q(\sub_141/carry[2] ));
  XNOR2X1 U612(.IN1(\sub_141/carry[1] ),.IN2(s_exp_10_i[1:1]),.Q(s_exp_10b[1:1]));
  OR2X1 U613(.IN1(s_exp_10_i[0:0]),.IN2(s_qutnt_i[26:26]),.Q(\sub_141/carry[1] ));
  XOR2X1 U614(.IN1(\add_105_I8_L14036_C191/carry[5] ),.IN2(n12),.Q(N358));
  XOR2X1 U615(.IN1(\add_105_I9_L14036_C191/carry[5] ),.IN2(N364),.Q(N375));
  XOR2X1 U616(.IN1(\add_105_I10_L14036_C191/carry[5] ),.IN2(N381),.Q(N392));
  XOR2X1 U617(.IN1(\add_105_I11_L14036_C191/carry[5] ),.IN2(N398),.Q(N409));
  XOR2X1 U618(.IN1(\add_105_I12_L14036_C191/carry[5] ),.IN2(N415),.Q(N426));
  XOR2X1 U619(.IN1(\add_105_I13_L14036_C191/carry[5] ),.IN2(N432),.Q(N443));
  XOR2X1 U620(.IN1(\add_105_I14_L14036_C191/carry[5] ),.IN2(N449),.Q(N460));
  XOR2X1 U621(.IN1(\add_105_I15_L14036_C191/carry[5] ),.IN2(N466),.Q(N477));
  XOR2X1 U622(.IN1(\add_105_I16_L14036_C191/carry[5] ),.IN2(N483),.Q(N494));
  XOR2X1 U623(.IN1(\add_105_I17_L14036_C191/carry[5] ),.IN2(N500),.Q(N511));
  XOR2X1 U624(.IN1(\add_105_I18_L14036_C191/carry[5] ),.IN2(N517),.Q(N528));
  XOR2X1 U625(.IN1(\add_105_I19_L14036_C191/carry[5] ),.IN2(N534),.Q(N545));
  XOR2X1 U626(.IN1(\add_105_I20_L14036_C191/carry[5] ),.IN2(N551),.Q(N562));
  XOR2X1 U627(.IN1(\add_105_I21_L14036_C191/carry[5] ),.IN2(N568),.Q(N579));
  XOR2X1 U628(.IN1(\add_105_I22_L14036_C191/carry[5] ),.IN2(N585),.Q(N596));
  XOR2X1 U629(.IN1(\add_105_I23_L14036_C191/carry[5] ),.IN2(N602),.Q(N613));
  XOR2X1 U630(.IN1(\add_105_I24_L14036_C191/carry[5] ),.IN2(N619),.Q(N630));
  XOR2X1 U631(.IN1(\add_105_I25_L14036_C191/carry[5] ),.IN2(N636),.Q(N647));
  XOR2X1 U632(.IN1(\add_105_I26_L14036_C191/carry[5] ),.IN2(N653),.Q(N664));
  XOR2X1 U633(.IN1(\add_105_I27_L14036_C191/carry[5] ),.IN2(N670),.Q(N681));
  AO22X1 U634(.IN1(N1024),.IN2(n7),.IN3(N1023),.IN4(n9),.Q(n50));
  OR2X1 U635(.IN1(n7),.IN2(N1024),.Q(n49));
  NOR2X0 U636(.IN1(n8),.IN2(N1022),.QN(n34));
  AOI21X1 U637(.IN1(n51),.IN2(s_r_zeros[2:2]),.IN3(n34),.QN(n40));
  NOR2X0 U638(.IN1(s_r_zeros[2:2]),.IN2(n34),.QN(n35));
  AO22X1 U639(.IN1(N1022),.IN2(n8),.IN3(n35),.IN4(N1021),.Q(n39));
  NOR2X0 U640(.IN1(N1020),.IN2(n10),.QN(n36));
  NOR2X0 U641(.IN1(s_r_zeros[0:0]),.IN2(n36),.QN(n37));
  AO221X1 U642(.IN1(N1020),.IN2(n10),.IN3(n37),.IN4(N1019),.IN5(n39),.Q(n38));
  OA21X1 U643(.IN1(n40),.IN2(n39),.IN3(n38),.Q(n48));
  OA21X1 U644(.IN1(N1023),.IN2(n9),.IN3(n49),.Q(n47));
  AO22X1 U645(.IN1(n50),.IN2(n49),.IN3(n48),.IN4(n47),.Q(N1025));
  AND2X1 U646(.IN1(N323),.IN2(n106),.Q(N329));
  MUX21X1 U647(.IN1(s_qutnt_i[3:3]),.IN2(s_qutnt_i[2:2]),.S(n20),.Q(n394));
  MUX21X1 U648(.IN1(s_qutnt_i[1:1]),.IN2(s_qutnt_i[0:0]),.S(n20),.Q(n330));
  MUX21X1 U649(.IN1(n394),.IN2(n330),.S(n18),.Q(n331));
  MUX21X1 U650(.IN1(s_qutnt_i[7:7]),.IN2(s_qutnt_i[6:6]),.S(n20),.Q(n392));
  MUX21X1 U651(.IN1(s_qutnt_i[5:5]),.IN2(s_qutnt_i[4:4]),.S(n20),.Q(n395));
  MUX21X1 U652(.IN1(n392),.IN2(n395),.S(n18),.Q(n412));
  MUX21X1 U653(.IN1(n331),.IN2(n412),.S(s_shr1[2:2]),.Q(n332));
  MUX21X1 U654(.IN1(s_qutnt_i[15:15]),.IN2(s_qutnt_i[14:14]),.S(n20),.Q(n333));
  MUX21X1 U655(.IN1(s_qutnt_i[13:13]),.IN2(s_qutnt_i[12:12]),.S(n20),.Q(n334));
  MUX21X1 U656(.IN1(n315),.IN2(n317),.S(n18),.Q(n349));
  MUX21X1 U657(.IN1(n99),.IN2(n100),.S(n20),.Q(n342));
  MUX21X1 U658(.IN1(n101),.IN2(n103),.S(n20),.Q(n393));
  MUX21X1 U659(.IN1(n342),.IN2(n393),.S(n18),.Q(n413));
  MUX21X1 U660(.IN1(n349),.IN2(n413),.S(n2),.Q(n439));
  MUX21X1 U661(.IN1(n322),.IN2(n439),.S(s_shr1[3:3]),.Q(n340));
  MUX21X1 U662(.IN1(s_qutnt_i[25:25]),.IN2(s_qutnt_i[24:24]),.S(n20),.Q(n335));
  MUX21X1 U663(.IN1(n343),.IN2(n80),.S(n18),.Q(n348));
  OR2X1 U664(.IN1(n348),.IN2(s_shr1[2:2]),.Q(n389));
  MUX21X1 U665(.IN1(s_qutnt_i[23:23]),.IN2(s_qutnt_i[22:22]),.S(n20),.Q(n336));
  MUX21X1 U666(.IN1(s_qutnt_i[21:21]),.IN2(s_qutnt_i[20:20]),.S(n19),.Q(n337));
  MUX21X1 U667(.IN1(n82),.IN2(n84),.S(n18),.Q(n347));
  MUX21X1 U668(.IN1(s_qutnt_i[19:19]),.IN2(s_qutnt_i[18:18]),.S(n19),.Q(n338));
  MUX21X1 U669(.IN1(s_qutnt_i[17:17]),.IN2(s_qutnt_i[16:16]),.S(n19),.Q(n339));
  MUX21X1 U670(.IN1(n109),.IN2(n125),.S(n18),.Q(n350));
  MUX21X1 U671(.IN1(n347),.IN2(n350),.S(n2),.Q(n440));
  MUX21X1 U672(.IN1(n389),.IN2(n440),.S(n3),.Q(n373));
  MUX21X1 U673(.IN1(n340),.IN2(n373),.S(n27),.Q(n341));
  MUX21X1 U674(.IN1(n80),.IN2(n82),.S(n18),.Q(n363));
  MUX21X1 U675(.IN1(n84),.IN2(n109),.S(n18),.Q(n366));
  MUX21X1 U676(.IN1(n363),.IN2(n366),.S(n2),.Q(n376));
  MUX21X1 U677(.IN1(n125),.IN2(n315),.S(n17),.Q(n365));
  MUX21X1 U678(.IN1(n317),.IN2(n342),.S(n17),.Q(n427));
  MUX21X1 U679(.IN1(n365),.IN2(n427),.S(n2),.Q(n398));
  MUX21X1 U680(.IN1(n376),.IN2(n398),.S(n3),.Q(n344));
  OR2X1 U681(.IN1(n343),.IN2(s_shr1[1:1]),.Q(n364));
  MUX21X1 U682(.IN1(n344),.IN2(n391),.S(n27),.Q(n345));
  MUX21X1 U683(.IN1(s_qutnt_i[26:26]),.IN2(s_qutnt_i[25:25]),.S(n19),.Q(n352));
  MUX21X1 U684(.IN1(s_qutnt_i[24:24]),.IN2(s_qutnt_i[23:23]),.S(n19),.Q(n354));
  MUX21X1 U685(.IN1(n352),.IN2(n354),.S(n17),.Q(n368));
  MUX21X1 U686(.IN1(s_qutnt_i[22:22]),.IN2(s_qutnt_i[21:21]),.S(n19),.Q(n353));
  MUX21X1 U687(.IN1(s_qutnt_i[20:20]),.IN2(s_qutnt_i[19:19]),.S(n19),.Q(n357));
  MUX21X1 U688(.IN1(n353),.IN2(n357),.S(n17),.Q(n370));
  MUX21X1 U689(.IN1(n368),.IN2(n370),.S(n2),.Q(n377));
  MUX21X1 U690(.IN1(s_qutnt_i[18:18]),.IN2(s_qutnt_i[17:17]),.S(n19),.Q(n356));
  MUX21X1 U691(.IN1(s_qutnt_i[16:16]),.IN2(s_qutnt_i[15:15]),.S(n19),.Q(n360));
  MUX21X1 U692(.IN1(n356),.IN2(n360),.S(n17),.Q(n369));
  MUX21X1 U693(.IN1(s_qutnt_i[14:14]),.IN2(s_qutnt_i[13:13]),.S(n19),.Q(n359));
  MUX21X1 U694(.IN1(n98),.IN2(n99),.S(n19),.Q(n378));
  MUX21X1 U695(.IN1(n316),.IN2(n378),.S(n17),.Q(n434));
  MUX21X1 U696(.IN1(n115),.IN2(n434),.S(n2),.Q(n408));
  MUX21X1 U697(.IN1(n77),.IN2(n408),.S(n3),.Q(n346));
  NOR3X0 U698(.IN1(n28),.IN2(n29),.IN3(n346),.QN(N195));
  MUX21X1 U699(.IN1(n348),.IN2(n347),.S(n2),.Q(n385));
  MUX21X1 U700(.IN1(n350),.IN2(n349),.S(n2),.Q(n415));
  MUX21X1 U701(.IN1(n385),.IN2(n415),.S(n3),.Q(n351));
  NOR3X0 U702(.IN1(n28),.IN2(n30),.IN3(n351),.QN(N196));
  MUX21X1 U703(.IN1(n354),.IN2(n353),.S(n17),.Q(n355));
  MUX21X1 U704(.IN1(n374),.IN2(n81),.S(n2),.Q(n386));
  MUX21X1 U705(.IN1(n357),.IN2(n356),.S(n17),.Q(n358));
  MUX21X1 U706(.IN1(n360),.IN2(n359),.S(n17),.Q(n361));
  MUX21X1 U707(.IN1(n90),.IN2(n299),.S(n2),.Q(n422));
  MUX21X1 U708(.IN1(n386),.IN2(n422),.S(n3),.Q(n362));
  NOR3X0 U709(.IN1(n28),.IN2(n30),.IN3(n362),.QN(N197));
  MUX21X1 U710(.IN1(n364),.IN2(n363),.S(n2),.Q(n387));
  MUX21X1 U711(.IN1(n366),.IN2(n365),.S(n2),.Q(n429));
  MUX21X1 U712(.IN1(n387),.IN2(n429),.S(n3),.Q(n367));
  NOR3X0 U713(.IN1(n367),.IN2(n30),.IN3(n28),.QN(N198));
  MUX21X1 U714(.IN1(n370),.IN2(n369),.S(n2),.Q(n371));
  MUX21X1 U715(.IN1(n388),.IN2(n83),.S(n3),.Q(n372));
  NOR3X0 U716(.IN1(n372),.IN2(n30),.IN3(n28),.QN(N199));
  NOR3X0 U717(.IN1(n373),.IN2(n30),.IN3(n28),.QN(N200));
  MUX21X1 U718(.IN1(n81),.IN2(n90),.S(n2),.Q(n445));
  MUX21X1 U719(.IN1(n78),.IN2(n445),.S(n3),.Q(n382));
  NOR3X0 U720(.IN1(n382),.IN2(n30),.IN3(n28),.QN(N201));
  MUX21X1 U721(.IN1(n76),.IN2(n376),.S(n3),.Q(n399));
  NOR3X0 U722(.IN1(n28),.IN2(n30),.IN3(n399),.QN(N202));
  NOR3X0 U723(.IN1(n409),.IN2(n30),.IN3(n28),.QN(N203));
  MUX21X1 U724(.IN1(n100),.IN2(n101),.S(n19),.Q(n403));
  MUX21X1 U725(.IN1(n378),.IN2(n403),.S(n17),.Q(n420));
  MUX21X1 U726(.IN1(n299),.IN2(n420),.S(n2),.Q(n444));
  MUX21X1 U727(.IN1(s_qutnt_i[8:8]),.IN2(s_qutnt_i[7:7]),.S(n19),.Q(n402));
  MUX21X1 U728(.IN1(s_qutnt_i[6:6]),.IN2(s_qutnt_i[5:5]),.S(n19),.Q(n405));
  MUX21X1 U729(.IN1(n402),.IN2(n405),.S(n17),.Q(n419));
  MUX21X1 U730(.IN1(s_qutnt_i[4:4]),.IN2(s_qutnt_i[3:3]),.S(n19),.Q(n404));
  MUX21X1 U731(.IN1(s_qutnt_i[2:2]),.IN2(s_qutnt_i[1:1]),.S(n19),.Q(n379));
  MUX21X1 U732(.IN1(n404),.IN2(n379),.S(n17),.Q(n380));
  MUX21X1 U733(.IN1(n419),.IN2(n380),.S(n2),.Q(n381));
  MUX21X1 U734(.IN1(n444),.IN2(n318),.S(n3),.Q(n383));
  MUX21X1 U735(.IN1(n383),.IN2(n382),.S(n27),.Q(n384));
  OR2X1 U736(.IN1(n385),.IN2(s_shr1[3:3]),.Q(n416));
  NOR3X0 U737(.IN1(n416),.IN2(n30),.IN3(n28),.QN(N204));
  OR2X1 U738(.IN1(n386),.IN2(s_shr1[3:3]),.Q(n423));
  NOR3X0 U739(.IN1(n423),.IN2(n30),.IN3(n28),.QN(N205));
  OR2X1 U740(.IN1(n387),.IN2(s_shr1[3:3]),.Q(n430));
  NOR3X0 U741(.IN1(n28),.IN2(n30),.IN3(n430),.QN(N206));
  OR2X1 U742(.IN1(n388),.IN2(s_shr1[3:3]),.Q(n436));
  NOR3X0 U743(.IN1(n28),.IN2(n30),.IN3(n436),.QN(N207));
  OR2X1 U744(.IN1(n389),.IN2(s_shr1[3:3]),.Q(n441));
  NOR3X0 U745(.IN1(n28),.IN2(n30),.IN3(n441),.QN(N208));
  NOR3X0 U746(.IN1(n446),.IN2(n30),.IN3(n28),.QN(N209));
  NOR3X0 U747(.IN1(n391),.IN2(n29),.IN3(n28),.QN(N210));
  MUX21X1 U748(.IN1(n393),.IN2(n324),.S(n17),.Q(n426));
  MUX21X1 U749(.IN1(n395),.IN2(n394),.S(n17),.Q(n396));
  MUX21X1 U750(.IN1(n426),.IN2(n326),.S(n2),.Q(n397));
  MUX21X1 U751(.IN1(n398),.IN2(n397),.S(n3),.Q(n400));
  MUX21X1 U752(.IN1(n400),.IN2(n399),.S(n27),.Q(n401));
  MUX21X1 U753(.IN1(n403),.IN2(n320),.S(n17),.Q(n433));
  MUX21X1 U754(.IN1(n405),.IN2(n404),.S(n17),.Q(n406));
  MUX21X1 U755(.IN1(n433),.IN2(n325),.S(n2),.Q(n407));
  MUX21X1 U756(.IN1(n408),.IN2(n407),.S(n3),.Q(n410));
  MUX21X1 U757(.IN1(n410),.IN2(n409),.S(n27),.Q(n411));
  MUX21X1 U758(.IN1(n413),.IN2(n323),.S(n2),.Q(n414));
  MUX21X1 U759(.IN1(n415),.IN2(n414),.S(n3),.Q(n417));
  MUX21X1 U760(.IN1(n417),.IN2(n416),.S(n27),.Q(n418));
  MUX21X1 U761(.IN1(n420),.IN2(n319),.S(n2),.Q(n421));
  MUX21X1 U762(.IN1(n422),.IN2(n421),.S(n3),.Q(n424));
  MUX21X1 U763(.IN1(n424),.IN2(n423),.S(n27),.Q(n425));
  MUX21X1 U764(.IN1(n427),.IN2(n426),.S(n2),.Q(n428));
  MUX21X1 U765(.IN1(n429),.IN2(n428),.S(n3),.Q(n431));
  MUX21X1 U766(.IN1(n431),.IN2(n430),.S(n27),.Q(n432));
  MUX21X1 U767(.IN1(n434),.IN2(n433),.S(n2),.Q(n435));
  MUX21X1 U768(.IN1(n83),.IN2(n435),.S(n3),.Q(n437));
  MUX21X1 U769(.IN1(n437),.IN2(n436),.S(n27),.Q(n438));
  MUX21X1 U770(.IN1(n440),.IN2(n439),.S(n3),.Q(n442));
  MUX21X1 U771(.IN1(n442),.IN2(n441),.S(n27),.Q(n443));
  MUX21X1 U772(.IN1(n445),.IN2(n444),.S(n3),.Q(n447));
  MUX21X1 U773(.IN1(n447),.IN2(n446),.S(n27),.Q(n448));
  MUX21X1 U774(.IN1(s_qutnt_i[10:10]),.IN2(s_qutnt_i[9:9]),.S(n25),.Q(N221));
  MUX21X1 U775(.IN1(s_qutnt_i[11:11]),.IN2(s_qutnt_i[10:10]),.S(n25),.Q(N222));
  MUX21X1 U776(.IN1(s_qutnt_i[12:12]),.IN2(s_qutnt_i[11:11]),.S(n25),.Q(N223));
  MUX21X1 U777(.IN1(s_qutnt_i[13:13]),.IN2(s_qutnt_i[12:12]),.S(n25),.Q(N224));
  MUX21X1 U778(.IN1(s_qutnt_i[14:14]),.IN2(s_qutnt_i[13:13]),.S(n25),.Q(N225));
  MUX21X1 U779(.IN1(s_qutnt_i[15:15]),.IN2(s_qutnt_i[14:14]),.S(n25),.Q(N226));
  MUX21X1 U780(.IN1(s_qutnt_i[16:16]),.IN2(s_qutnt_i[15:15]),.S(n25),.Q(N227));
  MUX21X1 U781(.IN1(s_qutnt_i[17:17]),.IN2(s_qutnt_i[16:16]),.S(n25),.Q(N228));
  MUX21X1 U782(.IN1(s_qutnt_i[18:18]),.IN2(s_qutnt_i[17:17]),.S(n25),.Q(N229));
  MUX21X1 U783(.IN1(s_qutnt_i[19:19]),.IN2(s_qutnt_i[18:18]),.S(n25),.Q(N230));
  MUX21X1 U784(.IN1(s_qutnt_i[1:1]),.IN2(s_qutnt_i[0:0]),.S(n25),.Q(N212));
  MUX21X1 U785(.IN1(s_qutnt_i[20:20]),.IN2(s_qutnt_i[19:19]),.S(n25),.Q(N231));
  MUX21X1 U786(.IN1(s_qutnt_i[21:21]),.IN2(s_qutnt_i[20:20]),.S(n25),.Q(N232));
  MUX21X1 U787(.IN1(s_qutnt_i[22:22]),.IN2(s_qutnt_i[21:21]),.S(n25),.Q(N233));
  MUX21X1 U788(.IN1(s_qutnt_i[23:23]),.IN2(s_qutnt_i[22:22]),.S(n25),.Q(N234));
  MUX21X1 U789(.IN1(s_qutnt_i[24:24]),.IN2(s_qutnt_i[23:23]),.S(n25),.Q(N235));
  MUX21X1 U790(.IN1(s_qutnt_i[25:25]),.IN2(s_qutnt_i[24:24]),.S(n25),.Q(N236));
  MUX21X1 U791(.IN1(s_qutnt_i[26:26]),.IN2(s_qutnt_i[25:25]),.S(n26),.Q(N237));
  MUX21X1 U792(.IN1(s_qutnt_i[2:2]),.IN2(s_qutnt_i[1:1]),.S(n26),.Q(N213));
  MUX21X1 U793(.IN1(s_qutnt_i[3:3]),.IN2(s_qutnt_i[2:2]),.S(n26),.Q(N214));
  MUX21X1 U794(.IN1(s_qutnt_i[4:4]),.IN2(s_qutnt_i[3:3]),.S(n26),.Q(N215));
  MUX21X1 U795(.IN1(s_qutnt_i[5:5]),.IN2(s_qutnt_i[4:4]),.S(n26),.Q(N216));
  MUX21X1 U796(.IN1(s_qutnt_i[6:6]),.IN2(s_qutnt_i[5:5]),.S(n26),.Q(N217));
  MUX21X1 U797(.IN1(s_qutnt_i[7:7]),.IN2(s_qutnt_i[6:6]),.S(n26),.Q(N218));
  MUX21X1 U798(.IN1(s_qutnt_i[8:8]),.IN2(s_qutnt_i[7:7]),.S(n26),.Q(N219));
  MUX21X1 U799(.IN1(s_qutnt_i[9:9]),.IN2(s_qutnt_i[8:8]),.S(n26),.Q(N220));
endmodule
module pre_norm_sqrt_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [8:0] A ;
input [8:0] B ;
output [8:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire [9:0] carry ;
// instances
  FADDX1 U2_5(.A(A[5:5]),.B(n6),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n7),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n10),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n9),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n8),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  INVX0 U1(.INP(A[6:6]),.ZN(n2));
  NAND2X0 U2(.IN1(n4),.IN2(n1),.QN(carry[8:8]));
  INVX0 U3(.INP(A[7:7]),.ZN(n4));
  AND2X1 U4(.IN1(n2),.IN2(n3),.Q(n1));
  INVX0 U5(.INP(carry[6:6]),.ZN(n3));
  XNOR2X1 U6(.IN1(carry[8:8]),.IN2(A[8:8]),.Q(DIFF[8:8]));
  INVX0 U7(.INP(B[1:1]),.ZN(n8));
  INVX0 U8(.INP(B[4:4]),.ZN(n7));
  INVX0 U9(.INP(B[3:3]),.ZN(n10));
  INVX0 U10(.INP(B[2:2]),.ZN(n9));
  INVX0 U11(.INP(B[5:5]),.ZN(n6));
  XOR2X1 U12(.IN1(n3),.IN2(A[6:6]),.Q(DIFF[6:6]));
  XOR2X1 U13(.IN1(n1),.IN2(A[7:7]),.Q(DIFF[7:7]));
  INVX0 U14(.INP(A[0:0]),.ZN(n5));
  NAND2X0 U15(.IN1(B[0:0]),.IN2(n5),.QN(carry[1:1]));
endmodule
module pre_norm_sqrt_inj (clk_i,opa_i,fracta_52_o,exp_o);
input [31:0] opa_i ;
output [51:0] fracta_52_o ;
output [7:0] exp_o ;
input clk_i ;
wire N125 ;
wire N126 ;
wire N127 ;
wire N134 ;
wire N135 ;
wire N136 ;
wire N137 ;
wire N139 ;
wire N140 ;
wire N141 ;
wire N142 ;
wire N149 ;
wire N150 ;
wire N151 ;
wire N152 ;
wire N153 ;
wire N155 ;
wire N156 ;
wire N157 ;
wire N158 ;
wire N159 ;
wire N166 ;
wire N167 ;
wire N168 ;
wire N169 ;
wire N170 ;
wire N171 ;
wire N172 ;
wire N173 ;
wire N174 ;
wire N175 ;
wire N176 ;
wire N183 ;
wire N184 ;
wire N185 ;
wire N186 ;
wire N187 ;
wire N188 ;
wire N189 ;
wire N190 ;
wire N191 ;
wire N192 ;
wire N193 ;
wire N194 ;
wire N200 ;
wire N201 ;
wire N202 ;
wire N203 ;
wire N204 ;
wire N205 ;
wire N206 ;
wire N207 ;
wire N208 ;
wire N209 ;
wire N210 ;
wire N211 ;
wire N217 ;
wire N218 ;
wire N219 ;
wire N220 ;
wire N221 ;
wire N222 ;
wire N223 ;
wire N224 ;
wire N225 ;
wire N226 ;
wire N227 ;
wire N228 ;
wire N234 ;
wire N235 ;
wire N236 ;
wire N237 ;
wire N238 ;
wire N239 ;
wire N240 ;
wire N241 ;
wire N242 ;
wire N243 ;
wire N244 ;
wire N245 ;
wire N251 ;
wire N252 ;
wire N253 ;
wire N254 ;
wire N255 ;
wire N256 ;
wire N257 ;
wire N258 ;
wire N259 ;
wire N260 ;
wire N261 ;
wire N262 ;
wire N268 ;
wire N269 ;
wire N270 ;
wire N271 ;
wire N272 ;
wire N273 ;
wire N274 ;
wire N275 ;
wire N276 ;
wire N277 ;
wire N278 ;
wire N279 ;
wire N285 ;
wire N286 ;
wire N287 ;
wire N288 ;
wire N289 ;
wire N290 ;
wire N291 ;
wire N292 ;
wire N293 ;
wire N294 ;
wire N295 ;
wire N296 ;
wire N302 ;
wire N303 ;
wire N304 ;
wire N305 ;
wire N306 ;
wire N307 ;
wire N308 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N313 ;
wire N319 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N324 ;
wire N325 ;
wire N326 ;
wire N327 ;
wire N328 ;
wire N329 ;
wire N330 ;
wire N336 ;
wire N337 ;
wire N338 ;
wire N339 ;
wire N340 ;
wire N341 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N345 ;
wire N346 ;
wire N347 ;
wire N353 ;
wire N354 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N361 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N370 ;
wire N371 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N375 ;
wire N376 ;
wire N377 ;
wire N378 ;
wire N379 ;
wire N380 ;
wire N381 ;
wire N387 ;
wire N388 ;
wire N389 ;
wire N390 ;
wire N391 ;
wire N392 ;
wire N393 ;
wire N394 ;
wire N395 ;
wire N396 ;
wire N397 ;
wire N398 ;
wire N404 ;
wire N405 ;
wire N406 ;
wire N407 ;
wire N408 ;
wire N409 ;
wire N410 ;
wire N411 ;
wire N412 ;
wire N413 ;
wire N414 ;
wire N415 ;
wire N421 ;
wire N422 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N438 ;
wire N439 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N455 ;
wire N456 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N774 ;
wire N799 ;
wire N800 ;
wire N801 ;
wire N802 ;
wire N803 ;
wire N804 ;
wire N805 ;
wire N806 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire N767 ;
wire N766 ;
wire N765 ;
wire N764 ;
wire N763 ;
wire N762 ;
wire N761 ;
wire N760 ;
wire \add_90_I24_L14036_C89/carry[5]  ;
wire \add_90_I24_L14036_C89/carry[4]  ;
wire \add_90_I24_L14036_C89/carry[3]  ;
wire \add_90_I24_L14036_C89/carry[2]  ;
wire \add_90_I23_L14036_C89/carry[5]  ;
wire \add_90_I23_L14036_C89/carry[4]  ;
wire \add_90_I23_L14036_C89/carry[3]  ;
wire \add_90_I23_L14036_C89/carry[2]  ;
wire \add_90_I22_L14036_C89/carry[5]  ;
wire \add_90_I22_L14036_C89/carry[4]  ;
wire \add_90_I22_L14036_C89/carry[3]  ;
wire \add_90_I22_L14036_C89/carry[2]  ;
wire \add_90_I21_L14036_C89/carry[5]  ;
wire \add_90_I21_L14036_C89/carry[4]  ;
wire \add_90_I21_L14036_C89/carry[3]  ;
wire \add_90_I21_L14036_C89/carry[2]  ;
wire \add_90_I20_L14036_C89/carry[5]  ;
wire \add_90_I20_L14036_C89/carry[4]  ;
wire \add_90_I20_L14036_C89/carry[3]  ;
wire \add_90_I20_L14036_C89/carry[2]  ;
wire \add_90_I19_L14036_C89/carry[5]  ;
wire \add_90_I19_L14036_C89/carry[4]  ;
wire \add_90_I19_L14036_C89/carry[3]  ;
wire \add_90_I19_L14036_C89/carry[2]  ;
wire \add_90_I18_L14036_C89/carry[5]  ;
wire \add_90_I18_L14036_C89/carry[4]  ;
wire \add_90_I18_L14036_C89/carry[3]  ;
wire \add_90_I18_L14036_C89/carry[2]  ;
wire \add_90_I17_L14036_C89/carry[5]  ;
wire \add_90_I17_L14036_C89/carry[4]  ;
wire \add_90_I17_L14036_C89/carry[3]  ;
wire \add_90_I17_L14036_C89/carry[2]  ;
wire \add_90_I16_L14036_C89/carry[5]  ;
wire \add_90_I16_L14036_C89/carry[4]  ;
wire \add_90_I16_L14036_C89/carry[3]  ;
wire \add_90_I16_L14036_C89/carry[2]  ;
wire \add_90_I15_L14036_C89/carry[5]  ;
wire \add_90_I15_L14036_C89/carry[4]  ;
wire \add_90_I15_L14036_C89/carry[3]  ;
wire \add_90_I15_L14036_C89/carry[2]  ;
wire \add_90_I14_L14036_C89/carry[5]  ;
wire \add_90_I14_L14036_C89/carry[4]  ;
wire \add_90_I14_L14036_C89/carry[3]  ;
wire \add_90_I14_L14036_C89/carry[2]  ;
wire \add_90_I13_L14036_C89/carry[5]  ;
wire \add_90_I13_L14036_C89/carry[4]  ;
wire \add_90_I13_L14036_C89/carry[3]  ;
wire \add_90_I13_L14036_C89/carry[2]  ;
wire \add_90_I12_L14036_C89/carry[5]  ;
wire \add_90_I12_L14036_C89/carry[4]  ;
wire \add_90_I12_L14036_C89/carry[3]  ;
wire \add_90_I12_L14036_C89/carry[2]  ;
wire \add_90_I11_L14036_C89/carry[5]  ;
wire \add_90_I11_L14036_C89/carry[4]  ;
wire \add_90_I11_L14036_C89/carry[3]  ;
wire \add_90_I11_L14036_C89/carry[2]  ;
wire \add_90_I10_L14036_C89/carry[5]  ;
wire \add_90_I10_L14036_C89/carry[4]  ;
wire \add_90_I10_L14036_C89/carry[3]  ;
wire \add_90_I10_L14036_C89/carry[2]  ;
wire \add_90_I9_L14036_C89/carry[5]  ;
wire \add_90_I9_L14036_C89/carry[4]  ;
wire \add_90_I9_L14036_C89/carry[3]  ;
wire \add_90_I9_L14036_C89/carry[2]  ;
wire \add_90_I8_L14036_C89/carry[5]  ;
wire \add_90_I8_L14036_C89/carry[4]  ;
wire \add_90_I8_L14036_C89/carry[3]  ;
wire \add_90_I8_L14036_C89/carry[2]  ;
wire \add_90_I7_L14036_C89/carry[4]  ;
wire \add_90_I7_L14036_C89/carry[3]  ;
wire \add_90_I7_L14036_C89/carry[2]  ;
wire \add_90_I6_L14036_C89/carry[2]  ;
wire \add_90_I6_L14036_C89/carry[3]  ;
wire \add_90_I5_L14036_C89/carry[2]  ;
wire \add_1_root_sub_0_root_sub_92/carry[2]  ;
wire \add_1_root_sub_0_root_sub_92/carry[3]  ;
wire \add_1_root_sub_0_root_sub_92/carry[4]  ;
wire \add_1_root_sub_0_root_sub_92/carry[5]  ;
wire \add_1_root_sub_0_root_sub_92/carry[6]  ;
wire \add_1_root_sub_0_root_sub_92/carry[7]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire [5:0] s_sqr_zeros_o ;
wire [8:1] s_exp_tem ;
wire [51:28] s_fracta1_52_o ;
wire SYNOPSYS_UNCONNECTED__0 ;
// instances
  DFFX1 desc1870(.D(N806),.CLK(clk_i),.Q(exp_o[7:7]));
  DFFX1 desc1871(.D(N805),.CLK(clk_i),.Q(exp_o[6:6]));
  DFFX1 desc1872(.D(N804),.CLK(clk_i),.Q(exp_o[5:5]));
  DFFX1 desc1873(.D(N803),.CLK(clk_i),.Q(exp_o[4:4]));
  DFFX1 desc1874(.D(N802),.CLK(clk_i),.Q(exp_o[3:3]));
  DFFX1 desc1875(.D(N801),.CLK(clk_i),.Q(exp_o[2:2]));
  DFFX1 desc1876(.D(N800),.CLK(clk_i),.Q(exp_o[1:1]));
  DFFX1 desc1877(.D(N799),.CLK(clk_i),.Q(exp_o[0:0]));
  NAND4X0 U112(.IN1(n84),.IN2(n85),.IN3(n86),.IN4(n87),.QN(s_sqr_zeros_o[5:5]));
  AOI222X1 U113(.IN1(N211),.IN2(n88),.IN3(n1),.IN4(n89),.IN5(N194),.IN6(n90),.QN(n87));
  AOI22X1 U114(.IN1(N228),.IN2(n91),.IN3(N245),.IN4(n92),.QN(n86));
  AO21X1 U115(.IN1(n94),.IN2(n95),.IN3(n96),.Q(n84));
  OA221X1 U116(.IN1(n43),.IN2(n97),.IN3(n44),.IN4(n98),.IN5(n99),.Q(n95));
  OA22X1 U117(.IN1(n100),.IN2(n47),.IN3(n46),.IN4(n101),.Q(n99));
  OA222X1 U118(.IN1(n45),.IN2(n102),.IN3(n42),.IN4(n103),.IN5(n104),.IN6(n105),.Q(n94));
  AO222X1 U119(.IN1(n108),.IN2(N449),.IN3(N460),.IN4(n83),.IN5(n109),.IN6(N415),.Q(n107));
  AO222X1 U120(.IN1(N381),.IN2(n110),.IN3(n111),.IN4(N432),.IN5(n112),.IN6(N398),.Q(n106));
  AO221X1 U121(.IN1(n88),.IN2(N210),.IN3(N159),.IN4(n115),.IN5(n116),.Q(n114));
  AO22X1 U122(.IN1(n90),.IN2(N193),.IN3(n89),.IN4(N176),.Q(n116));
  AO221X1 U123(.IN1(n93),.IN2(N261),.IN3(n82),.IN4(n117),.IN5(n118),.Q(n113));
  AO22X1 U124(.IN1(n92),.IN2(N244),.IN3(n91),.IN4(N227),.Q(n118));
  OA221X1 U125(.IN1(n50),.IN2(n97),.IN3(n51),.IN4(n98),.IN5(n121),.Q(n120));
  OA22X1 U126(.IN1(n100),.IN2(n54),.IN3(n53),.IN4(n101),.Q(n121));
  OA222X1 U127(.IN1(n52),.IN2(n102),.IN3(n49),.IN4(n103),.IN5(n122),.IN6(n105),.Q(n119));
  AO222X1 U128(.IN1(n108),.IN2(N448),.IN3(N459),.IN4(n83),.IN5(n109),.IN6(N414),.Q(n124));
  AO222X1 U129(.IN1(N380),.IN2(n110),.IN3(n111),.IN4(N431),.IN5(n112),.IN6(N397),.Q(n123));
  AO221X1 U130(.IN1(n88),.IN2(N209),.IN3(N158),.IN4(n115),.IN5(n127),.Q(n126));
  AO22X1 U131(.IN1(n90),.IN2(N192),.IN3(n89),.IN4(N175),.Q(n127));
  AO221X1 U132(.IN1(n93),.IN2(N260),.IN3(n82),.IN4(n128),.IN5(n129),.Q(n125));
  AO22X1 U133(.IN1(n92),.IN2(N243),.IN3(n91),.IN4(N226),.Q(n129));
  OA221X1 U134(.IN1(n198),.IN2(n97),.IN3(n199),.IN4(n98),.IN5(n132),.Q(n131));
  OA22X1 U135(.IN1(n100),.IN2(n202),.IN3(n201),.IN4(n101),.Q(n132));
  OA222X1 U136(.IN1(n200),.IN2(n102),.IN3(n197),.IN4(n103),.IN5(n133),.IN6(n105),.Q(n130));
  AO222X1 U137(.IN1(n108),.IN2(N447),.IN3(N458),.IN4(n83),.IN5(n109),.IN6(N413),.Q(n135));
  AO222X1 U138(.IN1(N379),.IN2(n110),.IN3(n111),.IN4(N430),.IN5(n112),.IN6(N396),.Q(n134));
  AO22X1 U139(.IN1(n196),.IN2(n136),.IN3(n137),.IN4(n138),.Q(s_sqr_zeros_o[2:2]));
  NAND4X0 U140(.IN1(n139),.IN2(n140),.IN3(n141),.IN4(n142),.QN(n136));
  AOI221X1 U141(.IN1(n115),.IN2(N157),.IN3(N208),.IN4(n88),.IN5(n143),.QN(n142));
  AO22X1 U142(.IN1(N174),.IN2(n89),.IN3(N191),.IN4(n90),.Q(n143));
  AOI22X1 U143(.IN1(N225),.IN2(n91),.IN3(N242),.IN4(n92),.QN(n141));
  AO21X1 U144(.IN1(n144),.IN2(n145),.IN3(n96),.Q(n139));
  OA221X1 U145(.IN1(n204),.IN2(n97),.IN3(n205),.IN4(n98),.IN5(n146),.Q(n145));
  OA22X1 U146(.IN1(n100),.IN2(n208),.IN3(n207),.IN4(n101),.Q(n146));
  OA222X1 U147(.IN1(n206),.IN2(n102),.IN3(n203),.IN4(n103),.IN5(n147),.IN6(n105),.Q(n144));
  AO222X1 U148(.IN1(n108),.IN2(N446),.IN3(N457),.IN4(n83),.IN5(n109),.IN6(N412),.Q(n149));
  AO222X1 U149(.IN1(N378),.IN2(n110),.IN3(n111),.IN4(N429),.IN5(n112),.IN6(N395),.Q(n148));
  AO22X1 U150(.IN1(n196),.IN2(n150),.IN3(n151),.IN4(N126),.Q(s_sqr_zeros_o[1:1]));
  NAND4X0 U151(.IN1(n152),.IN2(n153),.IN3(n154),.IN4(n155),.QN(n150));
  AOI221X1 U152(.IN1(n115),.IN2(N156),.IN3(N207),.IN4(n88),.IN5(n156),.QN(n155));
  AO22X1 U153(.IN1(N173),.IN2(n89),.IN3(N190),.IN4(n90),.Q(n156));
  AOI22X1 U154(.IN1(N224),.IN2(n91),.IN3(N241),.IN4(n92),.QN(n154));
  AO21X1 U155(.IN1(n157),.IN2(n158),.IN3(n96),.Q(n152));
  OA221X1 U156(.IN1(n210),.IN2(n97),.IN3(n211),.IN4(n98),.IN5(n159),.Q(n158));
  OA22X1 U157(.IN1(n100),.IN2(n214),.IN3(n213),.IN4(n101),.Q(n159));
  OA222X1 U158(.IN1(n212),.IN2(n102),.IN3(n209),.IN4(n103),.IN5(n160),.IN6(n105),.Q(n157));
  AO222X1 U159(.IN1(n108),.IN2(N445),.IN3(N456),.IN4(n83),.IN5(n109),.IN6(N411),.Q(n162));
  AO222X1 U160(.IN1(N377),.IN2(n110),.IN3(n111),.IN4(N428),.IN5(n112),.IN6(N394),.Q(n161));
  AO22X1 U161(.IN1(n163),.IN2(n78),.IN3(n196),.IN4(n164),.Q(s_sqr_zeros_o[0:0]));
  NAND4X0 U162(.IN1(n165),.IN2(n166),.IN3(n167),.IN4(n168),.QN(n164));
  AOI221X1 U163(.IN1(n115),.IN2(N155),.IN3(N206),.IN4(n88),.IN5(n169),.QN(n168));
  AO22X1 U164(.IN1(N172),.IN2(n89),.IN3(N189),.IN4(n90),.Q(n169));
  AND2X1 U165(.IN1(n170),.IN2(n171),.Q(n90));
  AOI22X1 U166(.IN1(N223),.IN2(n91),.IN3(N240),.IN4(n92),.QN(n167));
  AND2X1 U167(.IN1(n172),.IN2(n173),.Q(n91));
  AND2X1 U168(.IN1(n174),.IN2(n96),.Q(n93));
  AO21X1 U169(.IN1(n175),.IN2(n176),.IN3(n96),.Q(n165));
  OA221X1 U170(.IN1(N353),.IN2(n97),.IN3(N336),.IN4(n98),.IN5(n177),.Q(n176));
  OA22X1 U171(.IN1(n100),.IN2(N285),.IN3(N302),.IN4(n101),.Q(n177));
  OR2X1 U172(.IN1(n180),.IN2(n181),.Q(n97));
  OA222X1 U173(.IN1(N319),.IN2(n102),.IN3(N370),.IN4(n103),.IN5(n182),.IN6(n105),.Q(n175));
  AO222X1 U174(.IN1(n108),.IN2(N444),.IN3(N455),.IN4(n83),.IN5(n109),.IN6(N410),.Q(n184));
  AND2X1 U175(.IN1(n185),.IN2(n186),.Q(n109));
  AND2X1 U176(.IN1(n188),.IN2(n187),.Q(n108));
  AO222X1 U177(.IN1(N376),.IN2(n110),.IN3(n111),.IN4(N427),.IN5(n112),.IN6(N393),.Q(n183));
  OR2X1 U178(.IN1(n178),.IN2(n179),.Q(n102));
  OAI21X1 U179(.IN1(n189),.IN2(n137),.IN3(n215),.QN(n163));
  AND2X1 U180(.IN1(n39),.IN2(s_fracta1_52_o[51:51]),.Q(fracta_52_o[51:51]));
  AO22X1 U181(.IN1(n33),.IN2(s_fracta1_52_o[51:51]),.IN3(s_fracta1_52_o[50:50]),.IN4(n39),.Q(fracta_52_o[50:50]));
  AO22X1 U182(.IN1(n33),.IN2(s_fracta1_52_o[50:50]),.IN3(s_fracta1_52_o[49:49]),.IN4(n39),.Q(fracta_52_o[49:49]));
  AO22X1 U183(.IN1(s_fracta1_52_o[49:49]),.IN2(n33),.IN3(s_fracta1_52_o[48:48]),.IN4(n38),.Q(fracta_52_o[48:48]));
  AO22X1 U184(.IN1(s_fracta1_52_o[48:48]),.IN2(n34),.IN3(s_fracta1_52_o[47:47]),.IN4(n38),.Q(fracta_52_o[47:47]));
  AO22X1 U185(.IN1(s_fracta1_52_o[47:47]),.IN2(n34),.IN3(s_fracta1_52_o[46:46]),.IN4(n38),.Q(fracta_52_o[46:46]));
  AO22X1 U186(.IN1(s_fracta1_52_o[46:46]),.IN2(n34),.IN3(s_fracta1_52_o[45:45]),.IN4(n38),.Q(fracta_52_o[45:45]));
  AO22X1 U187(.IN1(s_fracta1_52_o[45:45]),.IN2(n34),.IN3(s_fracta1_52_o[44:44]),.IN4(n38),.Q(fracta_52_o[44:44]));
  AO22X1 U188(.IN1(s_fracta1_52_o[44:44]),.IN2(n34),.IN3(s_fracta1_52_o[43:43]),.IN4(n38),.Q(fracta_52_o[43:43]));
  AO22X1 U189(.IN1(s_fracta1_52_o[43:43]),.IN2(n34),.IN3(s_fracta1_52_o[42:42]),.IN4(n37),.Q(fracta_52_o[42:42]));
  AO22X1 U190(.IN1(s_fracta1_52_o[42:42]),.IN2(n34),.IN3(s_fracta1_52_o[41:41]),.IN4(n37),.Q(fracta_52_o[41:41]));
  AO22X1 U191(.IN1(s_fracta1_52_o[41:41]),.IN2(n34),.IN3(s_fracta1_52_o[40:40]),.IN4(n37),.Q(fracta_52_o[40:40]));
  AO22X1 U192(.IN1(s_fracta1_52_o[40:40]),.IN2(n34),.IN3(s_fracta1_52_o[39:39]),.IN4(n37),.Q(fracta_52_o[39:39]));
  AO22X1 U193(.IN1(s_fracta1_52_o[39:39]),.IN2(n33),.IN3(s_fracta1_52_o[38:38]),.IN4(n37),.Q(fracta_52_o[38:38]));
  AO22X1 U194(.IN1(s_fracta1_52_o[38:38]),.IN2(n33),.IN3(s_fracta1_52_o[37:37]),.IN4(n36),.Q(fracta_52_o[37:37]));
  AO22X1 U195(.IN1(s_fracta1_52_o[37:37]),.IN2(n33),.IN3(s_fracta1_52_o[36:36]),.IN4(n36),.Q(fracta_52_o[36:36]));
  AO22X1 U196(.IN1(s_fracta1_52_o[36:36]),.IN2(n33),.IN3(s_fracta1_52_o[35:35]),.IN4(n36),.Q(fracta_52_o[35:35]));
  AO22X1 U197(.IN1(s_fracta1_52_o[35:35]),.IN2(n33),.IN3(s_fracta1_52_o[34:34]),.IN4(n36),.Q(fracta_52_o[34:34]));
  AO22X1 U198(.IN1(s_fracta1_52_o[34:34]),.IN2(n33),.IN3(s_fracta1_52_o[33:33]),.IN4(n36),.Q(fracta_52_o[33:33]));
  AO22X1 U199(.IN1(s_fracta1_52_o[33:33]),.IN2(n33),.IN3(s_fracta1_52_o[32:32]),.IN4(n36),.Q(fracta_52_o[32:32]));
  AO22X1 U200(.IN1(s_fracta1_52_o[32:32]),.IN2(n33),.IN3(s_fracta1_52_o[31:31]),.IN4(n35),.Q(fracta_52_o[31:31]));
  AO22X1 U201(.IN1(s_fracta1_52_o[31:31]),.IN2(n33),.IN3(s_fracta1_52_o[30:30]),.IN4(n35),.Q(fracta_52_o[30:30]));
  AO22X1 U202(.IN1(s_fracta1_52_o[30:30]),.IN2(n33),.IN3(s_fracta1_52_o[29:29]),.IN4(n35),.Q(fracta_52_o[29:29]));
  AO22X1 U203(.IN1(s_fracta1_52_o[29:29]),.IN2(n33),.IN3(s_fracta1_52_o[28:28]),.IN4(n37),.Q(fracta_52_o[28:28]));
  AND2X1 U204(.IN1(n33),.IN2(s_fracta1_52_o[28:28]),.Q(fracta_52_o[27:27]));
  AND2X1 U205(.IN1(s_exp_tem[8:8]),.IN2(n187),.Q(N806));
  AND2X1 U206(.IN1(s_exp_tem[7:7]),.IN2(n187),.Q(N805));
  AND2X1 U207(.IN1(s_exp_tem[6:6]),.IN2(n187),.Q(N804));
  AND2X1 U208(.IN1(s_exp_tem[5:5]),.IN2(n187),.Q(N803));
  AND2X1 U209(.IN1(s_exp_tem[4:4]),.IN2(n187),.Q(N802));
  AND2X1 U210(.IN1(s_exp_tem[3:3]),.IN2(n187),.Q(N801));
  AND2X1 U211(.IN1(s_exp_tem[2:2]),.IN2(n187),.Q(N800));
  AND2X1 U212(.IN1(s_exp_tem[1:1]),.IN2(n187),.Q(N799));
  NAND3X0 U213(.IN1(n7),.IN2(n219),.IN3(n188),.QN(n187));
  OR2X1 U214(.IN1(n105),.IN2(n13),.Q(n110));
  AO22X1 U215(.IN1(N443),.IN2(n7),.IN3(n6),.IN4(N432),.Q(N449));
  AO22X1 U216(.IN1(N442),.IN2(n7),.IN3(n6),.IN4(N431),.Q(N448));
  AO22X1 U217(.IN1(N441),.IN2(n7),.IN3(n6),.IN4(N430),.Q(N447));
  AO22X1 U218(.IN1(N440),.IN2(n7),.IN3(n6),.IN4(N429),.Q(N446));
  AO22X1 U219(.IN1(N439),.IN2(n7),.IN3(n6),.IN4(N428),.Q(N445));
  AO22X1 U220(.IN1(N438),.IN2(n7),.IN3(n6),.IN4(N427),.Q(N444));
  AO22X1 U221(.IN1(N426),.IN2(n9),.IN3(n8),.IN4(N415),.Q(N432));
  AO22X1 U222(.IN1(N425),.IN2(n9),.IN3(n8),.IN4(N414),.Q(N431));
  AO22X1 U223(.IN1(N424),.IN2(n9),.IN3(n8),.IN4(N413),.Q(N430));
  AO22X1 U224(.IN1(N423),.IN2(n9),.IN3(n8),.IN4(N412),.Q(N429));
  AO22X1 U225(.IN1(N422),.IN2(n9),.IN3(n8),.IN4(N411),.Q(N428));
  AO22X1 U226(.IN1(N421),.IN2(n9),.IN3(n8),.IN4(N410),.Q(N427));
  AO22X1 U227(.IN1(N409),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N398),.Q(N415));
  AO22X1 U228(.IN1(N408),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N397),.Q(N414));
  AO22X1 U229(.IN1(N407),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N396),.Q(N413));
  AO22X1 U230(.IN1(N406),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N395),.Q(N412));
  AO22X1 U231(.IN1(N405),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N394),.Q(N411));
  AO22X1 U232(.IN1(N404),.IN2(n10),.IN3(opa_i[3:3]),.IN4(N393),.Q(N410));
  AO22X1 U233(.IN1(N392),.IN2(n12),.IN3(n11),.IN4(N381),.Q(N398));
  AO22X1 U234(.IN1(N391),.IN2(n12),.IN3(n11),.IN4(N380),.Q(N397));
  AO22X1 U235(.IN1(N390),.IN2(n12),.IN3(n11),.IN4(N379),.Q(N396));
  AO22X1 U236(.IN1(N389),.IN2(n12),.IN3(n11),.IN4(N378),.Q(N395));
  AO22X1 U237(.IN1(N388),.IN2(n12),.IN3(n11),.IN4(N377),.Q(N394));
  AO22X1 U238(.IN1(N387),.IN2(n12),.IN3(n11),.IN4(N376),.Q(N393));
  AO22X1 U239(.IN1(N375),.IN2(n14),.IN3(n13),.IN4(N364),.Q(N381));
  AO22X1 U240(.IN1(N374),.IN2(n14),.IN3(n13),.IN4(N363),.Q(N380));
  AO22X1 U241(.IN1(N373),.IN2(n14),.IN3(n13),.IN4(N362),.Q(N379));
  AO22X1 U242(.IN1(N372),.IN2(n14),.IN3(n13),.IN4(N361),.Q(N378));
  AO22X1 U243(.IN1(N371),.IN2(n14),.IN3(n13),.IN4(N360),.Q(N377));
  AO22X1 U244(.IN1(N370),.IN2(n14),.IN3(n13),.IN4(N359),.Q(N376));
  AO22X1 U245(.IN1(N358),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N347),.Q(N364));
  AO22X1 U246(.IN1(N357),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N346),.Q(N363));
  AO22X1 U247(.IN1(N356),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N345),.Q(N362));
  AO22X1 U248(.IN1(N355),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N344),.Q(N361));
  AO22X1 U249(.IN1(N354),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N343),.Q(N360));
  AO22X1 U250(.IN1(N353),.IN2(n15),.IN3(opa_i[6:6]),.IN4(N342),.Q(N359));
  AO22X1 U251(.IN1(N341),.IN2(n17),.IN3(n16),.IN4(N330),.Q(N347));
  AO22X1 U252(.IN1(N340),.IN2(n17),.IN3(n16),.IN4(N329),.Q(N346));
  AO22X1 U253(.IN1(N339),.IN2(n17),.IN3(n16),.IN4(N328),.Q(N345));
  AO22X1 U254(.IN1(N338),.IN2(n17),.IN3(n16),.IN4(N327),.Q(N344));
  AO22X1 U255(.IN1(N337),.IN2(n17),.IN3(n16),.IN4(N326),.Q(N343));
  AO22X1 U256(.IN1(N336),.IN2(n17),.IN3(n16),.IN4(N325),.Q(N342));
  AO22X1 U257(.IN1(N324),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N313),.Q(N330));
  AO22X1 U258(.IN1(N323),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N312),.Q(N329));
  AO22X1 U259(.IN1(N322),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N311),.Q(N328));
  AO22X1 U260(.IN1(N321),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N310),.Q(N327));
  AO22X1 U261(.IN1(N320),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N309),.Q(N326));
  AO22X1 U262(.IN1(N319),.IN2(n18),.IN3(opa_i[8:8]),.IN4(N308),.Q(N325));
  AO22X1 U263(.IN1(N307),.IN2(n20),.IN3(n19),.IN4(N296),.Q(N313));
  AO22X1 U264(.IN1(N306),.IN2(n20),.IN3(n19),.IN4(N295),.Q(N312));
  AO22X1 U265(.IN1(N305),.IN2(n20),.IN3(n19),.IN4(N294),.Q(N311));
  AO22X1 U266(.IN1(N304),.IN2(n20),.IN3(n19),.IN4(N293),.Q(N310));
  AO22X1 U267(.IN1(N303),.IN2(n20),.IN3(n19),.IN4(N292),.Q(N309));
  AO22X1 U268(.IN1(N302),.IN2(n20),.IN3(n19),.IN4(N291),.Q(N308));
  AO22X1 U269(.IN1(N290),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N279),.Q(N296));
  AO22X1 U270(.IN1(N289),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N278),.Q(N295));
  AO22X1 U271(.IN1(N288),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N277),.Q(N294));
  AO22X1 U272(.IN1(N287),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N276),.Q(N293));
  AO22X1 U273(.IN1(N286),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N275),.Q(N292));
  AO22X1 U274(.IN1(N285),.IN2(n21),.IN3(opa_i[10:10]),.IN4(N274),.Q(N291));
  AO22X1 U275(.IN1(N273),.IN2(n23),.IN3(n22),.IN4(N262),.Q(N279));
  AO22X1 U276(.IN1(N272),.IN2(n23),.IN3(n22),.IN4(N261),.Q(N278));
  AO22X1 U277(.IN1(N271),.IN2(n23),.IN3(n22),.IN4(N260),.Q(N277));
  AO22X1 U278(.IN1(N270),.IN2(n23),.IN3(n22),.IN4(N259),.Q(N276));
  AO22X1 U279(.IN1(N269),.IN2(n23),.IN3(n22),.IN4(N258),.Q(N275));
  AO22X1 U280(.IN1(N268),.IN2(n23),.IN3(n22),.IN4(N257),.Q(N274));
  AO22X1 U281(.IN1(N256),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N245),.Q(N262));
  AO22X1 U282(.IN1(N255),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N244),.Q(N261));
  AO22X1 U283(.IN1(N254),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N243),.Q(N260));
  AO22X1 U284(.IN1(N253),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N242),.Q(N259));
  AO22X1 U285(.IN1(N252),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N241),.Q(N258));
  AO22X1 U286(.IN1(N251),.IN2(n218),.IN3(opa_i[12:12]),.IN4(N240),.Q(N257));
  AO22X1 U287(.IN1(N239),.IN2(n25),.IN3(n24),.IN4(N228),.Q(N245));
  AO22X1 U288(.IN1(N238),.IN2(n25),.IN3(n24),.IN4(N227),.Q(N244));
  AO22X1 U289(.IN1(N237),.IN2(n25),.IN3(n24),.IN4(N226),.Q(N243));
  AO22X1 U290(.IN1(N236),.IN2(n25),.IN3(n24),.IN4(N225),.Q(N242));
  AO22X1 U291(.IN1(N235),.IN2(n25),.IN3(n24),.IN4(N224),.Q(N241));
  AO22X1 U292(.IN1(N234),.IN2(n25),.IN3(n24),.IN4(N223),.Q(N240));
  AO22X1 U293(.IN1(N222),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N211),.Q(N228));
  AO22X1 U294(.IN1(N221),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N210),.Q(N227));
  AO22X1 U295(.IN1(N220),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N209),.Q(N226));
  AO22X1 U296(.IN1(N219),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N208),.Q(N225));
  AO22X1 U297(.IN1(N218),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N207),.Q(N224));
  AO22X1 U298(.IN1(N217),.IN2(n26),.IN3(opa_i[14:14]),.IN4(N206),.Q(N223));
  AO22X1 U299(.IN1(N205),.IN2(n28),.IN3(n27),.IN4(N194),.Q(N211));
  AO22X1 U300(.IN1(N204),.IN2(n28),.IN3(n27),.IN4(N193),.Q(N210));
  AO22X1 U301(.IN1(N203),.IN2(n28),.IN3(n27),.IN4(N192),.Q(N209));
  AO22X1 U302(.IN1(N202),.IN2(n28),.IN3(n27),.IN4(N191),.Q(N208));
  AO22X1 U303(.IN1(N201),.IN2(n28),.IN3(n27),.IN4(N190),.Q(N207));
  AO22X1 U304(.IN1(N200),.IN2(n28),.IN3(n27),.IN4(N189),.Q(N206));
  AO22X1 U305(.IN1(N188),.IN2(n29),.IN3(opa_i[16:16]),.IN4(n1),.Q(N194));
  AO22X1 U306(.IN1(N187),.IN2(n29),.IN3(opa_i[16:16]),.IN4(N176),.Q(N193));
  AO22X1 U307(.IN1(N186),.IN2(n29),.IN3(opa_i[16:16]),.IN4(N175),.Q(N192));
  AO22X1 U308(.IN1(N185),.IN2(n29),.IN3(opa_i[16:16]),.IN4(N174),.Q(N191));
  AO22X1 U309(.IN1(N184),.IN2(n29),.IN3(opa_i[16:16]),.IN4(N173),.Q(N190));
  AO22X1 U310(.IN1(N183),.IN2(n29),.IN3(opa_i[16:16]),.IN4(N172),.Q(N189));
  AO22X1 U312(.IN1(N170),.IN2(n31),.IN3(n30),.IN4(N159),.Q(N176));
  AO22X1 U313(.IN1(N169),.IN2(n31),.IN3(n30),.IN4(N158),.Q(N175));
  AO22X1 U314(.IN1(N168),.IN2(n31),.IN3(n30),.IN4(N157),.Q(N174));
  AO22X1 U315(.IN1(N167),.IN2(n31),.IN3(n30),.IN4(N156),.Q(N173));
  AO22X1 U316(.IN1(N166),.IN2(n31),.IN3(n30),.IN4(N155),.Q(N172));
  AO22X1 U319(.IN1(N152),.IN2(n32),.IN3(N142),.IN4(opa_i[18:18]),.Q(N158));
  AO22X1 U320(.IN1(N151),.IN2(n32),.IN3(opa_i[18:18]),.IN4(N141),.Q(N157));
  AO22X1 U321(.IN1(N150),.IN2(n32),.IN3(opa_i[18:18]),.IN4(N140),.Q(N156));
  AO22X1 U322(.IN1(N149),.IN2(n32),.IN3(opa_i[18:18]),.IN4(N139),.Q(N155));
  AND2X1 U324(.IN1(N137),.IN2(n217),.Q(N142));
  AO22X1 U325(.IN1(N136),.IN2(n217),.IN3(opa_i[19:19]),.IN4(N127),.Q(N141));
  AO22X1 U326(.IN1(N135),.IN2(n217),.IN3(opa_i[19:19]),.IN4(N126),.Q(N140));
  AO22X1 U327(.IN1(N134),.IN2(n217),.IN3(N125),.IN4(opa_i[19:19]),.Q(N139));
  AND2X1 U329(.IN1(n191),.IN2(n192),.Q(N127));
  XOR2X1 U330(.IN1(n192),.IN2(n191),.Q(N126));
  AO21X1 U331(.IN1(n190),.IN2(n216),.IN3(n151),.Q(n192));
  XOR2X1 U332(.IN1(n193),.IN2(opa_i[20:20]),.Q(N125));
  XOR2X1 U333(.IN1(n190),.IN2(opa_i[21:21]),.Q(n193));
  XOR2X1 U334(.IN1(N774),.IN2(opa_i[22:22]),.Q(n190));
  NOR4X0 U335(.IN1(opa_i[30:30]),.IN2(opa_i[29:29]),.IN3(opa_i[28:28]),.IN4(opa_i[27:27]),.QN(n195));
  NOR4X0 U336(.IN1(opa_i[26:26]),.IN2(opa_i[25:25]),.IN3(opa_i[24:24]),.IN4(n33),.QN(n194));
  pre_norm_sqrt_DW01_sub_0_inj sub_0_root_sub_0_root_sub_92(.A({N767,N766,N765,N764,N763,N762,N761,N760,n35}),.B({1'b0,1'b0,1'b0,n3,s_sqr_zeros_o[4:0]}),.CI(1'b0),.DIFF({s_exp_tem,SYNOPSYS_UNCONNECTED__0}));
  HADDX1 desc1878(.A0(N445),.B0(N444),.C1(\add_90_I24_L14036_C89/carry[2] ),.SO(N456));
  HADDX1 desc1879(.A0(N446),.B0(\add_90_I24_L14036_C89/carry[2] ),.C1(\add_90_I24_L14036_C89/carry[3] ),.SO(N457));
  HADDX1 desc1880(.A0(N447),.B0(\add_90_I24_L14036_C89/carry[3] ),.C1(\add_90_I24_L14036_C89/carry[4] ),.SO(N458));
  HADDX1 desc1881(.A0(N448),.B0(\add_90_I24_L14036_C89/carry[4] ),.C1(\add_90_I24_L14036_C89/carry[5] ),.SO(N459));
  HADDX1 desc1882(.A0(N428),.B0(N427),.C1(\add_90_I23_L14036_C89/carry[2] ),.SO(N439));
  HADDX1 desc1883(.A0(N429),.B0(\add_90_I23_L14036_C89/carry[2] ),.C1(\add_90_I23_L14036_C89/carry[3] ),.SO(N440));
  HADDX1 desc1884(.A0(N430),.B0(\add_90_I23_L14036_C89/carry[3] ),.C1(\add_90_I23_L14036_C89/carry[4] ),.SO(N441));
  HADDX1 desc1885(.A0(N431),.B0(\add_90_I23_L14036_C89/carry[4] ),.C1(\add_90_I23_L14036_C89/carry[5] ),.SO(N442));
  HADDX1 desc1886(.A0(N411),.B0(N410),.C1(\add_90_I22_L14036_C89/carry[2] ),.SO(N422));
  HADDX1 desc1887(.A0(N412),.B0(\add_90_I22_L14036_C89/carry[2] ),.C1(\add_90_I22_L14036_C89/carry[3] ),.SO(N423));
  HADDX1 desc1888(.A0(N413),.B0(\add_90_I22_L14036_C89/carry[3] ),.C1(\add_90_I22_L14036_C89/carry[4] ),.SO(N424));
  HADDX1 desc1889(.A0(N414),.B0(\add_90_I22_L14036_C89/carry[4] ),.C1(\add_90_I22_L14036_C89/carry[5] ),.SO(N425));
  HADDX1 desc1890(.A0(N394),.B0(N393),.C1(\add_90_I21_L14036_C89/carry[2] ),.SO(N405));
  HADDX1 desc1891(.A0(N395),.B0(\add_90_I21_L14036_C89/carry[2] ),.C1(\add_90_I21_L14036_C89/carry[3] ),.SO(N406));
  HADDX1 desc1892(.A0(N396),.B0(\add_90_I21_L14036_C89/carry[3] ),.C1(\add_90_I21_L14036_C89/carry[4] ),.SO(N407));
  HADDX1 desc1893(.A0(N397),.B0(\add_90_I21_L14036_C89/carry[4] ),.C1(\add_90_I21_L14036_C89/carry[5] ),.SO(N408));
  HADDX1 desc1894(.A0(N377),.B0(N376),.C1(\add_90_I20_L14036_C89/carry[2] ),.SO(N388));
  HADDX1 desc1895(.A0(N378),.B0(\add_90_I20_L14036_C89/carry[2] ),.C1(\add_90_I20_L14036_C89/carry[3] ),.SO(N389));
  HADDX1 desc1896(.A0(N379),.B0(\add_90_I20_L14036_C89/carry[3] ),.C1(\add_90_I20_L14036_C89/carry[4] ),.SO(N390));
  HADDX1 desc1897(.A0(N380),.B0(\add_90_I20_L14036_C89/carry[4] ),.C1(\add_90_I20_L14036_C89/carry[5] ),.SO(N391));
  HADDX1 desc1898(.A0(N360),.B0(N359),.C1(\add_90_I19_L14036_C89/carry[2] ),.SO(N371));
  HADDX1 desc1899(.A0(N361),.B0(\add_90_I19_L14036_C89/carry[2] ),.C1(\add_90_I19_L14036_C89/carry[3] ),.SO(N372));
  HADDX1 desc1900(.A0(N362),.B0(\add_90_I19_L14036_C89/carry[3] ),.C1(\add_90_I19_L14036_C89/carry[4] ),.SO(N373));
  HADDX1 desc1901(.A0(N363),.B0(\add_90_I19_L14036_C89/carry[4] ),.C1(\add_90_I19_L14036_C89/carry[5] ),.SO(N374));
  HADDX1 desc1902(.A0(N343),.B0(N342),.C1(\add_90_I18_L14036_C89/carry[2] ),.SO(N354));
  HADDX1 desc1903(.A0(N344),.B0(\add_90_I18_L14036_C89/carry[2] ),.C1(\add_90_I18_L14036_C89/carry[3] ),.SO(N355));
  HADDX1 desc1904(.A0(N345),.B0(\add_90_I18_L14036_C89/carry[3] ),.C1(\add_90_I18_L14036_C89/carry[4] ),.SO(N356));
  HADDX1 desc1905(.A0(N346),.B0(\add_90_I18_L14036_C89/carry[4] ),.C1(\add_90_I18_L14036_C89/carry[5] ),.SO(N357));
  HADDX1 desc1906(.A0(N326),.B0(N325),.C1(\add_90_I17_L14036_C89/carry[2] ),.SO(N337));
  HADDX1 desc1907(.A0(N327),.B0(\add_90_I17_L14036_C89/carry[2] ),.C1(\add_90_I17_L14036_C89/carry[3] ),.SO(N338));
  HADDX1 desc1908(.A0(N328),.B0(\add_90_I17_L14036_C89/carry[3] ),.C1(\add_90_I17_L14036_C89/carry[4] ),.SO(N339));
  HADDX1 desc1909(.A0(N329),.B0(\add_90_I17_L14036_C89/carry[4] ),.C1(\add_90_I17_L14036_C89/carry[5] ),.SO(N340));
  HADDX1 desc1910(.A0(N309),.B0(N308),.C1(\add_90_I16_L14036_C89/carry[2] ),.SO(N320));
  HADDX1 desc1911(.A0(N310),.B0(\add_90_I16_L14036_C89/carry[2] ),.C1(\add_90_I16_L14036_C89/carry[3] ),.SO(N321));
  HADDX1 desc1912(.A0(N311),.B0(\add_90_I16_L14036_C89/carry[3] ),.C1(\add_90_I16_L14036_C89/carry[4] ),.SO(N322));
  HADDX1 desc1913(.A0(N312),.B0(\add_90_I16_L14036_C89/carry[4] ),.C1(\add_90_I16_L14036_C89/carry[5] ),.SO(N323));
  HADDX1 desc1914(.A0(N292),.B0(N291),.C1(\add_90_I15_L14036_C89/carry[2] ),.SO(N303));
  HADDX1 desc1915(.A0(N293),.B0(\add_90_I15_L14036_C89/carry[2] ),.C1(\add_90_I15_L14036_C89/carry[3] ),.SO(N304));
  HADDX1 desc1916(.A0(N294),.B0(\add_90_I15_L14036_C89/carry[3] ),.C1(\add_90_I15_L14036_C89/carry[4] ),.SO(N305));
  HADDX1 desc1917(.A0(N295),.B0(\add_90_I15_L14036_C89/carry[4] ),.C1(\add_90_I15_L14036_C89/carry[5] ),.SO(N306));
  HADDX1 desc1918(.A0(N275),.B0(N274),.C1(\add_90_I14_L14036_C89/carry[2] ),.SO(N286));
  HADDX1 desc1919(.A0(N276),.B0(\add_90_I14_L14036_C89/carry[2] ),.C1(\add_90_I14_L14036_C89/carry[3] ),.SO(N287));
  HADDX1 desc1920(.A0(N277),.B0(\add_90_I14_L14036_C89/carry[3] ),.C1(\add_90_I14_L14036_C89/carry[4] ),.SO(N288));
  HADDX1 desc1921(.A0(N278),.B0(\add_90_I14_L14036_C89/carry[4] ),.C1(\add_90_I14_L14036_C89/carry[5] ),.SO(N289));
  HADDX1 desc1922(.A0(N258),.B0(N257),.C1(\add_90_I13_L14036_C89/carry[2] ),.SO(N269));
  HADDX1 desc1923(.A0(N259),.B0(\add_90_I13_L14036_C89/carry[2] ),.C1(\add_90_I13_L14036_C89/carry[3] ),.SO(N270));
  HADDX1 desc1924(.A0(N260),.B0(\add_90_I13_L14036_C89/carry[3] ),.C1(\add_90_I13_L14036_C89/carry[4] ),.SO(N271));
  HADDX1 desc1925(.A0(N261),.B0(\add_90_I13_L14036_C89/carry[4] ),.C1(\add_90_I13_L14036_C89/carry[5] ),.SO(N272));
  HADDX1 desc1926(.A0(N241),.B0(N240),.C1(\add_90_I12_L14036_C89/carry[2] ),.SO(N252));
  HADDX1 desc1927(.A0(N242),.B0(\add_90_I12_L14036_C89/carry[2] ),.C1(\add_90_I12_L14036_C89/carry[3] ),.SO(N253));
  HADDX1 desc1928(.A0(N243),.B0(\add_90_I12_L14036_C89/carry[3] ),.C1(\add_90_I12_L14036_C89/carry[4] ),.SO(N254));
  HADDX1 desc1929(.A0(N244),.B0(\add_90_I12_L14036_C89/carry[4] ),.C1(\add_90_I12_L14036_C89/carry[5] ),.SO(N255));
  HADDX1 desc1930(.A0(N224),.B0(N223),.C1(\add_90_I11_L14036_C89/carry[2] ),.SO(N235));
  HADDX1 desc1931(.A0(N225),.B0(\add_90_I11_L14036_C89/carry[2] ),.C1(\add_90_I11_L14036_C89/carry[3] ),.SO(N236));
  HADDX1 desc1932(.A0(N226),.B0(\add_90_I11_L14036_C89/carry[3] ),.C1(\add_90_I11_L14036_C89/carry[4] ),.SO(N237));
  HADDX1 desc1933(.A0(N227),.B0(\add_90_I11_L14036_C89/carry[4] ),.C1(\add_90_I11_L14036_C89/carry[5] ),.SO(N238));
  HADDX1 desc1934(.A0(N207),.B0(N206),.C1(\add_90_I10_L14036_C89/carry[2] ),.SO(N218));
  HADDX1 desc1935(.A0(N208),.B0(\add_90_I10_L14036_C89/carry[2] ),.C1(\add_90_I10_L14036_C89/carry[3] ),.SO(N219));
  HADDX1 desc1936(.A0(N209),.B0(\add_90_I10_L14036_C89/carry[3] ),.C1(\add_90_I10_L14036_C89/carry[4] ),.SO(N220));
  HADDX1 desc1937(.A0(N210),.B0(\add_90_I10_L14036_C89/carry[4] ),.C1(\add_90_I10_L14036_C89/carry[5] ),.SO(N221));
  HADDX1 desc1938(.A0(N190),.B0(N189),.C1(\add_90_I9_L14036_C89/carry[2] ),.SO(N201));
  HADDX1 desc1939(.A0(N191),.B0(\add_90_I9_L14036_C89/carry[2] ),.C1(\add_90_I9_L14036_C89/carry[3] ),.SO(N202));
  HADDX1 desc1940(.A0(N192),.B0(\add_90_I9_L14036_C89/carry[3] ),.C1(\add_90_I9_L14036_C89/carry[4] ),.SO(N203));
  HADDX1 desc1941(.A0(N193),.B0(\add_90_I9_L14036_C89/carry[4] ),.C1(\add_90_I9_L14036_C89/carry[5] ),.SO(N204));
  HADDX1 desc1942(.A0(N173),.B0(N172),.C1(\add_90_I8_L14036_C89/carry[2] ),.SO(N184));
  HADDX1 desc1943(.A0(N174),.B0(\add_90_I8_L14036_C89/carry[2] ),.C1(\add_90_I8_L14036_C89/carry[3] ),.SO(N185));
  HADDX1 desc1944(.A0(N175),.B0(\add_90_I8_L14036_C89/carry[3] ),.C1(\add_90_I8_L14036_C89/carry[4] ),.SO(N186));
  HADDX1 desc1945(.A0(N176),.B0(\add_90_I8_L14036_C89/carry[4] ),.C1(\add_90_I8_L14036_C89/carry[5] ),.SO(N187));
  HADDX1 desc1946(.A0(N156),.B0(N155),.C1(\add_90_I7_L14036_C89/carry[2] ),.SO(N167));
  HADDX1 desc1947(.A0(N157),.B0(\add_90_I7_L14036_C89/carry[2] ),.C1(\add_90_I7_L14036_C89/carry[3] ),.SO(N168));
  HADDX1 desc1948(.A0(N158),.B0(\add_90_I7_L14036_C89/carry[3] ),.C1(\add_90_I7_L14036_C89/carry[4] ),.SO(N169));
  HADDX1 desc1949(.A0(N159),.B0(\add_90_I7_L14036_C89/carry[4] ),.C1(N171),.SO(N170));
  HADDX1 desc1950(.A0(N140),.B0(N139),.C1(\add_90_I6_L14036_C89/carry[2] ),.SO(N150));
  HADDX1 desc1951(.A0(N141),.B0(\add_90_I6_L14036_C89/carry[2] ),.C1(\add_90_I6_L14036_C89/carry[3] ),.SO(N151));
  HADDX1 desc1952(.A0(N142),.B0(\add_90_I6_L14036_C89/carry[3] ),.C1(N153),.SO(N152));
  HADDX1 desc1953(.A0(N126),.B0(N125),.C1(\add_90_I5_L14036_C89/carry[2] ),.SO(N135));
  HADDX1 desc1954(.A0(N127),.B0(\add_90_I5_L14036_C89/carry[2] ),.C1(N137),.SO(N136));
  NAND2X0 U3(.IN1(n181),.IN2(n15),.QN(n105));
  NAND2X0 U4(.IN1(n151),.IN2(n216),.QN(n189));
  NAND2X0 U5(.IN1(n174),.IN2(n218),.QN(n96));
  NOR2X0 U6(.IN1(s_sqr_zeros_o[5:5]),.IN2(n265),.QN(s_fracta1_52_o[45:45]));
  INVX0 U7(.INP(n306),.ZN(n66));
  INVX0 U8(.INP(s_sqr_zeros_o[5:5]),.ZN(n41));
  NOR2X0 U9(.IN1(n110),.IN2(n185),.QN(n112));
  INVX0 U10(.INP(s_sqr_zeros_o[2:2]),.ZN(n80));
  INVX0 U11(.INP(s_sqr_zeros_o[3:3]),.ZN(n81));
  INVX0 U12(.INP(s_sqr_zeros_o[4:4]),.ZN(n48));
  INVX0 U13(.INP(n323),.ZN(n62));
  NAND2X0 U14(.IN1(n323),.IN2(n81),.QN(n280));
  NAND2X0 U15(.IN1(n321),.IN2(n81),.QN(n258));
  INVX0 U16(.INP(n246),.ZN(n64));
  NOR2X0 U17(.IN1(n2),.IN2(n259),.QN(s_fracta1_52_o[44:44]));
  NOR2X0 U18(.IN1(n2),.IN2(n279),.QN(s_fracta1_52_o[47:47]));
  NOR2X0 U19(.IN1(n61),.IN2(s_sqr_zeros_o[3:3]),.QN(n319));
  NOR2X0 U20(.IN1(n3),.IN2(n272),.QN(s_fracta1_52_o[46:46]));
  NAND2X0 U21(.IN1(n119),.IN2(n120),.QN(n117));
  NAND2X0 U22(.IN1(n130),.IN2(n131),.QN(n128));
  INVX0 U23(.INP(n301),.ZN(n74));
  INVX0 U24(.INP(n292),.ZN(n72));
  INVX0 U25(.INP(n284),.ZN(n69));
  NBUFFX2 U26(.INP(n77),.Z(n4));
  NAND4X0 U27(.IN1(n84),.IN2(n85),.IN3(n86),.IN4(n87),.QN(n2));
  NBUFFX2 U28(.INP(n77),.Z(n5));
  INVX0 U29(.INP(n320),.ZN(n55));
  NOR2X0 U30(.IN1(n96),.IN2(n22),.QN(n100));
  NOR2X0 U31(.IN1(n178),.IN2(n19),.QN(n179));
  NOR2X0 U32(.IN1(n180),.IN2(n16),.QN(n181));
  NOR2X0 U33(.IN1(n110),.IN2(n11),.QN(n185));
  NOR2X0 U34(.IN1(n171),.IN2(n27),.QN(n172));
  NOR2X0 U35(.IN1(n115),.IN2(n30),.QN(n170));
  NOR2X0 U36(.IN1(n173),.IN2(n24),.QN(n174));
  NOR2X0 U37(.IN1(n186),.IN2(n8),.QN(n188));
  NOR2X0 U38(.IN1(n186),.IN2(n188),.QN(n111));
  INVX0 U39(.INP(n222),.ZN(n56));
  INVX0 U40(.INP(N343),.ZN(n210));
  INVX0 U41(.INP(N344),.ZN(n204));
  INVX0 U42(.INP(N345),.ZN(n198));
  INVX0 U43(.INP(N346),.ZN(n50));
  INVX0 U44(.INP(N347),.ZN(n43));
  NAND2X0 U45(.IN1(n179),.IN2(n180),.QN(n98));
  NAND2X0 U46(.IN1(n181),.IN2(n105),.QN(n103));
  INVX0 U47(.INP(N275),.ZN(n214));
  INVX0 U48(.INP(N276),.ZN(n208));
  INVX0 U49(.INP(N277),.ZN(n202));
  INVX0 U50(.INP(N278),.ZN(n54));
  INVX0 U51(.INP(N279),.ZN(n47));
  INVX0 U52(.INP(N309),.ZN(n212));
  INVX0 U53(.INP(N310),.ZN(n206));
  INVX0 U54(.INP(N311),.ZN(n200));
  INVX0 U55(.INP(N312),.ZN(n52));
  INVX0 U56(.INP(N313),.ZN(n45));
  NOR2X0 U57(.IN1(n173),.IN2(n174),.QN(n92));
  NAND2X0 U58(.IN1(n100),.IN2(n178),.QN(n101));
  NOR2X0 U59(.IN1(n171),.IN2(n172),.QN(n88));
  NOR2X0 U60(.IN1(n115),.IN2(n170),.QN(n89));
  INVX0 U61(.INP(n96),.ZN(n82));
  INVX0 U62(.INP(s_sqr_zeros_o[1:1]),.ZN(n79));
  OA21X1 U63(.IN1(n113),.IN2(n114),.IN3(n196),.Q(s_sqr_zeros_o[4:4]));
  NOR2X0 U64(.IN1(n3),.IN2(n296),.QN(s_fracta1_52_o[49:49]));
  INVX0 U65(.INP(n293),.ZN(n73));
  NAND2X0 U66(.IN1(n247),.IN2(n80),.QN(n273));
  NOR2X0 U67(.IN1(s_sqr_zeros_o[5:5]),.IN2(n288),.QN(s_fracta1_52_o[48:48]));
  INVX0 U68(.INP(n285),.ZN(n70));
  INVX0 U69(.INP(N291),.ZN(N302));
  INVX0 U70(.INP(N257),.ZN(N268));
  NOR2X0 U71(.IN1(n260),.IN2(s_sqr_zeros_o[2:2]),.QN(n323));
  INVX0 U72(.INP(N223),.ZN(N234));
  INVX0 U73(.INP(N155),.ZN(N166));
  INVX0 U74(.INP(N189),.ZN(N200));
  NOR2X0 U75(.IN1(n161),.IN2(n162),.QN(n160));
  NOR2X0 U76(.IN1(n148),.IN2(n149),.QN(n147));
  NOR2X0 U77(.IN1(n134),.IN2(n135),.QN(n133));
  NOR2X0 U78(.IN1(n123),.IN2(n124),.QN(n122));
  INVX0 U79(.INP(n261),.ZN(n71));
  INVX0 U80(.INP(n236),.ZN(n67));
  INVX0 U81(.INP(n254),.ZN(n68));
  OA21X1 U82(.IN1(n125),.IN2(n126),.IN3(n196),.Q(s_sqr_zeros_o[3:3]));
  INVX0 U83(.INP(n235),.ZN(n63));
  INVX0 U84(.INP(n238),.ZN(n65));
  INVX0 U85(.INP(n248),.ZN(n61));
  AND2X1 U86(.IN1(N171),.IN2(n31),.Q(n1));
  NOR2X0 U87(.IN1(n106),.IN2(n107),.QN(n104));
  INVX0 U88(.INP(n310),.ZN(n76));
  INVX0 U89(.INP(N325),.ZN(N336));
  INVX0 U90(.INP(N410),.ZN(N421));
  INVX0 U91(.INP(N376),.ZN(N387));
  INVX0 U92(.INP(N359),.ZN(N370));
  NOR2X0 U93(.IN1(n230),.IN2(s_sqr_zeros_o[2:2]),.QN(n321));
  INVX0 U94(.INP(N427),.ZN(N438));
  NOR2X0 U95(.IN1(n183),.IN2(n184),.QN(n182));
  INVX0 U96(.INP(N444),.ZN(N455));
  INVX0 U97(.INP(s_sqr_zeros_o[0:0]),.ZN(n77));
  NAND2X0 U98(.IN1(n196),.IN2(n32),.QN(n115));
  NAND2X0 U99(.IN1(n100),.IN2(n21),.QN(n178));
  NAND2X0 U100(.IN1(n172),.IN2(n26),.QN(n173));
  NAND2X0 U101(.IN1(n170),.IN2(n29),.QN(n171));
  NAND2X0 U102(.IN1(n179),.IN2(n18),.QN(n180));
  NAND2X0 U103(.IN1(n185),.IN2(n10),.QN(n186));
  INVX0 U104(.INP(n138),.ZN(n196));
  INVX0 U105(.INP(N326),.ZN(n211));
  INVX0 U106(.INP(N327),.ZN(n205));
  INVX0 U107(.INP(N328),.ZN(n199));
  INVX0 U108(.INP(N329),.ZN(n51));
  INVX0 U109(.INP(N360),.ZN(n209));
  INVX0 U110(.INP(N361),.ZN(n203));
  INVX0 U111(.INP(N362),.ZN(n197));
  INVX0 U311(.INP(N363),.ZN(n49));
  INVX0 U317(.INP(N364),.ZN(n42));
  NBUFFX2 U318(.INP(n40),.Z(n35));
  INVX0 U323(.INP(N292),.ZN(n213));
  INVX0 U328(.INP(N293),.ZN(n207));
  INVX0 U337(.INP(N294),.ZN(n201));
  INVX0 U338(.INP(N295),.ZN(n53));
  INVX0 U339(.INP(N296),.ZN(n46));
  INVX0 U340(.INP(N330),.ZN(n44));
  NAND2X0 U341(.IN1(n93),.IN2(N262),.QN(n85));
  NAND2X0 U342(.IN1(n93),.IN2(N257),.QN(n166));
  NAND2X0 U343(.IN1(n93),.IN2(N259),.QN(n140));
  NAND2X0 U344(.IN1(n93),.IN2(N258),.QN(n153));
  NBUFFX2 U345(.INP(n40),.Z(n36));
  NBUFFX2 U346(.INP(n40),.Z(n37));
  NBUFFX2 U347(.INP(n40),.Z(n38));
  NBUFFX2 U348(.INP(n40),.Z(n39));
  NAND2X0 U349(.IN1(n232),.IN2(n79),.QN(n260));
  INVX0 U350(.INP(N240),.ZN(N251));
  INVX0 U351(.INP(N274),.ZN(N285));
  INVX0 U352(.INP(N172),.ZN(N183));
  INVX0 U353(.INP(N139),.ZN(N149));
  INVX0 U354(.INP(N206),.ZN(N217));
  NOR2X0 U355(.IN1(n193),.IN2(opa_i[20:20]),.QN(n191));
  NOR2X0 U356(.IN1(n2),.IN2(n305),.QN(s_fracta1_52_o[50:50]));
  INVX0 U357(.INP(n302),.ZN(n75));
  INVX0 U358(.INP(N342),.ZN(N353));
  INVX0 U359(.INP(N308),.ZN(N319));
  INVX0 U360(.INP(N393),.ZN(N404));
  INVX0 U361(.INP(N774),.ZN(n78));
  INVX0 U362(.INP(n187),.ZN(n83));
  NOR2X0 U363(.IN1(n189),.IN2(opa_i[20:20]),.QN(n137));
  INVX0 U364(.INP(opa_i[13:13]),.ZN(n25));
  NAND2X0 U365(.IN1(n137),.IN2(n217),.QN(n138));
  INVX0 U366(.INP(n224),.ZN(n57));
  INVX0 U367(.INP(n225),.ZN(n58));
  INVX0 U368(.INP(n227),.ZN(n60));
  INVX0 U369(.INP(n226),.ZN(n59));
  INVX0 U370(.INP(opa_i[23:23]),.ZN(n40));
  INVX0 U371(.INP(opa_i[12:12]),.ZN(n218));
  INVX0 U372(.INP(opa_i[17:17]),.ZN(n31));
  INVX0 U373(.INP(opa_i[15:15]),.ZN(n28));
  INVX0 U374(.INP(opa_i[11:11]),.ZN(n23));
  INVX0 U375(.INP(opa_i[4:4]),.ZN(n12));
  INVX0 U376(.INP(opa_i[7:7]),.ZN(n17));
  INVX0 U377(.INP(opa_i[9:9]),.ZN(n20));
  INVX0 U378(.INP(n190),.ZN(n215));
  INVX0 U379(.INP(opa_i[2:2]),.ZN(n9));
  INVX0 U380(.INP(opa_i[5:5]),.ZN(n14));
  INVX0 U381(.INP(opa_i[1:1]),.ZN(n7));
  NAND2X0 U382(.IN1(n194),.IN2(n195),.QN(N774));
  NOR2X0 U383(.IN1(N774),.IN2(opa_i[22:22]),.QN(n151));
  INVX0 U384(.INP(N125),.ZN(N134));
  INVX0 U385(.INP(opa_i[0:0]),.ZN(n219));
  NAND2X0 U386(.IN1(opa_i[0:0]),.IN2(n4),.QN(n223));
  INVX0 U387(.INP(opa_i[19:19]),.ZN(n217));
  INVX0 U388(.INP(opa_i[21:21]),.ZN(n216));
  NAND4X0 U389(.IN1(n84),.IN2(n85),.IN3(n86),.IN4(n87),.QN(n3));
  INVX0 U390(.INP(n7),.ZN(n6));
  INVX0 U391(.INP(n9),.ZN(n8));
  INVX0 U392(.INP(opa_i[3:3]),.ZN(n10));
  INVX0 U393(.INP(n12),.ZN(n11));
  INVX0 U394(.INP(n14),.ZN(n13));
  INVX0 U395(.INP(opa_i[6:6]),.ZN(n15));
  INVX0 U396(.INP(n17),.ZN(n16));
  INVX0 U397(.INP(opa_i[8:8]),.ZN(n18));
  INVX0 U398(.INP(n20),.ZN(n19));
  INVX0 U399(.INP(opa_i[10:10]),.ZN(n21));
  INVX0 U400(.INP(n23),.ZN(n22));
  INVX0 U401(.INP(n25),.ZN(n24));
  INVX0 U402(.INP(opa_i[14:14]),.ZN(n26));
  INVX0 U403(.INP(n28),.ZN(n27));
  INVX0 U404(.INP(opa_i[16:16]),.ZN(n29));
  INVX0 U405(.INP(n31),.ZN(n30));
  INVX0 U406(.INP(opa_i[18:18]),.ZN(n32));
  INVX0 U407(.INP(n35),.ZN(n33));
  INVX0 U408(.INP(n35),.ZN(n34));
  AND2X1 U409(.IN1(\add_1_root_sub_0_root_sub_92/carry[7] ),.IN2(opa_i[30:30]),.Q(N767));
  XOR2X1 U410(.IN1(opa_i[30:30]),.IN2(\add_1_root_sub_0_root_sub_92/carry[7] ),.Q(N766));
  OR2X1 U411(.IN1(opa_i[29:29]),.IN2(\add_1_root_sub_0_root_sub_92/carry[6] ),.Q(\add_1_root_sub_0_root_sub_92/carry[7] ));
  XNOR2X1 U412(.IN1(\add_1_root_sub_0_root_sub_92/carry[6] ),.IN2(opa_i[29:29]),.Q(N765));
  OR2X1 U413(.IN1(opa_i[28:28]),.IN2(\add_1_root_sub_0_root_sub_92/carry[5] ),.Q(\add_1_root_sub_0_root_sub_92/carry[6] ));
  XNOR2X1 U414(.IN1(\add_1_root_sub_0_root_sub_92/carry[5] ),.IN2(opa_i[28:28]),.Q(N764));
  OR2X1 U415(.IN1(opa_i[27:27]),.IN2(\add_1_root_sub_0_root_sub_92/carry[4] ),.Q(\add_1_root_sub_0_root_sub_92/carry[5] ));
  XNOR2X1 U416(.IN1(\add_1_root_sub_0_root_sub_92/carry[4] ),.IN2(opa_i[27:27]),.Q(N763));
  OR2X1 U417(.IN1(opa_i[26:26]),.IN2(\add_1_root_sub_0_root_sub_92/carry[3] ),.Q(\add_1_root_sub_0_root_sub_92/carry[4] ));
  XNOR2X1 U418(.IN1(\add_1_root_sub_0_root_sub_92/carry[3] ),.IN2(opa_i[26:26]),.Q(N762));
  OR2X1 U419(.IN1(opa_i[25:25]),.IN2(\add_1_root_sub_0_root_sub_92/carry[2] ),.Q(\add_1_root_sub_0_root_sub_92/carry[3] ));
  XNOR2X1 U420(.IN1(\add_1_root_sub_0_root_sub_92/carry[2] ),.IN2(opa_i[25:25]),.Q(N761));
  OR2X1 U421(.IN1(opa_i[24:24]),.IN2(n33),.Q(\add_1_root_sub_0_root_sub_92/carry[2] ));
  XNOR2X1 U422(.IN1(n33),.IN2(opa_i[24:24]),.Q(N760));
  XOR2X1 U423(.IN1(\add_90_I8_L14036_C89/carry[5] ),.IN2(n1),.Q(N188));
  XOR2X1 U424(.IN1(\add_90_I9_L14036_C89/carry[5] ),.IN2(N194),.Q(N205));
  XOR2X1 U425(.IN1(\add_90_I10_L14036_C89/carry[5] ),.IN2(N211),.Q(N222));
  XOR2X1 U426(.IN1(\add_90_I11_L14036_C89/carry[5] ),.IN2(N228),.Q(N239));
  XOR2X1 U427(.IN1(\add_90_I12_L14036_C89/carry[5] ),.IN2(N245),.Q(N256));
  XOR2X1 U428(.IN1(\add_90_I13_L14036_C89/carry[5] ),.IN2(N262),.Q(N273));
  XOR2X1 U429(.IN1(\add_90_I14_L14036_C89/carry[5] ),.IN2(N279),.Q(N290));
  XOR2X1 U430(.IN1(\add_90_I15_L14036_C89/carry[5] ),.IN2(N296),.Q(N307));
  XOR2X1 U431(.IN1(\add_90_I16_L14036_C89/carry[5] ),.IN2(N313),.Q(N324));
  XOR2X1 U432(.IN1(\add_90_I17_L14036_C89/carry[5] ),.IN2(N330),.Q(N341));
  XOR2X1 U433(.IN1(\add_90_I18_L14036_C89/carry[5] ),.IN2(N347),.Q(N358));
  XOR2X1 U434(.IN1(\add_90_I19_L14036_C89/carry[5] ),.IN2(N364),.Q(N375));
  XOR2X1 U435(.IN1(\add_90_I20_L14036_C89/carry[5] ),.IN2(N381),.Q(N392));
  XOR2X1 U436(.IN1(\add_90_I21_L14036_C89/carry[5] ),.IN2(N398),.Q(N409));
  XOR2X1 U437(.IN1(\add_90_I22_L14036_C89/carry[5] ),.IN2(N415),.Q(N426));
  XOR2X1 U438(.IN1(\add_90_I23_L14036_C89/carry[5] ),.IN2(N432),.Q(N443));
  XOR2X1 U439(.IN1(\add_90_I24_L14036_C89/carry[5] ),.IN2(N449),.Q(N460));
  AND2X1 U440(.IN1(N153),.IN2(n32),.Q(N159));
  OR2X1 U443(.IN1(n223),.IN2(s_sqr_zeros_o[1:1]),.Q(n230));
  NOR3X0 U444(.IN1(n258),.IN2(n2),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[28:28]));
  MUX21X1 U445(.IN1(n6),.IN2(n8),.S(n5),.Q(n222));
  MUX21X1 U446(.IN1(n223),.IN2(n56),.S(n79),.Q(n242));
  OR2X1 U447(.IN1(n242),.IN2(s_sqr_zeros_o[2:2]),.Q(n266));
  MUX21X1 U448(.IN1(opa_i[3:3]),.IN2(n11),.S(n5),.Q(n224));
  MUX21X1 U449(.IN1(n13),.IN2(opa_i[6:6]),.S(n5),.Q(n225));
  MUX21X1 U450(.IN1(n57),.IN2(n58),.S(n79),.Q(n241));
  MUX21X1 U451(.IN1(n16),.IN2(opa_i[8:8]),.S(n5),.Q(n226));
  MUX21X1 U452(.IN1(n19),.IN2(opa_i[10:10]),.S(n5),.Q(n227));
  MUX21X1 U453(.IN1(n59),.IN2(n60),.S(n79),.Q(n244));
  MUX21X1 U454(.IN1(n241),.IN2(n244),.S(n80),.Q(n270));
  MUX21X1 U455(.IN1(n266),.IN2(n270),.S(n81),.Q(n228));
  NOR3X0 U456(.IN1(n228),.IN2(n3),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[38:38]));
  MUX21X1 U457(.IN1(opa_i[0:0]),.IN2(n6),.S(n5),.Q(n232));
  MUX21X1 U458(.IN1(n8),.IN2(opa_i[3:3]),.S(n5),.Q(n234));
  MUX21X1 U459(.IN1(n232),.IN2(n234),.S(n79),.Q(n247));
  MUX21X1 U460(.IN1(n11),.IN2(n13),.S(n5),.Q(n233));
  MUX21X1 U461(.IN1(opa_i[6:6]),.IN2(n16),.S(n5),.Q(n237));
  MUX21X1 U462(.IN1(n233),.IN2(n237),.S(n79),.Q(n246));
  MUX21X1 U463(.IN1(opa_i[8:8]),.IN2(n19),.S(n5),.Q(n236));
  MUX21X1 U464(.IN1(n21),.IN2(n23),.S(n5),.Q(n239));
  MUX21X1 U465(.IN1(n67),.IN2(n239),.S(n79),.Q(n250));
  MUX21X1 U466(.IN1(n64),.IN2(n250),.S(n80),.Q(n277));
  MUX21X1 U467(.IN1(n273),.IN2(n277),.S(n81),.Q(n229));
  NOR3X0 U468(.IN1(n229),.IN2(n2),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[39:39]));
  MUX21X1 U469(.IN1(n56),.IN2(n57),.S(n79),.Q(n253));
  MUX21X1 U470(.IN1(n230),.IN2(n253),.S(n80),.Q(n281));
  MUX21X1 U471(.IN1(n58),.IN2(n59),.S(n79),.Q(n252));
  MUX21X1 U472(.IN1(n23),.IN2(n218),.S(n5),.Q(n243));
  MUX21X1 U473(.IN1(n60),.IN2(n243),.S(n79),.Q(n255));
  MUX21X1 U474(.IN1(n252),.IN2(n255),.S(n80),.Q(n286));
  MUX21X1 U475(.IN1(n281),.IN2(n286),.S(n81),.Q(n231));
  NOR3X0 U476(.IN1(n231),.IN2(n3),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[40:40]));
  MUX21X1 U477(.IN1(n234),.IN2(n233),.S(n79),.Q(n235));
  MUX21X1 U478(.IN1(n260),.IN2(n63),.S(n80),.Q(n289));
  MUX21X1 U479(.IN1(n237),.IN2(n236),.S(n79),.Q(n238));
  MUX21X1 U480(.IN1(n218),.IN2(n25),.S(n4),.Q(n249));
  MUX21X1 U481(.IN1(n239),.IN2(n249),.S(n79),.Q(n262));
  MUX21X1 U482(.IN1(n65),.IN2(n262),.S(n80),.Q(n294));
  MUX21X1 U483(.IN1(n289),.IN2(n294),.S(n81),.Q(n240));
  NOR3X0 U484(.IN1(n240),.IN2(s_sqr_zeros_o[5:5]),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[41:41]));
  MUX21X1 U485(.IN1(n242),.IN2(n241),.S(n80),.Q(n297));
  MUX21X1 U486(.IN1(n24),.IN2(opa_i[14:14]),.S(n4),.Q(n254));
  MUX21X1 U487(.IN1(n243),.IN2(n68),.S(n79),.Q(n268));
  MUX21X1 U488(.IN1(n244),.IN2(n268),.S(n80),.Q(n303));
  MUX21X1 U489(.IN1(n297),.IN2(n303),.S(n81),.Q(n245));
  NOR3X0 U490(.IN1(s_sqr_zeros_o[4:4]),.IN2(n2),.IN3(n245),.QN(s_fracta1_52_o[42:42]));
  MUX21X1 U491(.IN1(n247),.IN2(n246),.S(n80),.Q(n248));
  MUX21X1 U492(.IN1(opa_i[14:14]),.IN2(n27),.S(n4),.Q(n261));
  MUX21X1 U493(.IN1(n249),.IN2(n71),.S(n79),.Q(n275));
  MUX21X1 U494(.IN1(n250),.IN2(n275),.S(n80),.Q(n306));
  MUX21X1 U495(.IN1(n61),.IN2(n306),.S(n81),.Q(n251));
  NOR3X0 U496(.IN1(s_sqr_zeros_o[4:4]),.IN2(n3),.IN3(n251),.QN(s_fracta1_52_o[43:43]));
  MUX21X1 U497(.IN1(n253),.IN2(n252),.S(n80),.Q(n320));
  MUX21X1 U498(.IN1(n27),.IN2(opa_i[16:16]),.S(n4),.Q(n267));
  MUX21X1 U499(.IN1(n254),.IN2(n267),.S(n79),.Q(n284));
  MUX21X1 U500(.IN1(n255),.IN2(n69),.S(n80),.Q(n256));
  MUX21X1 U501(.IN1(n320),.IN2(n256),.S(n81),.Q(n257));
  MUX21X1 U502(.IN1(n258),.IN2(n257),.S(n48),.Q(n259));
  MUX21X1 U503(.IN1(n63),.IN2(n65),.S(n80),.Q(n324));
  MUX21X1 U504(.IN1(opa_i[16:16]),.IN2(n30),.S(n4),.Q(n274));
  MUX21X1 U505(.IN1(n261),.IN2(n274),.S(n79),.Q(n292));
  MUX21X1 U506(.IN1(n262),.IN2(n72),.S(n80),.Q(n263));
  MUX21X1 U507(.IN1(n324),.IN2(n263),.S(n81),.Q(n264));
  MUX21X1 U508(.IN1(n280),.IN2(n264),.S(n48),.Q(n265));
  OR2X1 U509(.IN1(n266),.IN2(s_sqr_zeros_o[3:3]),.Q(n314));
  MUX21X1 U510(.IN1(n30),.IN2(opa_i[18:18]),.S(n4),.Q(n282));
  MUX21X1 U511(.IN1(n267),.IN2(n282),.S(n79),.Q(n301));
  MUX21X1 U512(.IN1(n268),.IN2(n74),.S(n80),.Q(n269));
  MUX21X1 U513(.IN1(n270),.IN2(n269),.S(n81),.Q(n271));
  MUX21X1 U514(.IN1(n314),.IN2(n271),.S(n48),.Q(n272));
  OR2X1 U515(.IN1(n273),.IN2(s_sqr_zeros_o[3:3]),.Q(n315));
  MUX21X1 U516(.IN1(opa_i[18:18]),.IN2(opa_i[19:19]),.S(n4),.Q(n290));
  MUX21X1 U517(.IN1(n274),.IN2(n290),.S(n79),.Q(n310));
  MUX21X1 U518(.IN1(n275),.IN2(n76),.S(n80),.Q(n276));
  MUX21X1 U519(.IN1(n277),.IN2(n276),.S(n81),.Q(n278));
  MUX21X1 U520(.IN1(n315),.IN2(n278),.S(n48),.Q(n279));
  NOR3X0 U521(.IN1(n280),.IN2(s_sqr_zeros_o[5:5]),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[29:29]));
  OR2X1 U522(.IN1(n281),.IN2(s_sqr_zeros_o[3:3]),.Q(n316));
  MUX21X1 U523(.IN1(opa_i[19:19]),.IN2(opa_i[20:20]),.S(n4),.Q(n299));
  MUX21X1 U524(.IN1(n282),.IN2(n299),.S(n79),.Q(n283));
  MUX21X1 U525(.IN1(n284),.IN2(n283),.S(n80),.Q(n285));
  MUX21X1 U526(.IN1(n286),.IN2(n70),.S(n81),.Q(n287));
  MUX21X1 U527(.IN1(n316),.IN2(n287),.S(n48),.Q(n288));
  OR2X1 U528(.IN1(n289),.IN2(s_sqr_zeros_o[3:3]),.Q(n317));
  MUX21X1 U529(.IN1(opa_i[20:20]),.IN2(opa_i[21:21]),.S(n4),.Q(n308));
  MUX21X1 U530(.IN1(n290),.IN2(n308),.S(n79),.Q(n291));
  MUX21X1 U531(.IN1(n292),.IN2(n291),.S(n80),.Q(n293));
  MUX21X1 U532(.IN1(n294),.IN2(n73),.S(n81),.Q(n295));
  MUX21X1 U533(.IN1(n317),.IN2(n295),.S(n48),.Q(n296));
  OR2X1 U534(.IN1(n297),.IN2(s_sqr_zeros_o[3:3]),.Q(n318));
  MUX21X1 U535(.IN1(opa_i[21:21]),.IN2(opa_i[22:22]),.S(n4),.Q(n298));
  MUX21X1 U536(.IN1(n299),.IN2(n298),.S(n79),.Q(n300));
  MUX21X1 U537(.IN1(n301),.IN2(n300),.S(n80),.Q(n302));
  MUX21X1 U538(.IN1(n303),.IN2(n75),.S(n81),.Q(n304));
  MUX21X1 U539(.IN1(n318),.IN2(n304),.S(n48),.Q(n305));
  MUX21X1 U540(.IN1(opa_i[22:22]),.IN2(N774),.S(n4),.Q(n307));
  MUX21X1 U541(.IN1(n308),.IN2(n307),.S(n79),.Q(n309));
  MUX21X1 U542(.IN1(n310),.IN2(n309),.S(n80),.Q(n311));
  MUX21X1 U543(.IN1(n66),.IN2(n311),.S(n81),.Q(n312));
  MUX21X1 U544(.IN1(n319),.IN2(n312),.S(n48),.Q(n313));
  AND2X1 U545(.IN1(n313),.IN2(n41),.Q(s_fracta1_52_o[51:51]));
  NOR3X0 U546(.IN1(s_sqr_zeros_o[4:4]),.IN2(n2),.IN3(n314),.QN(s_fracta1_52_o[30:30]));
  NOR3X0 U547(.IN1(s_sqr_zeros_o[4:4]),.IN2(n3),.IN3(n315),.QN(s_fracta1_52_o[31:31]));
  NOR3X0 U548(.IN1(s_sqr_zeros_o[4:4]),.IN2(s_sqr_zeros_o[5:5]),.IN3(n316),.QN(s_fracta1_52_o[32:32]));
  NOR3X0 U549(.IN1(n317),.IN2(n2),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[33:33]));
  NOR3X0 U550(.IN1(n318),.IN2(n3),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[34:34]));
  AND3X1 U551(.IN1(n319),.IN2(n41),.IN3(n48),.Q(s_fracta1_52_o[35:35]));
  MUX21X1 U552(.IN1(n321),.IN2(n55),.S(n81),.Q(n322));
  AND3X1 U553(.IN1(n48),.IN2(n41),.IN3(n322),.Q(s_fracta1_52_o[36:36]));
  MUX21X1 U554(.IN1(n62),.IN2(n324),.S(n81),.Q(n325));
  NOR3X0 U555(.IN1(n325),.IN2(s_sqr_zeros_o[5:5]),.IN3(s_sqr_zeros_o[4:4]),.QN(s_fracta1_52_o[37:37]));
assign fracta_52_o[0:0]=1'b0;
assign fracta_52_o[1:1]=1'b0;
assign fracta_52_o[2:2]=1'b0;
assign fracta_52_o[3:3]=1'b0;
assign fracta_52_o[4:4]=1'b0;
assign fracta_52_o[5:5]=1'b0;
assign fracta_52_o[6:6]=1'b0;
assign fracta_52_o[7:7]=1'b0;
assign fracta_52_o[8:8]=1'b0;
assign fracta_52_o[9:9]=1'b0;
assign fracta_52_o[10:10]=1'b0;
assign fracta_52_o[11:11]=1'b0;
assign fracta_52_o[12:12]=1'b0;
assign fracta_52_o[13:13]=1'b0;
assign fracta_52_o[14:14]=1'b0;
assign fracta_52_o[15:15]=1'b0;
assign fracta_52_o[16:16]=1'b0;
assign fracta_52_o[17:17]=1'b0;
assign fracta_52_o[18:18]=1'b0;
assign fracta_52_o[19:19]=1'b0;
assign fracta_52_o[20:20]=1'b0;
assign fracta_52_o[21:21]=1'b0;
assign fracta_52_o[22:22]=1'b0;
assign fracta_52_o[23:23]=1'b0;
assign fracta_52_o[24:24]=1'b0;
assign fracta_52_o[25:25]=1'b0;
assign fracta_52_o[26:26]=1'b0;
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_0_inj (A,B,CI,DIFF,CO);
input [25:0] A ;
input [25:0] B ;
output [25:0] DIFF ;
input CI ;
output CO ;
wire \carry[25]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
// instances
  INVX0 U1(.INP(A[0:0]),.ZN(n49));
  INVX0 U2(.INP(A[1:1]),.ZN(n35));
  INVX0 U3(.INP(A[2:2]),.ZN(n41));
  INVX0 U4(.INP(A[3:3]),.ZN(n42));
  INVX0 U5(.INP(A[4:4]),.ZN(n43));
  INVX0 U6(.INP(A[5:5]),.ZN(n44));
  INVX0 U7(.INP(A[6:6]),.ZN(n45));
  INVX0 U8(.INP(A[7:7]),.ZN(n46));
  INVX0 U9(.INP(A[8:8]),.ZN(n47));
  INVX0 U10(.INP(A[9:9]),.ZN(n48));
  INVX0 U11(.INP(A[10:10]),.ZN(n25));
  INVX0 U12(.INP(A[11:11]),.ZN(n26));
  INVX0 U13(.INP(A[12:12]),.ZN(n27));
  INVX0 U14(.INP(A[13:13]),.ZN(n28));
  INVX0 U15(.INP(A[14:14]),.ZN(n29));
  INVX0 U16(.INP(A[15:15]),.ZN(n30));
  INVX0 U17(.INP(A[16:16]),.ZN(n31));
  INVX0 U18(.INP(A[17:17]),.ZN(n32));
  INVX0 U19(.INP(A[18:18]),.ZN(n33));
  INVX0 U20(.INP(A[19:19]),.ZN(n34));
  INVX0 U21(.INP(A[20:20]),.ZN(n36));
  INVX0 U22(.INP(A[21:21]),.ZN(n37));
  INVX0 U23(.INP(A[22:22]),.ZN(n38));
  INVX0 U24(.INP(A[23:23]),.ZN(n39));
  AND2X1 U25(.IN1(n32),.IN2(n3),.Q(n1));
  AND2X1 U26(.IN1(n33),.IN2(n1),.Q(n2));
  AND2X1 U27(.IN1(n31),.IN2(n5),.Q(n3));
  AND2X1 U28(.IN1(n34),.IN2(n2),.Q(n4));
  AND2X1 U29(.IN1(n30),.IN2(n8),.Q(n5));
  AND2X1 U30(.IN1(n36),.IN2(n4),.Q(n6));
  AND2X1 U31(.IN1(n37),.IN2(n6),.Q(n7));
  AND2X1 U32(.IN1(n29),.IN2(n10),.Q(n8));
  AND2X1 U33(.IN1(n38),.IN2(n7),.Q(n9));
  AND2X1 U34(.IN1(n28),.IN2(n11),.Q(n10));
  AND2X1 U35(.IN1(n27),.IN2(n24),.Q(n11));
  AND2X1 U36(.IN1(n39),.IN2(n9),.Q(n12));
  AND2X1 U37(.IN1(n49),.IN2(B[0:0]),.Q(n13));
  AND2X1 U38(.IN1(n35),.IN2(n13),.Q(n14));
  AND2X1 U39(.IN1(n41),.IN2(n14),.Q(n15));
  AND2X1 U40(.IN1(n42),.IN2(n15),.Q(n16));
  AND2X1 U41(.IN1(n43),.IN2(n16),.Q(n17));
  AND2X1 U42(.IN1(n44),.IN2(n17),.Q(n18));
  AND2X1 U43(.IN1(n45),.IN2(n18),.Q(n19));
  AND2X1 U44(.IN1(n46),.IN2(n19),.Q(n20));
  AND2X1 U45(.IN1(n47),.IN2(n20),.Q(n21));
  AND2X1 U46(.IN1(n48),.IN2(n21),.Q(n22));
  AND2X1 U47(.IN1(n25),.IN2(n22),.Q(n23));
  AND2X1 U48(.IN1(n26),.IN2(n23),.Q(n24));
  XNOR2X1 U49(.IN1(\carry[25] ),.IN2(A[25:25]),.Q(DIFF[25:25]));
  NAND2X0 U50(.IN1(n40),.IN2(n12),.QN(\carry[25] ));
  INVX0 U51(.INP(A[24:24]),.ZN(n40));
  XOR2X1 U52(.IN1(n22),.IN2(A[10:10]),.Q(DIFF[10:10]));
  XOR2X1 U53(.IN1(n23),.IN2(A[11:11]),.Q(DIFF[11:11]));
  XOR2X1 U54(.IN1(n24),.IN2(A[12:12]),.Q(DIFF[12:12]));
  XOR2X1 U55(.IN1(n11),.IN2(A[13:13]),.Q(DIFF[13:13]));
  XOR2X1 U56(.IN1(n10),.IN2(A[14:14]),.Q(DIFF[14:14]));
  XOR2X1 U57(.IN1(n8),.IN2(A[15:15]),.Q(DIFF[15:15]));
  XOR2X1 U58(.IN1(n5),.IN2(A[16:16]),.Q(DIFF[16:16]));
  XOR2X1 U59(.IN1(n3),.IN2(A[17:17]),.Q(DIFF[17:17]));
  XOR2X1 U60(.IN1(n1),.IN2(A[18:18]),.Q(DIFF[18:18]));
  XOR2X1 U61(.IN1(n2),.IN2(A[19:19]),.Q(DIFF[19:19]));
  XOR2X1 U62(.IN1(n13),.IN2(A[1:1]),.Q(DIFF[1:1]));
  XOR2X1 U63(.IN1(n4),.IN2(A[20:20]),.Q(DIFF[20:20]));
  XOR2X1 U64(.IN1(n6),.IN2(A[21:21]),.Q(DIFF[21:21]));
  XOR2X1 U65(.IN1(n7),.IN2(A[22:22]),.Q(DIFF[22:22]));
  XOR2X1 U66(.IN1(n9),.IN2(A[23:23]),.Q(DIFF[23:23]));
  XOR2X1 U67(.IN1(n12),.IN2(A[24:24]),.Q(DIFF[24:24]));
  XOR2X1 U68(.IN1(n14),.IN2(A[2:2]),.Q(DIFF[2:2]));
  XOR2X1 U69(.IN1(n15),.IN2(A[3:3]),.Q(DIFF[3:3]));
  XOR2X1 U70(.IN1(n16),.IN2(A[4:4]),.Q(DIFF[4:4]));
  XOR2X1 U71(.IN1(n17),.IN2(A[5:5]),.Q(DIFF[5:5]));
  XOR2X1 U72(.IN1(n18),.IN2(A[6:6]),.Q(DIFF[6:6]));
  XOR2X1 U73(.IN1(n19),.IN2(A[7:7]),.Q(DIFF[7:7]));
  XOR2X1 U74(.IN1(n20),.IN2(A[8:8]),.Q(DIFF[8:8]));
  XOR2X1 U75(.IN1(n21),.IN2(A[9:9]),.Q(DIFF[9:9]));
  XOR2X1 U76(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW_cmp_0_inj (A,B,TC,GE_LT,GE_GT_EQ,GE_LT_GT_LE,EQ_NE);
input [51:0] A ;
input [51:0] B ;
input TC ;
input GE_LT ;
input GE_GT_EQ ;
output GE_LT_GT_LE ;
output EQ_NE ;
wire n2148 ;
wire n2149 ;
wire n2150 ;
wire n2151 ;
wire n2152 ;
wire n2153 ;
wire n2154 ;
wire n2155 ;
wire n2156 ;
wire n2157 ;
wire n2158 ;
wire n2159 ;
wire n2160 ;
wire n2161 ;
wire n2162 ;
wire n2163 ;
wire n2164 ;
wire n2165 ;
wire n2166 ;
wire n2167 ;
wire n2168 ;
wire n2169 ;
wire n2170 ;
wire n2171 ;
wire n2172 ;
wire n2173 ;
wire n2174 ;
wire n2175 ;
wire n2176 ;
wire n2177 ;
wire n2178 ;
wire n2179 ;
wire n2180 ;
wire n2181 ;
wire n2182 ;
wire n2183 ;
wire n2184 ;
wire n2185 ;
wire n2186 ;
wire n2187 ;
wire n2188 ;
wire n2189 ;
wire n2190 ;
wire n2191 ;
wire n2192 ;
wire n2193 ;
wire n2194 ;
wire n2195 ;
wire n2196 ;
wire n2197 ;
wire n2198 ;
wire n2199 ;
wire n2200 ;
wire n2201 ;
wire n2202 ;
wire n2203 ;
wire n2204 ;
wire n2205 ;
wire n2206 ;
wire n2207 ;
wire n2208 ;
wire n2209 ;
wire n2210 ;
wire n2211 ;
wire n2212 ;
wire n2213 ;
wire n2214 ;
wire n2215 ;
wire n2216 ;
wire n2217 ;
wire n2218 ;
wire n2219 ;
wire n2220 ;
wire n2221 ;
wire n2222 ;
wire n2223 ;
wire n2224 ;
wire n2225 ;
wire n2226 ;
wire n2227 ;
wire n2228 ;
wire n2229 ;
wire n2230 ;
wire n2231 ;
wire n2232 ;
wire n2233 ;
wire n2234 ;
wire n2235 ;
wire n2236 ;
wire n2237 ;
wire n2238 ;
wire n2239 ;
wire n2240 ;
wire n2241 ;
wire n2242 ;
wire n2243 ;
wire n2244 ;
wire n2245 ;
wire n2246 ;
wire n2247 ;
wire n2248 ;
wire n2249 ;
wire n2250 ;
wire n2251 ;
wire n2252 ;
wire n2253 ;
wire n2254 ;
wire n2255 ;
wire n2256 ;
wire n2257 ;
wire n2258 ;
wire n2259 ;
wire n2260 ;
wire n2261 ;
wire n2262 ;
wire n2263 ;
wire n2264 ;
wire n2265 ;
wire n2266 ;
wire n2267 ;
wire n2268 ;
wire n2269 ;
wire n2270 ;
wire n2271 ;
wire n2272 ;
wire n2273 ;
wire n2274 ;
wire n2275 ;
wire n2276 ;
wire n2277 ;
wire n2278 ;
wire n2279 ;
wire n2280 ;
wire n2281 ;
wire n2282 ;
wire n2283 ;
wire n2284 ;
wire n2285 ;
wire n2286 ;
wire n2287 ;
wire n2288 ;
wire n2289 ;
wire n2290 ;
wire n2291 ;
wire n2292 ;
wire n2293 ;
wire n2294 ;
wire n2295 ;
wire n2296 ;
wire n2297 ;
wire n2298 ;
wire n2299 ;
wire n2300 ;
wire n2301 ;
wire n2302 ;
wire n2303 ;
wire n2304 ;
wire n2305 ;
wire n2306 ;
wire n2307 ;
wire n2308 ;
wire n2309 ;
wire n2310 ;
wire n2311 ;
wire n2312 ;
wire n2313 ;
wire n2314 ;
wire n2315 ;
wire n2316 ;
wire n2317 ;
wire n2318 ;
wire n2319 ;
wire n2320 ;
wire n2321 ;
wire n2322 ;
wire n2323 ;
wire n2324 ;
wire n2325 ;
wire n2326 ;
wire n2327 ;
wire n2328 ;
wire n2329 ;
wire n2330 ;
wire n2331 ;
wire n2332 ;
wire n2333 ;
wire n2334 ;
wire n2335 ;
wire n2336 ;
wire n2337 ;
wire n2338 ;
wire n2339 ;
wire n2340 ;
wire n2341 ;
wire n2342 ;
wire n2343 ;
wire n2344 ;
wire n2345 ;
wire n2346 ;
wire n2347 ;
wire n2348 ;
wire n2349 ;
wire n2350 ;
wire n2351 ;
wire n2352 ;
wire n2353 ;
wire n2354 ;
wire n2355 ;
// instances
  INVX0 U1187(.INP(n2278),.ZN(n2162));
  INVX0 U1188(.INP(n2285),.ZN(n2178));
  INVX0 U1189(.INP(n2277),.ZN(n2170));
  INVX0 U1190(.INP(n2309),.ZN(n2187));
  INVX0 U1191(.INP(n2286),.ZN(n2182));
  INVX0 U1192(.INP(n2317),.ZN(n2185));
  INVX0 U1193(.INP(n2308),.ZN(n2188));
  INVX0 U1194(.INP(n2226),.ZN(n2149));
  INVX0 U1195(.INP(n2259),.ZN(n2156));
  INVX0 U1196(.INP(n2282),.ZN(n2176));
  INVX0 U1197(.INP(n2327),.ZN(n2172));
  INVX0 U1198(.INP(A[20:20]),.ZN(n2173));
  INVX0 U1199(.INP(n2264),.ZN(n2152));
  OR2X1 U1200(.IN1(n2287),.IN2(n2148),.Q(n2280));
  AND4X1 U1201(.IN1(n2182),.IN2(n2178),.IN3(n2283),.IN4(n2284),.Q(n2148));
  INVX0 U1202(.INP(A[18:18]),.ZN(n2175));
  INVX0 U1203(.INP(A[1:1]),.ZN(n2190));
  INVX0 U1204(.INP(A[14:14]),.ZN(n2180));
  INVX0 U1205(.INP(A[30:30]),.ZN(n2165));
  INVX0 U1206(.INP(A[46:46]),.ZN(n2153));
  INVX0 U1207(.INP(A[10:10]),.ZN(n2183));
  INVX0 U1208(.INP(A[26:26]),.ZN(n2168));
  INVX0 U1209(.INP(A[42:42]),.ZN(n2155));
  INVX0 U1210(.INP(n2242),.ZN(n2159));
  INVX0 U1211(.INP(A[36:36]),.ZN(n2160));
  INVX0 U1212(.INP(A[6:6]),.ZN(n2186));
  INVX0 U1213(.INP(B[12:12]),.ZN(n2199));
  INVX0 U1214(.INP(B[8:8]),.ZN(n2197));
  INVX0 U1215(.INP(B[28:28]),.ZN(n2207));
  INVX0 U1216(.INP(B[44:44]),.ZN(n2216));
  INVX0 U1217(.INP(B[24:24]),.ZN(n2205));
  INVX0 U1218(.INP(B[40:40]),.ZN(n2214));
  INVX0 U1219(.INP(B[33:33]),.ZN(n2210));
  INVX0 U1220(.INP(B[21:21]),.ZN(n2203));
  INVX0 U1221(.INP(B[5:5]),.ZN(n2195));
  INVX0 U1222(.INP(B[17:17]),.ZN(n2201));
  INVX0 U1223(.INP(B[37:37]),.ZN(n2212));
  INVX0 U1224(.INP(n2276),.ZN(n2174));
  INVX0 U1225(.INP(B[3:3]),.ZN(n2193));
  INVX0 U1226(.INP(B[7:7]),.ZN(n2196));
  INVX0 U1227(.INP(B[23:23]),.ZN(n2204));
  INVX0 U1228(.INP(B[39:39]),.ZN(n2213));
  INVX0 U1229(.INP(B[19:19]),.ZN(n2202));
  INVX0 U1230(.INP(B[35:35]),.ZN(n2211));
  INVX0 U1231(.INP(A[22:22]),.ZN(n2171));
  INVX0 U1232(.INP(B[11:11]),.ZN(n2198));
  INVX0 U1233(.INP(B[15:15]),.ZN(n2200));
  INVX0 U1234(.INP(B[27:27]),.ZN(n2206));
  INVX0 U1235(.INP(B[31:31]),.ZN(n2208));
  INVX0 U1236(.INP(B[43:43]),.ZN(n2215));
  INVX0 U1237(.INP(B[47:47]),.ZN(n2217));
  INVX0 U1238(.INP(n2340),.ZN(n2167));
  INVX0 U1239(.INP(n2342),.ZN(n2163));
  INVX0 U1240(.INP(A[38:38]),.ZN(n2158));
  INVX0 U1241(.INP(A[34:34]),.ZN(n2161));
  INVX0 U1242(.INP(A[13:13]),.ZN(n2181));
  INVX0 U1243(.INP(A[25:25]),.ZN(n2169));
  INVX0 U1244(.INP(A[41:41]),.ZN(n2157));
  INVX0 U1245(.INP(A[45:45]),.ZN(n2154));
  INVX0 U1246(.INP(B[0:0]),.ZN(n2191));
  INVX0 U1247(.INP(B[4:4]),.ZN(n2194));
  INVX0 U1248(.INP(A[9:9]),.ZN(n2184));
  INVX0 U1249(.INP(A[29:29]),.ZN(n2166));
  INVX0 U1250(.INP(n2298),.ZN(n2179));
  INVX0 U1251(.INP(n2349),.ZN(n2164));
  INVX0 U1252(.INP(A[2:2]),.ZN(n2189));
  INVX0 U1253(.INP(B[32:32]),.ZN(n2209));
  INVX0 U1254(.INP(B[50:50]),.ZN(n2218));
  INVX0 U1255(.INP(B[51:51]),.ZN(n2192));
  INVX0 U1256(.INP(A[49:49]),.ZN(n2150));
  INVX0 U1257(.INP(A[48:48]),.ZN(n2151));
  INVX0 U1258(.INP(A[16:16]),.ZN(n2177));
  AO22X1 U1259(.IN1(n2219),.IN2(n2220),.IN3(n2220),.IN4(n2221),.Q(GE_LT_GT_LE));
  NAND4X0 U1260(.IN1(n2222),.IN2(n2223),.IN3(n2224),.IN4(n2225),.QN(n2221));
  NOR3X0 U1261(.IN1(n2226),.IN2(n2227),.IN3(n2228),.QN(n2225));
  NOR2X0 U1262(.IN1(A[32:32]),.IN2(n2209),.QN(n2227));
  AOI22X1 U1263(.IN1(n2229),.IN2(n2230),.IN3(n2231),.IN4(n2149),.QN(n2220));
  NAND4X0 U1264(.IN1(n2230),.IN2(n2232),.IN3(n2233),.IN4(n2234),.QN(n2226));
  NAND2X0 U1265(.IN1(B[48:48]),.IN2(n2151),.QN(n2234));
  OA21X1 U1266(.IN1(n2222),.IN2(n2235),.IN3(n2236),.Q(n2231));
  AO221X1 U1267(.IN1(n2237),.IN2(n2238),.IN3(n2239),.IN4(n2223),.IN5(n2235),.Q(n2236));
  AND3X1 U1268(.IN1(n2159),.IN2(n2240),.IN3(n2241),.Q(n2223));
  NAND2X0 U1269(.IN1(B[36:36]),.IN2(n2160),.QN(n2240));
  OA21X1 U1270(.IN1(n2224),.IN2(n2243),.IN3(n2244),.Q(n2239));
  AO221X1 U1271(.IN1(A[33:33]),.IN2(n2210),.IN3(n2245),.IN4(A[32:32]),.IN5(n2243),.Q(n2244));
  NOR2X0 U1272(.IN1(B[32:32]),.IN2(n2228),.QN(n2245));
  NOR2X0 U1273(.IN1(n2210),.IN2(A[33:33]),.QN(n2228));
  AO22X1 U1274(.IN1(A[35:35]),.IN2(n2211),.IN3(n2246),.IN4(A[34:34]),.Q(n2243));
  NOR2X0 U1275(.IN1(B[34:34]),.IN2(n2247),.QN(n2246));
  AOI21X1 U1276(.IN1(B[34:34]),.IN2(n2161),.IN3(n2247),.QN(n2224));
  NOR2X0 U1277(.IN1(n2211),.IN2(A[35:35]),.QN(n2247));
  OR2X1 U1278(.IN1(n2248),.IN2(n2241),.Q(n2238));
  AOI21X1 U1279(.IN1(B[38:38]),.IN2(n2158),.IN3(n2249),.QN(n2241));
  AO221X1 U1280(.IN1(A[37:37]),.IN2(n2212),.IN3(n2250),.IN4(A[36:36]),.IN5(n2248),.Q(n2237));
  AO22X1 U1281(.IN1(A[39:39]),.IN2(n2213),.IN3(n2251),.IN4(A[38:38]),.Q(n2248));
  NOR2X0 U1282(.IN1(B[38:38]),.IN2(n2249),.QN(n2251));
  NOR2X0 U1283(.IN1(n2213),.IN2(A[39:39]),.QN(n2249));
  NOR2X0 U1284(.IN1(B[36:36]),.IN2(n2242),.QN(n2250));
  NOR2X0 U1285(.IN1(n2212),.IN2(A[37:37]),.QN(n2242));
  NAND2X0 U1286(.IN1(n2252),.IN2(n2253),.QN(n2235));
  AO221X1 U1287(.IN1(n2254),.IN2(n2255),.IN3(n2256),.IN4(n2254),.IN5(n2257),.Q(n2253));
  OA21X1 U1288(.IN1(B[41:41]),.IN2(n2157),.IN3(n2258),.Q(n2256));
  NAND3X0 U1289(.IN1(n2259),.IN2(n2214),.IN3(A[40:40]),.QN(n2258));
  AOI22X1 U1290(.IN1(A[43:43]),.IN2(n2215),.IN3(n2260),.IN4(A[42:42]),.QN(n2254));
  NOR2X0 U1291(.IN1(B[42:42]),.IN2(n2261),.QN(n2260));
  AO22X1 U1292(.IN1(n2262),.IN2(n2263),.IN3(n2263),.IN4(n2264),.Q(n2252));
  AOI22X1 U1293(.IN1(A[47:47]),.IN2(n2217),.IN3(n2265),.IN4(A[46:46]),.QN(n2263));
  NOR2X0 U1294(.IN1(B[46:46]),.IN2(n2266),.QN(n2265));
  OA21X1 U1295(.IN1(B[45:45]),.IN2(n2154),.IN3(n2267),.Q(n2262));
  NAND3X0 U1296(.IN1(n2268),.IN2(n2216),.IN3(A[44:44]),.QN(n2267));
  NOR4X0 U1297(.IN1(n2255),.IN2(n2257),.IN3(n2156),.IN4(n2269),.QN(n2222));
  NOR2X0 U1298(.IN1(n2214),.IN2(A[40:40]),.QN(n2269));
  NAND2X0 U1299(.IN1(B[41:41]),.IN2(n2157),.QN(n2259));
  NAND3X0 U1300(.IN1(n2268),.IN2(n2270),.IN3(n2152),.QN(n2257));
  AO21X1 U1301(.IN1(B[46:46]),.IN2(n2153),.IN3(n2266),.Q(n2264));
  NOR2X0 U1302(.IN1(n2217),.IN2(A[47:47]),.QN(n2266));
  OR2X1 U1303(.IN1(n2216),.IN2(A[44:44]),.Q(n2270));
  NAND2X0 U1304(.IN1(B[45:45]),.IN2(n2154),.QN(n2268));
  AO21X1 U1305(.IN1(B[42:42]),.IN2(n2155),.IN3(n2261),.Q(n2255));
  NOR2X0 U1306(.IN1(n2215),.IN2(A[43:43]),.QN(n2261));
  OR2X1 U1307(.IN1(n2192),.IN2(A[51:51]),.Q(n2230));
  AO221X1 U1308(.IN1(A[50:50]),.IN2(n2218),.IN3(A[51:51]),.IN4(n2192),.IN5(n2271),.Q(n2229));
  AND3X1 U1309(.IN1(n2272),.IN2(n2233),.IN3(n2232),.Q(n2271));
  OR2X1 U1310(.IN1(n2218),.IN2(A[50:50]),.Q(n2232));
  NAND2X0 U1311(.IN1(B[49:49]),.IN2(n2150),.QN(n2233));
  OAI22X1 U1312(.IN1(B[48:48]),.IN2(n2151),.IN3(B[49:49]),.IN4(n2150),.QN(n2272));
  NOR2X0 U1313(.IN1(n2273),.IN2(n2274),.QN(n2219));
  NOR4X0 U1314(.IN1(n2275),.IN2(n2276),.IN3(n2277),.IN4(n2278),.QN(n2274));
  NAND4X0 U1315(.IN1(n2279),.IN2(n2280),.IN3(n2176),.IN4(n2281),.QN(n2275));
  NAND2X0 U1316(.IN1(B[16:16]),.IN2(n2177),.QN(n2281));
  OR2X1 U1317(.IN1(n2197),.IN2(A[8:8]),.Q(n2284));
  AO221X1 U1318(.IN1(n2288),.IN2(n2289),.IN3(n2290),.IN4(n2291),.IN5(n2287),.Q(n2279));
  NAND2X0 U1319(.IN1(n2292),.IN2(n2293),.QN(n2287));
  AO221X1 U1320(.IN1(n2294),.IN2(n2286),.IN3(n2295),.IN4(n2294),.IN5(n2285),.Q(n2293));
  NAND3X0 U1321(.IN1(n2296),.IN2(n2297),.IN3(n2179),.QN(n2285));
  OR2X1 U1322(.IN1(n2199),.IN2(A[12:12]),.Q(n2297));
  OA21X1 U1323(.IN1(B[9:9]),.IN2(n2184),.IN3(n2299),.Q(n2295));
  NAND3X0 U1324(.IN1(n2283),.IN2(n2197),.IN3(A[8:8]),.QN(n2299));
  NAND2X0 U1325(.IN1(B[9:9]),.IN2(n2184),.QN(n2283));
  AO21X1 U1326(.IN1(B[10:10]),.IN2(n2183),.IN3(n2300),.Q(n2286));
  AOI22X1 U1327(.IN1(A[11:11]),.IN2(n2198),.IN3(n2301),.IN4(A[10:10]),.QN(n2294));
  NOR2X0 U1328(.IN1(B[10:10]),.IN2(n2300),.QN(n2301));
  NOR2X0 U1329(.IN1(n2198),.IN2(A[11:11]),.QN(n2300));
  AO22X1 U1330(.IN1(n2302),.IN2(n2303),.IN3(n2303),.IN4(n2298),.Q(n2292));
  AO21X1 U1331(.IN1(B[14:14]),.IN2(n2180),.IN3(n2304),.Q(n2298));
  AOI22X1 U1332(.IN1(A[15:15]),.IN2(n2200),.IN3(n2305),.IN4(A[14:14]),.QN(n2303));
  NOR2X0 U1333(.IN1(B[14:14]),.IN2(n2304),.QN(n2305));
  NOR2X0 U1334(.IN1(n2200),.IN2(A[15:15]),.QN(n2304));
  OA21X1 U1335(.IN1(B[13:13]),.IN2(n2181),.IN3(n2306),.Q(n2302));
  NAND3X0 U1336(.IN1(n2296),.IN2(n2199),.IN3(A[12:12]),.QN(n2306));
  NAND2X0 U1337(.IN1(B[13:13]),.IN2(n2181),.QN(n2296));
  OA221X1 U1338(.IN1(n2307),.IN2(n2308),.IN3(A[4:4]),.IN4(n2194),.IN5(n2187),.Q(n2291));
  AOI21X1 U1339(.IN1(n2189),.IN2(B[2:2]),.IN3(n2310),.QN(n2307));
  NOR2X0 U1340(.IN1(n2311),.IN2(n2312),.QN(n2290));
  OA221X1 U1341(.IN1(n2313),.IN2(n2314),.IN3(B[1:1]),.IN4(n2190),.IN5(n2188),.Q(n2311));
  AO22X1 U1342(.IN1(A[3:3]),.IN2(n2193),.IN3(n2315),.IN4(A[2:2]),.Q(n2308));
  NOR2X0 U1343(.IN1(B[2:2]),.IN2(n2310),.QN(n2315));
  NOR2X0 U1344(.IN1(n2193),.IN2(A[3:3]),.QN(n2310));
  NOR2X0 U1345(.IN1(A[0:0]),.IN2(n2191),.QN(n2314));
  AND2X1 U1346(.IN1(n2190),.IN2(B[1:1]),.Q(n2313));
  NAND2X0 U1347(.IN1(n2185),.IN2(n2312),.QN(n2289));
  AO21X1 U1348(.IN1(B[6:6]),.IN2(n2186),.IN3(n2316),.Q(n2312));
  AO221X1 U1349(.IN1(A[5:5]),.IN2(n2195),.IN3(n2318),.IN4(A[4:4]),.IN5(n2317),.Q(n2288));
  AO22X1 U1350(.IN1(A[7:7]),.IN2(n2196),.IN3(n2319),.IN4(A[6:6]),.Q(n2317));
  NOR2X0 U1351(.IN1(B[6:6]),.IN2(n2316),.QN(n2319));
  NOR2X0 U1352(.IN1(n2196),.IN2(A[7:7]),.QN(n2316));
  NOR2X0 U1353(.IN1(B[4:4]),.IN2(n2309),.QN(n2318));
  NOR2X0 U1354(.IN1(n2195),.IN2(A[5:5]),.QN(n2309));
  OA21X1 U1355(.IN1(n2162),.IN2(n2320),.IN3(n2321),.Q(n2273));
  AO221X1 U1356(.IN1(n2322),.IN2(n2323),.IN3(n2324),.IN4(n2170),.IN5(n2320),.Q(n2321));
  NAND3X0 U1357(.IN1(n2172),.IN2(n2325),.IN3(n2326),.QN(n2277));
  NAND2X0 U1358(.IN1(B[20:20]),.IN2(n2173),.QN(n2325));
  OA21X1 U1359(.IN1(n2174),.IN2(n2328),.IN3(n2329),.Q(n2324));
  AO221X1 U1360(.IN1(A[17:17]),.IN2(n2201),.IN3(n2330),.IN4(A[16:16]),.IN5(n2328),.Q(n2329));
  NOR2X0 U1361(.IN1(B[16:16]),.IN2(n2282),.QN(n2330));
  NOR2X0 U1362(.IN1(n2201),.IN2(A[17:17]),.QN(n2282));
  AO22X1 U1363(.IN1(A[19:19]),.IN2(n2202),.IN3(n2331),.IN4(A[18:18]),.Q(n2328));
  NOR2X0 U1364(.IN1(B[18:18]),.IN2(n2332),.QN(n2331));
  AO21X1 U1365(.IN1(B[18:18]),.IN2(n2175),.IN3(n2332),.Q(n2276));
  NOR2X0 U1366(.IN1(n2202),.IN2(A[19:19]),.QN(n2332));
  OR2X1 U1367(.IN1(n2333),.IN2(n2326),.Q(n2323));
  AOI21X1 U1368(.IN1(B[22:22]),.IN2(n2171),.IN3(n2334),.QN(n2326));
  AO221X1 U1369(.IN1(A[21:21]),.IN2(n2203),.IN3(n2335),.IN4(A[20:20]),.IN5(n2333),.Q(n2322));
  AO22X1 U1370(.IN1(A[23:23]),.IN2(n2204),.IN3(n2336),.IN4(A[22:22]),.Q(n2333));
  NOR2X0 U1371(.IN1(B[22:22]),.IN2(n2334),.QN(n2336));
  NOR2X0 U1372(.IN1(n2204),.IN2(A[23:23]),.QN(n2334));
  NOR2X0 U1373(.IN1(B[20:20]),.IN2(n2327),.QN(n2335));
  NOR2X0 U1374(.IN1(n2203),.IN2(A[21:21]),.QN(n2327));
  NAND2X0 U1375(.IN1(n2337),.IN2(n2338),.QN(n2320));
  AO221X1 U1376(.IN1(n2339),.IN2(n2340),.IN3(n2341),.IN4(n2339),.IN5(n2342),.Q(n2338));
  OA21X1 U1377(.IN1(B[25:25]),.IN2(n2169),.IN3(n2343),.Q(n2341));
  NAND3X0 U1378(.IN1(n2344),.IN2(n2205),.IN3(A[24:24]),.QN(n2343));
  AOI22X1 U1379(.IN1(A[27:27]),.IN2(n2206),.IN3(n2345),.IN4(A[26:26]),.QN(n2339));
  NOR2X0 U1380(.IN1(B[26:26]),.IN2(n2346),.QN(n2345));
  AO22X1 U1381(.IN1(n2347),.IN2(n2348),.IN3(n2348),.IN4(n2349),.Q(n2337));
  AOI22X1 U1382(.IN1(A[31:31]),.IN2(n2208),.IN3(n2350),.IN4(A[30:30]),.QN(n2348));
  NOR2X0 U1383(.IN1(B[30:30]),.IN2(n2351),.QN(n2350));
  OA21X1 U1384(.IN1(B[29:29]),.IN2(n2166),.IN3(n2352),.Q(n2347));
  NAND3X0 U1385(.IN1(n2353),.IN2(n2207),.IN3(A[28:28]),.QN(n2352));
  NAND4X0 U1386(.IN1(n2167),.IN2(n2163),.IN3(n2344),.IN4(n2354),.QN(n2278));
  OR2X1 U1387(.IN1(n2205),.IN2(A[24:24]),.Q(n2354));
  NAND2X0 U1388(.IN1(B[25:25]),.IN2(n2169),.QN(n2344));
  NAND3X0 U1389(.IN1(n2353),.IN2(n2355),.IN3(n2164),.QN(n2342));
  AO21X1 U1390(.IN1(B[30:30]),.IN2(n2165),.IN3(n2351),.Q(n2349));
  NOR2X0 U1391(.IN1(n2208),.IN2(A[31:31]),.QN(n2351));
  OR2X1 U1392(.IN1(n2207),.IN2(A[28:28]),.Q(n2355));
  NAND2X0 U1393(.IN1(B[29:29]),.IN2(n2166),.QN(n2353));
  AO21X1 U1394(.IN1(B[26:26]),.IN2(n2168),.IN3(n2346),.Q(n2340));
  NOR2X0 U1395(.IN1(n2206),.IN2(A[27:27]),.QN(n2346));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_0_inj (A,B,CI,SUM,CO);
input [51:0] A ;
input [51:0] B ;
output [51:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire [51:1] carry ;
// instances
  FADDX1 U1_50(.A(A[50:50]),.B(B[50:50]),.CI(carry[50:50]),.CO(carry[51:51]),.S(SUM[50:50]));
  FADDX1 U1_49(.A(A[49:49]),.B(B[49:49]),.CI(carry[49:49]),.CO(carry[50:50]),.S(SUM[49:49]));
  FADDX1 U1_48(.A(A[48:48]),.B(B[48:48]),.CI(carry[48:48]),.CO(carry[49:49]),.S(SUM[48:48]));
  FADDX1 U1_47(.A(A[47:47]),.B(B[47:47]),.CI(carry[47:47]),.CO(carry[48:48]),.S(SUM[47:47]));
  FADDX1 U1_46(.A(A[46:46]),.B(B[46:46]),.CI(carry[46:46]),.CO(carry[47:47]),.S(SUM[46:46]));
  FADDX1 U1_45(.A(A[45:45]),.B(B[45:45]),.CI(carry[45:45]),.CO(carry[46:46]),.S(SUM[45:45]));
  FADDX1 U1_44(.A(A[44:44]),.B(B[44:44]),.CI(carry[44:44]),.CO(carry[45:45]),.S(SUM[44:44]));
  FADDX1 U1_43(.A(A[43:43]),.B(B[43:43]),.CI(carry[43:43]),.CO(carry[44:44]),.S(SUM[43:43]));
  FADDX1 U1_42(.A(A[42:42]),.B(B[42:42]),.CI(carry[42:42]),.CO(carry[43:43]),.S(SUM[42:42]));
  FADDX1 U1_41(.A(A[41:41]),.B(B[41:41]),.CI(carry[41:41]),.CO(carry[42:42]),.S(SUM[41:41]));
  FADDX1 U1_40(.A(A[40:40]),.B(B[40:40]),.CI(carry[40:40]),.CO(carry[41:41]),.S(SUM[40:40]));
  FADDX1 U1_39(.A(A[39:39]),.B(B[39:39]),.CI(carry[39:39]),.CO(carry[40:40]),.S(SUM[39:39]));
  FADDX1 U1_38(.A(A[38:38]),.B(B[38:38]),.CI(carry[38:38]),.CO(carry[39:39]),.S(SUM[38:38]));
  FADDX1 U1_37(.A(A[37:37]),.B(B[37:37]),.CI(carry[37:37]),.CO(carry[38:38]),.S(SUM[37:37]));
  FADDX1 U1_36(.A(A[36:36]),.B(B[36:36]),.CI(carry[36:36]),.CO(carry[37:37]),.S(SUM[36:36]));
  FADDX1 U1_35(.A(A[35:35]),.B(B[35:35]),.CI(carry[35:35]),.CO(carry[36:36]),.S(SUM[35:35]));
  FADDX1 U1_34(.A(A[34:34]),.B(B[34:34]),.CI(carry[34:34]),.CO(carry[35:35]),.S(SUM[34:34]));
  FADDX1 U1_33(.A(A[33:33]),.B(B[33:33]),.CI(carry[33:33]),.CO(carry[34:34]),.S(SUM[33:33]));
  FADDX1 U1_32(.A(A[32:32]),.B(B[32:32]),.CI(carry[32:32]),.CO(carry[33:33]),.S(SUM[32:32]));
  FADDX1 U1_31(.A(A[31:31]),.B(B[31:31]),.CI(carry[31:31]),.CO(carry[32:32]),.S(SUM[31:31]));
  FADDX1 U1_30(.A(A[30:30]),.B(B[30:30]),.CI(carry[30:30]),.CO(carry[31:31]),.S(SUM[30:30]));
  FADDX1 U1_29(.A(A[29:29]),.B(B[29:29]),.CI(carry[29:29]),.CO(carry[30:30]),.S(SUM[29:29]));
  FADDX1 U1_28(.A(A[28:28]),.B(B[28:28]),.CI(carry[28:28]),.CO(carry[29:29]),.S(SUM[28:28]));
  FADDX1 U1_27(.A(A[27:27]),.B(B[27:27]),.CI(carry[27:27]),.CO(carry[28:28]),.S(SUM[27:27]));
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(carry[26:26]),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_25(.A(A[25:25]),.B(B[25:25]),.CI(carry[25:25]),.CO(carry[26:26]),.S(SUM[25:25]));
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(carry[24:24]),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(carry[13:13]),.CO(carry[14:14]),.S(SUM[13:13]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(carry[12:12]),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_11(.A(A[11:11]),.B(B[11:11]),.CI(carry[11:11]),.CO(carry[12:12]),.S(SUM[11:11]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(carry[10:10]),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_9(.A(A[9:9]),.B(B[9:9]),.CI(carry[9:9]),.CO(carry[10:10]),.S(SUM[9:9]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(carry[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  XOR3X1 U1_51(.IN1(A[51:51]),.IN2(B[51:51]),.IN3(carry[51:51]),.Q(SUM[51:51]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  XOR2X1 U2(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_1_inj (A,B,CI,DIFF,CO);
input [51:0] A ;
input [51:0] B ;
output [51:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire [52:0] carry ;
// instances
  FADDX1 U2_50(.A(A[50:50]),.B(n51),.CI(carry[50:50]),.CO(carry[51:51]),.S(DIFF[50:50]));
  FADDX1 U2_49(.A(A[49:49]),.B(n50),.CI(carry[49:49]),.CO(carry[50:50]),.S(DIFF[49:49]));
  FADDX1 U2_48(.A(A[48:48]),.B(n49),.CI(carry[48:48]),.CO(carry[49:49]),.S(DIFF[48:48]));
  FADDX1 U2_47(.A(A[47:47]),.B(n48),.CI(carry[47:47]),.CO(carry[48:48]),.S(DIFF[47:47]));
  FADDX1 U2_46(.A(A[46:46]),.B(n47),.CI(carry[46:46]),.CO(carry[47:47]),.S(DIFF[46:46]));
  FADDX1 U2_45(.A(A[45:45]),.B(n46),.CI(carry[45:45]),.CO(carry[46:46]),.S(DIFF[45:45]));
  FADDX1 U2_44(.A(A[44:44]),.B(n45),.CI(carry[44:44]),.CO(carry[45:45]),.S(DIFF[44:44]));
  FADDX1 U2_43(.A(A[43:43]),.B(n44),.CI(carry[43:43]),.CO(carry[44:44]),.S(DIFF[43:43]));
  FADDX1 U2_42(.A(A[42:42]),.B(n43),.CI(carry[42:42]),.CO(carry[43:43]),.S(DIFF[42:42]));
  FADDX1 U2_41(.A(A[41:41]),.B(n42),.CI(carry[41:41]),.CO(carry[42:42]),.S(DIFF[41:41]));
  FADDX1 U2_40(.A(A[40:40]),.B(n21),.CI(carry[40:40]),.CO(carry[41:41]),.S(DIFF[40:40]));
  FADDX1 U2_39(.A(A[39:39]),.B(n41),.CI(carry[39:39]),.CO(carry[40:40]),.S(DIFF[39:39]));
  FADDX1 U2_38(.A(A[38:38]),.B(n20),.CI(carry[38:38]),.CO(carry[39:39]),.S(DIFF[38:38]));
  FADDX1 U2_37(.A(A[37:37]),.B(n40),.CI(carry[37:37]),.CO(carry[38:38]),.S(DIFF[37:37]));
  FADDX1 U2_36(.A(A[36:36]),.B(n19),.CI(carry[36:36]),.CO(carry[37:37]),.S(DIFF[36:36]));
  FADDX1 U2_35(.A(A[35:35]),.B(n39),.CI(carry[35:35]),.CO(carry[36:36]),.S(DIFF[35:35]));
  FADDX1 U2_34(.A(A[34:34]),.B(n18),.CI(carry[34:34]),.CO(carry[35:35]),.S(DIFF[34:34]));
  FADDX1 U2_33(.A(A[33:33]),.B(n38),.CI(carry[33:33]),.CO(carry[34:34]),.S(DIFF[33:33]));
  FADDX1 U2_32(.A(A[32:32]),.B(n17),.CI(carry[32:32]),.CO(carry[33:33]),.S(DIFF[32:32]));
  FADDX1 U2_31(.A(A[31:31]),.B(n27),.CI(carry[31:31]),.CO(carry[32:32]),.S(DIFF[31:31]));
  FADDX1 U2_30(.A(A[30:30]),.B(n14),.CI(carry[30:30]),.CO(carry[31:31]),.S(DIFF[30:30]));
  FADDX1 U2_29(.A(A[29:29]),.B(n31),.CI(carry[29:29]),.CO(carry[30:30]),.S(DIFF[29:29]));
  FADDX1 U2_28(.A(A[28:28]),.B(n6),.CI(carry[28:28]),.CO(carry[29:29]),.S(DIFF[28:28]));
  FADDX1 U2_27(.A(A[27:27]),.B(n23),.CI(carry[27:27]),.CO(carry[28:28]),.S(DIFF[27:27]));
  FADDX1 U2_26(.A(A[26:26]),.B(n10),.CI(carry[26:26]),.CO(carry[27:27]),.S(DIFF[26:26]));
  FADDX1 U2_25(.A(A[25:25]),.B(n36),.CI(carry[25:25]),.CO(carry[26:26]),.S(DIFF[25:25]));
  FADDX1 U2_24(.A(A[24:24]),.B(n3),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n28),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n15),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n32),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n7),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n24),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n11),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n34),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n2),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n26),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n13),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n30),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n5),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n22),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n9),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n37),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n4),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n29),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n16),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n33),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n8),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n25),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n12),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n35),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_51(.IN1(A[51:51]),.IN2(n52),.IN3(carry[51:51]),.Q(DIFF[51:51]));
  INVX0 U1(.INP(B[32:32]),.ZN(n17));
  INVX0 U2(.INP(B[4:4]),.ZN(n8));
  INVX0 U3(.INP(B[48:48]),.ZN(n49));
  INVX0 U4(.INP(B[46:46]),.ZN(n47));
  INVX0 U5(.INP(B[44:44]),.ZN(n45));
  INVX0 U6(.INP(B[50:50]),.ZN(n51));
  INVX0 U7(.INP(B[42:42]),.ZN(n43));
  INVX0 U8(.INP(B[40:40]),.ZN(n21));
  INVX0 U9(.INP(B[38:38]),.ZN(n20));
  INVX0 U10(.INP(B[36:36]),.ZN(n19));
  INVX0 U11(.INP(B[34:34]),.ZN(n18));
  INVX0 U12(.INP(B[30:30]),.ZN(n14));
  INVX0 U13(.INP(B[2:2]),.ZN(n12));
  INVX0 U14(.INP(B[6:6]),.ZN(n16));
  INVX0 U15(.INP(B[8:8]),.ZN(n4));
  INVX0 U16(.INP(B[10:10]),.ZN(n9));
  INVX0 U17(.INP(B[12:12]),.ZN(n5));
  INVX0 U18(.INP(B[14:14]),.ZN(n13));
  INVX0 U19(.INP(B[16:16]),.ZN(n2));
  INVX0 U20(.INP(B[18:18]),.ZN(n11));
  INVX0 U21(.INP(B[20:20]),.ZN(n7));
  INVX0 U22(.INP(B[22:22]),.ZN(n15));
  INVX0 U23(.INP(B[24:24]),.ZN(n3));
  INVX0 U24(.INP(B[26:26]),.ZN(n10));
  INVX0 U25(.INP(B[28:28]),.ZN(n6));
  INVX0 U26(.INP(B[47:47]),.ZN(n48));
  INVX0 U27(.INP(B[49:49]),.ZN(n50));
  INVX0 U28(.INP(B[45:45]),.ZN(n46));
  INVX0 U29(.INP(B[43:43]),.ZN(n44));
  INVX0 U30(.INP(B[41:41]),.ZN(n42));
  INVX0 U31(.INP(B[39:39]),.ZN(n41));
  INVX0 U32(.INP(B[37:37]),.ZN(n40));
  INVX0 U33(.INP(B[35:35]),.ZN(n39));
  INVX0 U34(.INP(B[33:33]),.ZN(n38));
  INVX0 U35(.INP(B[31:31]),.ZN(n27));
  INVX0 U36(.INP(B[29:29]),.ZN(n31));
  INVX0 U37(.INP(B[3:3]),.ZN(n25));
  INVX0 U38(.INP(B[5:5]),.ZN(n33));
  INVX0 U39(.INP(B[7:7]),.ZN(n29));
  INVX0 U40(.INP(B[9:9]),.ZN(n37));
  INVX0 U41(.INP(B[11:11]),.ZN(n22));
  INVX0 U42(.INP(B[13:13]),.ZN(n30));
  INVX0 U43(.INP(B[15:15]),.ZN(n26));
  INVX0 U44(.INP(B[17:17]),.ZN(n34));
  INVX0 U45(.INP(B[19:19]),.ZN(n24));
  INVX0 U46(.INP(B[21:21]),.ZN(n32));
  INVX0 U47(.INP(B[23:23]),.ZN(n28));
  INVX0 U48(.INP(B[25:25]),.ZN(n36));
  INVX0 U49(.INP(B[27:27]),.ZN(n23));
  INVX0 U50(.INP(B[1:1]),.ZN(n35));
  NAND2X0 U51(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U52(.INP(A[0:0]),.ZN(n1));
  INVX0 U53(.INP(B[51:51]),.ZN(n52));
  XOR2X1 U54(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_1_inj (A,B,CI,SUM,CO);
input [25:0] A ;
input [25:0] B ;
output [25:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire [25:1] carry ;
// instances
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(carry[24:24]),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_23(.A(A[23:23]),.B(B[23:23]),.CI(carry[23:23]),.CO(carry[24:24]),.S(SUM[23:23]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(carry[22:22]),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_21(.A(A[21:21]),.B(B[21:21]),.CI(carry[21:21]),.CO(carry[22:22]),.S(SUM[21:21]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(carry[20:20]),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_19(.A(A[19:19]),.B(B[19:19]),.CI(carry[19:19]),.CO(carry[20:20]),.S(SUM[19:19]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(carry[18:18]),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_17(.A(A[17:17]),.B(B[17:17]),.CI(carry[17:17]),.CO(carry[18:18]),.S(SUM[17:17]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(carry[16:16]),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_15(.A(A[15:15]),.B(B[15:15]),.CI(carry[15:15]),.CO(carry[16:16]),.S(SUM[15:15]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(carry[14:14]),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_13(.A(A[13:13]),.B(B[13:13]),.CI(carry[13:13]),.CO(carry[14:14]),.S(SUM[13:13]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(carry[12:12]),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_11(.A(A[11:11]),.B(B[11:11]),.CI(carry[11:11]),.CO(carry[12:12]),.S(SUM[11:11]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(carry[10:10]),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_9(.A(A[9:9]),.B(B[9:9]),.CI(carry[9:9]),.CO(carry[10:10]),.S(SUM[9:9]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(carry[8:8]),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_7(.A(A[7:7]),.B(B[7:7]),.CI(carry[7:7]),.CO(carry[8:8]),.S(SUM[7:7]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(carry[6:6]),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_5(.A(A[5:5]),.B(B[5:5]),.CI(carry[5:5]),.CO(carry[6:6]),.S(SUM[5:5]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(carry[4:4]),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_3(.A(A[3:3]),.B(B[3:3]),.CI(carry[3:3]),.CO(carry[4:4]),.S(SUM[3:3]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(carry[2:2]),.CO(carry[3:3]),.S(SUM[2:2]));
  FADDX1 U1_1(.A(A[1:1]),.B(B[1:1]),.CI(n1),.CO(carry[2:2]),.S(SUM[1:1]));
  XOR3X1 U1_25(.IN1(A[25:25]),.IN2(B[25:25]),.IN3(carry[25:25]),.Q(SUM[25:25]));
  AND2X1 U1(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n1));
  XOR2X1 U2(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_2_inj (A,B,CI,DIFF,CO);
input [25:0] A ;
input [25:0] B ;
output [25:0] DIFF ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire [26:0] carry ;
// instances
  FADDX1 U2_24(.A(A[24:24]),.B(n3),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n4),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n5),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n6),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n7),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n8),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n9),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n10),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n11),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n12),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n13),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n14),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n15),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n16),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n17),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n18),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n19),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n20),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n21),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n22),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n23),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n24),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n25),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  FADDX1 U2_1(.A(A[1:1]),.B(n26),.CI(carry[1:1]),.CO(carry[2:2]),.S(DIFF[1:1]));
  XOR3X1 U2_25(.IN1(A[25:25]),.IN2(n2),.IN3(carry[25:25]),.Q(DIFF[25:25]));
  INVX0 U1(.INP(B[1:1]),.ZN(n26));
  NAND2X1 U2(.IN1(n1),.IN2(B[0:0]),.QN(carry[1:1]));
  INVX0 U3(.INP(A[0:0]),.ZN(n1));
  INVX0 U4(.INP(B[2:2]),.ZN(n25));
  INVX0 U5(.INP(B[3:3]),.ZN(n24));
  INVX0 U6(.INP(B[4:4]),.ZN(n23));
  INVX0 U7(.INP(B[5:5]),.ZN(n22));
  INVX0 U8(.INP(B[6:6]),.ZN(n21));
  INVX0 U9(.INP(B[7:7]),.ZN(n20));
  INVX0 U10(.INP(B[8:8]),.ZN(n19));
  INVX0 U11(.INP(B[9:9]),.ZN(n18));
  INVX0 U12(.INP(B[10:10]),.ZN(n17));
  INVX0 U13(.INP(B[11:11]),.ZN(n16));
  INVX0 U14(.INP(B[12:12]),.ZN(n15));
  INVX0 U15(.INP(B[13:13]),.ZN(n14));
  INVX0 U16(.INP(B[14:14]),.ZN(n13));
  INVX0 U17(.INP(B[15:15]),.ZN(n12));
  INVX0 U18(.INP(B[16:16]),.ZN(n11));
  INVX0 U19(.INP(B[17:17]),.ZN(n10));
  INVX0 U20(.INP(B[18:18]),.ZN(n9));
  INVX0 U21(.INP(B[19:19]),.ZN(n8));
  INVX0 U22(.INP(B[20:20]),.ZN(n7));
  INVX0 U23(.INP(B[21:21]),.ZN(n6));
  INVX0 U24(.INP(B[22:22]),.ZN(n5));
  INVX0 U25(.INP(B[23:23]),.ZN(n4));
  INVX0 U26(.INP(B[24:24]),.ZN(n3));
  INVX0 U27(.INP(B[25:25]),.ZN(n2));
  XOR2X1 U28(.IN1(B[0:0]),.IN2(A[0:0]),.Q(DIFF[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_2_inj (A,B,CI,SUM,CO);
input [51:0] A ;
input [51:0] B ;
output [51:0] SUM ;
input CI ;
output CO ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire [51:1] carry ;
// instances
  FADDX1 U1_50(.A(A[50:50]),.B(B[50:50]),.CI(n8),.CO(carry[51:51]),.S(SUM[50:50]));
  FADDX1 U1_48(.A(A[48:48]),.B(B[48:48]),.CI(n6),.CO(carry[49:49]),.S(SUM[48:48]));
  FADDX1 U1_46(.A(A[46:46]),.B(B[46:46]),.CI(n26),.CO(carry[47:47]),.S(SUM[46:46]));
  FADDX1 U1_44(.A(A[44:44]),.B(B[44:44]),.CI(n5),.CO(carry[45:45]),.S(SUM[44:44]));
  FADDX1 U1_42(.A(A[42:42]),.B(B[42:42]),.CI(n25),.CO(carry[43:43]),.S(SUM[42:42]));
  FADDX1 U1_40(.A(A[40:40]),.B(B[40:40]),.CI(n3),.CO(carry[41:41]),.S(SUM[40:40]));
  FADDX1 U1_38(.A(A[38:38]),.B(B[38:38]),.CI(n11),.CO(carry[39:39]),.S(SUM[38:38]));
  FADDX1 U1_36(.A(A[36:36]),.B(B[36:36]),.CI(n13),.CO(carry[37:37]),.S(SUM[36:36]));
  FADDX1 U1_34(.A(A[34:34]),.B(B[34:34]),.CI(n10),.CO(carry[35:35]),.S(SUM[34:34]));
  FADDX1 U1_32(.A(A[32:32]),.B(B[32:32]),.CI(n1),.CO(carry[33:33]),.S(SUM[32:32]));
  FADDX1 U1_30(.A(A[30:30]),.B(B[30:30]),.CI(n24),.CO(carry[31:31]),.S(SUM[30:30]));
  FADDX1 U1_28(.A(A[28:28]),.B(B[28:28]),.CI(n21),.CO(carry[29:29]),.S(SUM[28:28]));
  FADDX1 U1_26(.A(A[26:26]),.B(B[26:26]),.CI(n22),.CO(carry[27:27]),.S(SUM[26:26]));
  FADDX1 U1_24(.A(A[24:24]),.B(B[24:24]),.CI(n20),.CO(carry[25:25]),.S(SUM[24:24]));
  FADDX1 U1_22(.A(A[22:22]),.B(B[22:22]),.CI(n19),.CO(carry[23:23]),.S(SUM[22:22]));
  FADDX1 U1_20(.A(A[20:20]),.B(B[20:20]),.CI(n17),.CO(carry[21:21]),.S(SUM[20:20]));
  FADDX1 U1_18(.A(A[18:18]),.B(B[18:18]),.CI(n16),.CO(carry[19:19]),.S(SUM[18:18]));
  FADDX1 U1_16(.A(A[16:16]),.B(B[16:16]),.CI(n18),.CO(carry[17:17]),.S(SUM[16:16]));
  FADDX1 U1_14(.A(A[14:14]),.B(B[14:14]),.CI(n12),.CO(carry[15:15]),.S(SUM[14:14]));
  FADDX1 U1_12(.A(A[12:12]),.B(B[12:12]),.CI(n4),.CO(carry[13:13]),.S(SUM[12:12]));
  FADDX1 U1_10(.A(A[10:10]),.B(B[10:10]),.CI(n23),.CO(carry[11:11]),.S(SUM[10:10]));
  FADDX1 U1_8(.A(A[8:8]),.B(B[8:8]),.CI(n7),.CO(carry[9:9]),.S(SUM[8:8]));
  FADDX1 U1_6(.A(A[6:6]),.B(B[6:6]),.CI(n14),.CO(carry[7:7]),.S(SUM[6:6]));
  FADDX1 U1_4(.A(A[4:4]),.B(B[4:4]),.CI(n2),.CO(carry[5:5]),.S(SUM[4:4]));
  FADDX1 U1_2(.A(A[2:2]),.B(B[2:2]),.CI(n9),.CO(carry[3:3]),.S(SUM[2:2]));
  AND2X1 U1(.IN1(A[31:31]),.IN2(carry[31:31]),.Q(n1));
  AND2X1 U2(.IN1(A[3:3]),.IN2(carry[3:3]),.Q(n2));
  AND2X1 U3(.IN1(A[39:39]),.IN2(carry[39:39]),.Q(n3));
  AND2X1 U4(.IN1(A[11:11]),.IN2(carry[11:11]),.Q(n4));
  AND2X1 U5(.IN1(A[43:43]),.IN2(carry[43:43]),.Q(n5));
  AND2X1 U6(.IN1(A[47:47]),.IN2(carry[47:47]),.Q(n6));
  AND2X1 U7(.IN1(A[7:7]),.IN2(carry[7:7]),.Q(n7));
  AND2X1 U8(.IN1(A[49:49]),.IN2(carry[49:49]),.Q(n8));
  AND2X1 U9(.IN1(A[1:1]),.IN2(n15),.Q(n9));
  AND2X1 U10(.IN1(A[33:33]),.IN2(carry[33:33]),.Q(n10));
  AND2X1 U11(.IN1(A[37:37]),.IN2(carry[37:37]),.Q(n11));
  AND2X1 U12(.IN1(A[13:13]),.IN2(carry[13:13]),.Q(n12));
  AND2X1 U13(.IN1(A[35:35]),.IN2(carry[35:35]),.Q(n13));
  AND2X1 U14(.IN1(A[5:5]),.IN2(carry[5:5]),.Q(n14));
  AND2X1 U15(.IN1(A[0:0]),.IN2(B[0:0]),.Q(n15));
  AND2X1 U16(.IN1(A[17:17]),.IN2(carry[17:17]),.Q(n16));
  AND2X1 U17(.IN1(A[19:19]),.IN2(carry[19:19]),.Q(n17));
  AND2X1 U18(.IN1(A[15:15]),.IN2(carry[15:15]),.Q(n18));
  AND2X1 U19(.IN1(A[21:21]),.IN2(carry[21:21]),.Q(n19));
  AND2X1 U20(.IN1(A[23:23]),.IN2(carry[23:23]),.Q(n20));
  AND2X1 U21(.IN1(A[27:27]),.IN2(carry[27:27]),.Q(n21));
  AND2X1 U22(.IN1(A[25:25]),.IN2(carry[25:25]),.Q(n22));
  AND2X1 U23(.IN1(A[9:9]),.IN2(carry[9:9]),.Q(n23));
  AND2X1 U24(.IN1(A[29:29]),.IN2(carry[29:29]),.Q(n24));
  AND2X1 U25(.IN1(A[41:41]),.IN2(carry[41:41]),.Q(n25));
  AND2X1 U26(.IN1(A[45:45]),.IN2(carry[45:45]),.Q(n26));
  XOR2X1 U27(.IN1(A[51:51]),.IN2(carry[51:51]),.Q(SUM[51:51]));
  XOR2X1 U28(.IN1(A[49:49]),.IN2(carry[49:49]),.Q(SUM[49:49]));
  XOR2X1 U29(.IN1(A[47:47]),.IN2(carry[47:47]),.Q(SUM[47:47]));
  XOR2X1 U30(.IN1(A[45:45]),.IN2(carry[45:45]),.Q(SUM[45:45]));
  XOR2X1 U31(.IN1(A[43:43]),.IN2(carry[43:43]),.Q(SUM[43:43]));
  XOR2X1 U32(.IN1(A[41:41]),.IN2(carry[41:41]),.Q(SUM[41:41]));
  XOR2X1 U33(.IN1(A[39:39]),.IN2(carry[39:39]),.Q(SUM[39:39]));
  XOR2X1 U34(.IN1(A[37:37]),.IN2(carry[37:37]),.Q(SUM[37:37]));
  XOR2X1 U35(.IN1(A[35:35]),.IN2(carry[35:35]),.Q(SUM[35:35]));
  XOR2X1 U36(.IN1(A[33:33]),.IN2(carry[33:33]),.Q(SUM[33:33]));
  XOR2X1 U37(.IN1(A[31:31]),.IN2(carry[31:31]),.Q(SUM[31:31]));
  XOR2X1 U38(.IN1(A[29:29]),.IN2(carry[29:29]),.Q(SUM[29:29]));
  XOR2X1 U39(.IN1(A[27:27]),.IN2(carry[27:27]),.Q(SUM[27:27]));
  XOR2X1 U40(.IN1(A[25:25]),.IN2(carry[25:25]),.Q(SUM[25:25]));
  XOR2X1 U41(.IN1(A[23:23]),.IN2(carry[23:23]),.Q(SUM[23:23]));
  XOR2X1 U42(.IN1(A[21:21]),.IN2(carry[21:21]),.Q(SUM[21:21]));
  XOR2X1 U43(.IN1(A[19:19]),.IN2(carry[19:19]),.Q(SUM[19:19]));
  XOR2X1 U44(.IN1(A[17:17]),.IN2(carry[17:17]),.Q(SUM[17:17]));
  XOR2X1 U45(.IN1(A[15:15]),.IN2(carry[15:15]),.Q(SUM[15:15]));
  XOR2X1 U46(.IN1(A[13:13]),.IN2(carry[13:13]),.Q(SUM[13:13]));
  XOR2X1 U47(.IN1(A[11:11]),.IN2(carry[11:11]),.Q(SUM[11:11]));
  XOR2X1 U48(.IN1(A[9:9]),.IN2(carry[9:9]),.Q(SUM[9:9]));
  XOR2X1 U49(.IN1(A[7:7]),.IN2(carry[7:7]),.Q(SUM[7:7]));
  XOR2X1 U50(.IN1(A[5:5]),.IN2(carry[5:5]),.Q(SUM[5:5]));
  XOR2X1 U51(.IN1(A[3:3]),.IN2(carry[3:3]),.Q(SUM[3:3]));
  XOR2X1 U52(.IN1(A[1:1]),.IN2(n15),.Q(SUM[1:1]));
  XOR2X1 U53(.IN1(A[0:0]),.IN2(B[0:0]),.Q(SUM[0:0]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp6_0_inj (A,B,TC,LT,GT,EQ,LE,GE,NE);
input [51:0] A ;
input [51:0] B ;
input TC ;
output LT ;
output GT ;
output EQ ;
output LE ;
output GE ;
output NE ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n129 ;
wire n130 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
// instances
  INVX0 U1(.INP(n58),.ZN(LT));
  INVX0 U2(.INP(n90),.ZN(n4));
  INVX0 U3(.INP(n91),.ZN(n3));
  INVX0 U4(.INP(n106),.ZN(n2));
  INVX0 U5(.INP(A[3:3]),.ZN(n5));
  INVX0 U6(.INP(B[15:15]),.ZN(n44));
  INVX0 U7(.INP(B[7:7]),.ZN(n52));
  INVX0 U8(.INP(B[9:9]),.ZN(n50));
  INVX0 U9(.INP(B[11:11]),.ZN(n48));
  INVX0 U10(.INP(B[13:13]),.ZN(n46));
  INVX0 U11(.INP(B[17:17]),.ZN(n42));
  INVX0 U12(.INP(B[19:19]),.ZN(n40));
  INVX0 U13(.INP(B[21:21]),.ZN(n38));
  INVX0 U14(.INP(B[23:23]),.ZN(n36));
  INVX0 U15(.INP(B[25:25]),.ZN(n34));
  INVX0 U16(.INP(B[0:0]),.ZN(n57));
  INVX0 U17(.INP(B[4:4]),.ZN(n55));
  INVX0 U18(.INP(B[5:5]),.ZN(n54));
  INVX0 U19(.INP(A[2:2]),.ZN(n6));
  INVX0 U20(.INP(B[6:6]),.ZN(n53));
  INVX0 U21(.INP(B[16:16]),.ZN(n43));
  INVX0 U22(.INP(B[8:8]),.ZN(n51));
  INVX0 U23(.INP(B[10:10]),.ZN(n49));
  INVX0 U24(.INP(B[12:12]),.ZN(n47));
  INVX0 U25(.INP(B[14:14]),.ZN(n45));
  INVX0 U26(.INP(B[20:20]),.ZN(n39));
  INVX0 U27(.INP(B[18:18]),.ZN(n41));
  INVX0 U28(.INP(B[22:22]),.ZN(n37));
  INVX0 U29(.INP(B[26:26]),.ZN(n33));
  INVX0 U30(.INP(B[24:24]),.ZN(n35));
  INVX0 U31(.INP(B[27:27]),.ZN(n32));
  INVX0 U32(.INP(B[29:29]),.ZN(n30));
  INVX0 U33(.INP(B[28:28]),.ZN(n31));
  INVX0 U34(.INP(B[30:30]),.ZN(n29));
  INVX0 U35(.INP(A[1:1]),.ZN(n7));
  INVX0 U36(.INP(B[31:31]),.ZN(n28));
  INVX0 U37(.INP(B[33:33]),.ZN(n26));
  INVX0 U38(.INP(B[35:35]),.ZN(n24));
  INVX0 U39(.INP(B[37:37]),.ZN(n22));
  INVX0 U40(.INP(B[39:39]),.ZN(n20));
  INVX0 U41(.INP(B[41:41]),.ZN(n18));
  INVX0 U42(.INP(B[43:43]),.ZN(n16));
  INVX0 U43(.INP(B[45:45]),.ZN(n14));
  INVX0 U44(.INP(B[34:34]),.ZN(n25));
  INVX0 U45(.INP(B[32:32]),.ZN(n27));
  INVX0 U46(.INP(B[36:36]),.ZN(n23));
  INVX0 U47(.INP(B[40:40]),.ZN(n19));
  INVX0 U48(.INP(B[38:38]),.ZN(n21));
  INVX0 U49(.INP(B[42:42]),.ZN(n17));
  INVX0 U50(.INP(B[44:44]),.ZN(n15));
  INVX0 U51(.INP(B[46:46]),.ZN(n13));
  INVX0 U52(.INP(B[50:50]),.ZN(n9));
  INVX0 U53(.INP(B[47:47]),.ZN(n12));
  INVX0 U54(.INP(B[49:49]),.ZN(n10));
  INVX0 U55(.INP(B[48:48]),.ZN(n11));
  INVX0 U56(.INP(B[51:51]),.ZN(n8));
  INVX0 U57(.INP(B[1:1]),.ZN(n56));
  NOR2X0 U58(.IN1(n59),.IN2(n60),.QN(EQ));
  NAND4X0 U59(.IN1(n61),.IN2(n62),.IN3(n63),.IN4(n64),.QN(n60));
  AND4X1 U60(.IN1(n65),.IN2(n66),.IN3(n67),.IN4(n68),.Q(n64));
  AND4X1 U61(.IN1(n69),.IN2(n70),.IN3(n71),.IN4(n72),.Q(n65));
  AND4X1 U62(.IN1(n73),.IN2(n74),.IN3(n75),.IN4(n76),.Q(n63));
  AND3X1 U63(.IN1(n77),.IN2(n78),.IN3(n79),.Q(n73));
  AND4X1 U64(.IN1(n80),.IN2(n81),.IN3(n82),.IN4(n83),.Q(n62));
  AND4X1 U65(.IN1(n84),.IN2(n85),.IN3(n86),.IN4(n87),.Q(n80));
  NOR4X0 U66(.IN1(n88),.IN2(n89),.IN3(n3),.IN4(n4),.QN(n61));
  OA22X1 U67(.IN1(n92),.IN2(n56),.IN3(A[1:1]),.IN4(n92),.Q(n89));
  AND2X1 U68(.IN1(A[0:0]),.IN2(n57),.Q(n92));
  NAND3X0 U69(.IN1(n93),.IN2(n94),.IN3(n95),.QN(n88));
  NAND4X0 U70(.IN1(n96),.IN2(n97),.IN3(n98),.IN4(n99),.QN(n59));
  AND4X1 U71(.IN1(n100),.IN2(n101),.IN3(n102),.IN4(n103),.Q(n99));
  AND4X1 U72(.IN1(n104),.IN2(n105),.IN3(n106),.IN4(n58),.Q(n100));
  OA22X1 U73(.IN1(A[51:51]),.IN2(n8),.IN3(n2),.IN4(n107),.Q(n58));
  OA22X1 U74(.IN1(A[50:50]),.IN2(n9),.IN3(n108),.IN4(n109),.Q(n107));
  NAND2X0 U75(.IN1(n90),.IN2(n91),.QN(n109));
  NAND2X0 U76(.IN1(A[50:50]),.IN2(n9),.QN(n91));
  NAND2X0 U77(.IN1(A[49:49]),.IN2(n10),.QN(n90));
  OA222X1 U78(.IN1(A[49:49]),.IN2(n10),.IN3(A[48:48]),.IN4(n11),.IN5(n110),.IN6(n111),.Q(n108));
  NAND2X0 U79(.IN1(n95),.IN2(n93),.QN(n111));
  NAND2X0 U80(.IN1(A[47:47]),.IN2(n12),.QN(n93));
  NAND2X0 U81(.IN1(A[48:48]),.IN2(n11),.QN(n95));
  OA222X1 U82(.IN1(A[47:47]),.IN2(n12),.IN3(A[46:46]),.IN4(n13),.IN5(n112),.IN6(n113),.Q(n110));
  NAND2X0 U83(.IN1(n94),.IN2(n81),.QN(n113));
  NAND2X0 U84(.IN1(A[45:45]),.IN2(n14),.QN(n81));
  NAND2X0 U85(.IN1(A[46:46]),.IN2(n13),.QN(n94));
  OA222X1 U86(.IN1(A[45:45]),.IN2(n14),.IN3(A[44:44]),.IN4(n15),.IN5(n114),.IN6(n115),.Q(n112));
  NAND2X0 U87(.IN1(n83),.IN2(n82),.QN(n115));
  NAND2X0 U88(.IN1(A[43:43]),.IN2(n16),.QN(n82));
  NAND2X0 U89(.IN1(A[44:44]),.IN2(n15),.QN(n83));
  OA222X1 U90(.IN1(A[43:43]),.IN2(n16),.IN3(A[42:42]),.IN4(n17),.IN5(n116),.IN6(n117),.Q(n114));
  NAND2X0 U91(.IN1(n84),.IN2(n85),.QN(n117));
  NAND2X0 U92(.IN1(A[41:41]),.IN2(n18),.QN(n85));
  NAND2X0 U93(.IN1(A[42:42]),.IN2(n17),.QN(n84));
  OA222X1 U94(.IN1(A[41:41]),.IN2(n18),.IN3(A[40:40]),.IN4(n19),.IN5(n118),.IN6(n119),.Q(n116));
  NAND2X0 U95(.IN1(n86),.IN2(n87),.QN(n119));
  NAND2X0 U96(.IN1(A[39:39]),.IN2(n20),.QN(n87));
  NAND2X0 U97(.IN1(A[40:40]),.IN2(n19),.QN(n86));
  OA222X1 U98(.IN1(A[39:39]),.IN2(n20),.IN3(A[38:38]),.IN4(n21),.IN5(n120),.IN6(n121),.Q(n118));
  NAND2X0 U99(.IN1(n74),.IN2(n76),.QN(n121));
  NAND2X0 U100(.IN1(A[37:37]),.IN2(n22),.QN(n76));
  NAND2X0 U101(.IN1(A[38:38]),.IN2(n21),.QN(n74));
  OA222X1 U102(.IN1(A[37:37]),.IN2(n22),.IN3(A[36:36]),.IN4(n23),.IN5(n122),.IN6(n123),.Q(n120));
  NAND2X0 U103(.IN1(n75),.IN2(n79),.QN(n123));
  NAND2X0 U104(.IN1(A[35:35]),.IN2(n24),.QN(n79));
  NAND2X0 U105(.IN1(A[36:36]),.IN2(n23),.QN(n75));
  OA222X1 U106(.IN1(A[35:35]),.IN2(n24),.IN3(A[34:34]),.IN4(n25),.IN5(n124),.IN6(n125),.Q(n122));
  NAND2X0 U107(.IN1(n77),.IN2(n78),.QN(n125));
  NAND2X0 U108(.IN1(A[33:33]),.IN2(n26),.QN(n78));
  NAND2X0 U109(.IN1(A[34:34]),.IN2(n25),.QN(n77));
  OA222X1 U110(.IN1(A[33:33]),.IN2(n26),.IN3(A[32:32]),.IN4(n27),.IN5(n126),.IN6(n127),.Q(n124));
  NAND2X0 U111(.IN1(n66),.IN2(n68),.QN(n127));
  NAND2X0 U112(.IN1(A[31:31]),.IN2(n28),.QN(n68));
  NAND2X0 U113(.IN1(A[32:32]),.IN2(n27),.QN(n66));
  OA222X1 U114(.IN1(A[31:31]),.IN2(n28),.IN3(A[30:30]),.IN4(n29),.IN5(n128),.IN6(n129),.Q(n126));
  NAND2X0 U115(.IN1(n67),.IN2(n69),.QN(n129));
  NAND2X0 U116(.IN1(A[29:29]),.IN2(n30),.QN(n69));
  NAND2X0 U117(.IN1(A[30:30]),.IN2(n29),.QN(n67));
  OA222X1 U118(.IN1(A[29:29]),.IN2(n30),.IN3(A[28:28]),.IN4(n31),.IN5(n130),.IN6(n131),.Q(n128));
  NAND2X0 U119(.IN1(n70),.IN2(n71),.QN(n131));
  NAND2X0 U120(.IN1(A[27:27]),.IN2(n32),.QN(n71));
  NAND2X0 U121(.IN1(A[28:28]),.IN2(n31),.QN(n70));
  OA222X1 U122(.IN1(A[27:27]),.IN2(n32),.IN3(A[26:26]),.IN4(n33),.IN5(n132),.IN6(n133),.Q(n130));
  NAND2X0 U123(.IN1(n72),.IN2(n134),.QN(n133));
  NAND2X0 U124(.IN1(A[26:26]),.IN2(n33),.QN(n72));
  OA222X1 U125(.IN1(A[25:25]),.IN2(n34),.IN3(A[24:24]),.IN4(n35),.IN5(n135),.IN6(n136),.Q(n132));
  NAND2X0 U126(.IN1(n137),.IN2(n138),.QN(n136));
  OA222X1 U127(.IN1(A[23:23]),.IN2(n36),.IN3(A[22:22]),.IN4(n37),.IN5(n139),.IN6(n140),.Q(n135));
  NAND2X0 U128(.IN1(n141),.IN2(n142),.QN(n140));
  OA222X1 U129(.IN1(A[21:21]),.IN2(n38),.IN3(A[20:20]),.IN4(n39),.IN5(n143),.IN6(n144),.Q(n139));
  NAND2X0 U130(.IN1(n145),.IN2(n146),.QN(n144));
  OA222X1 U131(.IN1(A[19:19]),.IN2(n40),.IN3(A[18:18]),.IN4(n41),.IN5(n147),.IN6(n148),.Q(n143));
  NAND2X0 U132(.IN1(n149),.IN2(n150),.QN(n148));
  OA222X1 U133(.IN1(A[17:17]),.IN2(n42),.IN3(A[16:16]),.IN4(n43),.IN5(n151),.IN6(n152),.Q(n147));
  NAND2X0 U134(.IN1(n153),.IN2(n154),.QN(n152));
  OA222X1 U135(.IN1(A[15:15]),.IN2(n44),.IN3(A[14:14]),.IN4(n45),.IN5(n155),.IN6(n156),.Q(n151));
  NAND2X0 U136(.IN1(n157),.IN2(n158),.QN(n156));
  OA222X1 U137(.IN1(A[13:13]),.IN2(n46),.IN3(A[12:12]),.IN4(n47),.IN5(n159),.IN6(n160),.Q(n155));
  NAND2X0 U138(.IN1(n161),.IN2(n162),.QN(n160));
  OA222X1 U139(.IN1(A[11:11]),.IN2(n48),.IN3(A[10:10]),.IN4(n49),.IN5(n163),.IN6(n164),.Q(n159));
  NAND2X0 U140(.IN1(n165),.IN2(n166),.QN(n164));
  OA222X1 U141(.IN1(A[9:9]),.IN2(n50),.IN3(A[8:8]),.IN4(n51),.IN5(n167),.IN6(n168),.Q(n163));
  NAND2X0 U142(.IN1(n169),.IN2(n170),.QN(n168));
  OA222X1 U143(.IN1(A[7:7]),.IN2(n52),.IN3(A[6:6]),.IN4(n53),.IN5(n171),.IN6(n172),.Q(n167));
  NAND2X0 U144(.IN1(n101),.IN2(n103),.QN(n172));
  NAND2X0 U145(.IN1(A[5:5]),.IN2(n54),.QN(n103));
  NAND2X0 U146(.IN1(A[6:6]),.IN2(n53),.QN(n101));
  OA221X1 U147(.IN1(A[5:5]),.IN2(n54),.IN3(A[4:4]),.IN4(n55),.IN5(n173),.Q(n171));
  NAND3X0 U148(.IN1(n102),.IN2(n104),.IN3(n174),.QN(n173));
  AO221X1 U149(.IN1(B[2:2]),.IN2(n6),.IN3(B[3:3]),.IN4(n5),.IN5(n175),.Q(n174));
  OA221X1 U150(.IN1(n176),.IN2(n7),.IN3(B[1:1]),.IN4(n177),.IN5(n105),.Q(n175));
  AND2X1 U151(.IN1(n7),.IN2(n176),.Q(n177));
  NOR2X0 U152(.IN1(n57),.IN2(A[0:0]),.QN(n176));
  NAND2X0 U153(.IN1(A[4:4]),.IN2(n55),.QN(n102));
  NAND2X0 U154(.IN1(A[51:51]),.IN2(n8),.QN(n106));
  OR2X1 U155(.IN1(n6),.IN2(B[2:2]),.Q(n105));
  OR2X1 U156(.IN1(n5),.IN2(B[3:3]),.Q(n104));
  AND4X1 U157(.IN1(n178),.IN2(n161),.IN3(n165),.IN4(n162),.Q(n98));
  NAND2X0 U158(.IN1(A[11:11]),.IN2(n48),.QN(n162));
  NAND2X0 U159(.IN1(A[10:10]),.IN2(n49),.QN(n165));
  NAND2X0 U160(.IN1(A[12:12]),.IN2(n47),.QN(n161));
  AND3X1 U161(.IN1(n169),.IN2(n170),.IN3(n166),.Q(n178));
  NAND2X0 U162(.IN1(A[9:9]),.IN2(n50),.QN(n166));
  NAND2X0 U163(.IN1(A[7:7]),.IN2(n52),.QN(n170));
  NAND2X0 U164(.IN1(A[8:8]),.IN2(n51),.QN(n169));
  AND4X1 U165(.IN1(n179),.IN2(n146),.IN3(n150),.IN4(n149),.Q(n97));
  NAND2X0 U166(.IN1(A[18:18]),.IN2(n41),.QN(n149));
  NAND2X0 U167(.IN1(A[17:17]),.IN2(n42),.QN(n150));
  NAND2X0 U168(.IN1(A[19:19]),.IN2(n40),.QN(n146));
  AND4X1 U169(.IN1(n153),.IN2(n154),.IN3(n157),.IN4(n158),.Q(n179));
  NAND2X0 U170(.IN1(A[13:13]),.IN2(n46),.QN(n158));
  NAND2X0 U171(.IN1(A[14:14]),.IN2(n45),.QN(n157));
  NAND2X0 U172(.IN1(A[15:15]),.IN2(n44),.QN(n154));
  NAND2X0 U173(.IN1(A[16:16]),.IN2(n43),.QN(n153));
  AND4X1 U174(.IN1(n180),.IN2(n134),.IN3(n138),.IN4(n137),.Q(n96));
  NAND2X0 U175(.IN1(A[24:24]),.IN2(n35),.QN(n137));
  NAND2X0 U176(.IN1(A[23:23]),.IN2(n36),.QN(n138));
  NAND2X0 U177(.IN1(A[25:25]),.IN2(n34),.QN(n134));
  AND3X1 U178(.IN1(n142),.IN2(n145),.IN3(n141),.Q(n180));
  NAND2X0 U179(.IN1(A[22:22]),.IN2(n37),.QN(n141));
  NAND2X0 U180(.IN1(A[20:20]),.IN2(n39),.QN(n145));
  NAND2X0 U181(.IN1(A[21:21]),.IN2(n38),.QN(n142));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_3_inj (A,B,CI,DIFF,CO);
input [51:0] A ;
input [51:0] B ;
output [51:0] DIFF ;
input CI ;
output CO ;
wire \A[0]  ;
wire n1 ;
wire n2 ;
wire n3 ;
wire n4 ;
wire n5 ;
wire n6 ;
wire n7 ;
wire n8 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire [52:0] carry ;
// instances
  FADDX1 U2_26(.A(A[26:26]),.B(n50),.CI(carry[26:26]),.CO(carry[27:27]),.S(DIFF[26:26]));
  FADDX1 U2_25(.A(A[25:25]),.B(n51),.CI(carry[25:25]),.CO(carry[26:26]),.S(DIFF[25:25]));
  FADDX1 U2_24(.A(A[24:24]),.B(n52),.CI(carry[24:24]),.CO(carry[25:25]),.S(DIFF[24:24]));
  FADDX1 U2_23(.A(A[23:23]),.B(n53),.CI(carry[23:23]),.CO(carry[24:24]),.S(DIFF[23:23]));
  FADDX1 U2_22(.A(A[22:22]),.B(n54),.CI(carry[22:22]),.CO(carry[23:23]),.S(DIFF[22:22]));
  FADDX1 U2_21(.A(A[21:21]),.B(n55),.CI(carry[21:21]),.CO(carry[22:22]),.S(DIFF[21:21]));
  FADDX1 U2_20(.A(A[20:20]),.B(n56),.CI(carry[20:20]),.CO(carry[21:21]),.S(DIFF[20:20]));
  FADDX1 U2_19(.A(A[19:19]),.B(n57),.CI(carry[19:19]),.CO(carry[20:20]),.S(DIFF[19:19]));
  FADDX1 U2_18(.A(A[18:18]),.B(n58),.CI(carry[18:18]),.CO(carry[19:19]),.S(DIFF[18:18]));
  FADDX1 U2_17(.A(A[17:17]),.B(n59),.CI(carry[17:17]),.CO(carry[18:18]),.S(DIFF[17:17]));
  FADDX1 U2_16(.A(A[16:16]),.B(n60),.CI(carry[16:16]),.CO(carry[17:17]),.S(DIFF[16:16]));
  FADDX1 U2_15(.A(A[15:15]),.B(n61),.CI(carry[15:15]),.CO(carry[16:16]),.S(DIFF[15:15]));
  FADDX1 U2_14(.A(A[14:14]),.B(n62),.CI(carry[14:14]),.CO(carry[15:15]),.S(DIFF[14:14]));
  FADDX1 U2_13(.A(A[13:13]),.B(n63),.CI(carry[13:13]),.CO(carry[14:14]),.S(DIFF[13:13]));
  FADDX1 U2_12(.A(A[12:12]),.B(n64),.CI(carry[12:12]),.CO(carry[13:13]),.S(DIFF[12:12]));
  FADDX1 U2_11(.A(A[11:11]),.B(n65),.CI(carry[11:11]),.CO(carry[12:12]),.S(DIFF[11:11]));
  FADDX1 U2_10(.A(A[10:10]),.B(n66),.CI(carry[10:10]),.CO(carry[11:11]),.S(DIFF[10:10]));
  FADDX1 U2_9(.A(A[9:9]),.B(n67),.CI(carry[9:9]),.CO(carry[10:10]),.S(DIFF[9:9]));
  FADDX1 U2_8(.A(A[8:8]),.B(n68),.CI(carry[8:8]),.CO(carry[9:9]),.S(DIFF[8:8]));
  FADDX1 U2_7(.A(A[7:7]),.B(n69),.CI(carry[7:7]),.CO(carry[8:8]),.S(DIFF[7:7]));
  FADDX1 U2_6(.A(A[6:6]),.B(n70),.CI(carry[6:6]),.CO(carry[7:7]),.S(DIFF[6:6]));
  FADDX1 U2_5(.A(A[5:5]),.B(n71),.CI(carry[5:5]),.CO(carry[6:6]),.S(DIFF[5:5]));
  FADDX1 U2_4(.A(A[4:4]),.B(n72),.CI(carry[4:4]),.CO(carry[5:5]),.S(DIFF[4:4]));
  FADDX1 U2_3(.A(A[3:3]),.B(n73),.CI(carry[3:3]),.CO(carry[4:4]),.S(DIFF[3:3]));
  FADDX1 U2_2(.A(A[2:2]),.B(n74),.CI(carry[2:2]),.CO(carry[3:3]),.S(DIFF[2:2]));
  INVX0 U1(.INP(A[36:36]),.ZN(n27));
  INVX0 U2(.INP(A[31:31]),.ZN(n32));
  INVX0 U3(.INP(A[44:44]),.ZN(n44));
  INVX0 U4(.INP(A[35:35]),.ZN(n28));
  INVX0 U5(.INP(A[47:47]),.ZN(n41));
  INVX0 U6(.INP(A[30:30]),.ZN(n33));
  INVX0 U7(.INP(A[41:41]),.ZN(n47));
  INVX0 U8(.INP(A[34:34]),.ZN(n29));
  INVX0 U9(.INP(A[29:29]),.ZN(n34));
  INVX0 U10(.INP(A[40:40]),.ZN(n48));
  INVX0 U11(.INP(A[45:45]),.ZN(n43));
  INVX0 U12(.INP(A[38:38]),.ZN(n25));
  INVX0 U13(.INP(A[32:32]),.ZN(n31));
  INVX0 U14(.INP(A[28:28]),.ZN(n35));
  INVX0 U15(.INP(A[48:48]),.ZN(n40));
  INVX0 U16(.INP(A[42:42]),.ZN(n46));
  INVX0 U17(.INP(A[27:27]),.ZN(n36));
  INVX0 U18(.INP(A[49:49]),.ZN(n39));
  INVX0 U19(.INP(A[43:43]),.ZN(n45));
  INVX0 U20(.INP(A[39:39]),.ZN(n49));
  INVX0 U21(.INP(A[33:33]),.ZN(n30));
  INVX0 U22(.INP(carry[27:27]),.ZN(n37));
  INVX0 U23(.INP(B[2:2]),.ZN(n74));
  NAND2X0 U24(.IN1(n24),.IN2(B[1:1]),.QN(carry[2:2]));
  INVX0 U25(.INP(A[1:1]),.ZN(n24));
  INVX0 U26(.INP(B[3:3]),.ZN(n73));
  INVX0 U27(.INP(B[19:19]),.ZN(n57));
  INVX0 U28(.INP(B[20:20]),.ZN(n56));
  INVX0 U29(.INP(B[21:21]),.ZN(n55));
  INVX0 U30(.INP(B[22:22]),.ZN(n54));
  INVX0 U31(.INP(B[23:23]),.ZN(n53));
  INVX0 U32(.INP(B[18:18]),.ZN(n58));
  INVX0 U33(.INP(B[24:24]),.ZN(n52));
  INVX0 U34(.INP(B[25:25]),.ZN(n51));
  INVX0 U35(.INP(B[17:17]),.ZN(n59));
  INVX0 U36(.INP(B[16:16]),.ZN(n60));
  INVX0 U37(.INP(B[15:15]),.ZN(n61));
  INVX0 U38(.INP(B[14:14]),.ZN(n62));
  INVX0 U39(.INP(B[13:13]),.ZN(n63));
  INVX0 U40(.INP(B[12:12]),.ZN(n64));
  INVX0 U41(.INP(B[11:11]),.ZN(n65));
  INVX0 U42(.INP(B[10:10]),.ZN(n66));
  INVX0 U43(.INP(B[9:9]),.ZN(n67));
  INVX0 U44(.INP(B[5:5]),.ZN(n71));
  INVX0 U45(.INP(B[6:6]),.ZN(n70));
  INVX0 U46(.INP(B[8:8]),.ZN(n68));
  INVX0 U47(.INP(B[7:7]),.ZN(n69));
  INVX0 U48(.INP(B[4:4]),.ZN(n72));
  INVX0 U49(.INP(B[26:26]),.ZN(n50));
  AND2X1 U50(.IN1(n36),.IN2(n37),.Q(n1));
  AND2X1 U51(.IN1(n35),.IN2(n1),.Q(n2));
  AND2X1 U52(.IN1(n34),.IN2(n2),.Q(n3));
  AND2X1 U53(.IN1(n33),.IN2(n3),.Q(n4));
  AND2X1 U54(.IN1(n31),.IN2(n23),.Q(n5));
  AND2X1 U55(.IN1(n30),.IN2(n5),.Q(n6));
  AND2X1 U56(.IN1(n29),.IN2(n6),.Q(n7));
  AND2X1 U57(.IN1(n28),.IN2(n7),.Q(n8));
  AND2X1 U58(.IN1(n27),.IN2(n8),.Q(n9));
  AND2X1 U59(.IN1(n26),.IN2(n9),.Q(n10));
  AND2X1 U60(.IN1(n25),.IN2(n10),.Q(n11));
  AND2X1 U61(.IN1(n49),.IN2(n11),.Q(n12));
  AND2X1 U62(.IN1(n48),.IN2(n12),.Q(n13));
  AND2X1 U63(.IN1(n47),.IN2(n13),.Q(n14));
  AND2X1 U64(.IN1(n46),.IN2(n14),.Q(n15));
  AND2X1 U65(.IN1(n45),.IN2(n15),.Q(n16));
  AND2X1 U66(.IN1(n44),.IN2(n16),.Q(n17));
  AND2X1 U67(.IN1(n43),.IN2(n17),.Q(n18));
  AND2X1 U68(.IN1(n42),.IN2(n18),.Q(n19));
  AND2X1 U69(.IN1(n41),.IN2(n19),.Q(n20));
  AND2X1 U70(.IN1(n40),.IN2(n20),.Q(n21));
  AND2X1 U71(.IN1(n39),.IN2(n21),.Q(n22));
  XNOR2X1 U72(.IN1(carry[51:51]),.IN2(A[51:51]),.Q(DIFF[51:51]));
  AND2X1 U73(.IN1(n32),.IN2(n4),.Q(n23));
  NAND2X0 U74(.IN1(n38),.IN2(n22),.QN(carry[51:51]));
  INVX0 U75(.INP(A[50:50]),.ZN(n38));
  XOR2X1 U76(.IN1(B[1:1]),.IN2(A[1:1]),.Q(DIFF[1:1]));
  XOR2X1 U77(.IN1(n10),.IN2(A[38:38]),.Q(DIFF[38:38]));
  XOR2X1 U78(.IN1(n9),.IN2(A[37:37]),.Q(DIFF[37:37]));
  INVX1 U79(.INP(A[37:37]),.ZN(n26));
  XOR2X1 U80(.IN1(n8),.IN2(A[36:36]),.Q(DIFF[36:36]));
  XOR2X1 U81(.IN1(n7),.IN2(A[35:35]),.Q(DIFF[35:35]));
  XOR2X1 U82(.IN1(n6),.IN2(A[34:34]),.Q(DIFF[34:34]));
  XOR2X1 U83(.IN1(n5),.IN2(A[33:33]),.Q(DIFF[33:33]));
  XOR2X1 U84(.IN1(n23),.IN2(A[32:32]),.Q(DIFF[32:32]));
  XOR2X1 U85(.IN1(n4),.IN2(A[31:31]),.Q(DIFF[31:31]));
  XOR2X1 U86(.IN1(n3),.IN2(A[30:30]),.Q(DIFF[30:30]));
  XOR2X1 U87(.IN1(n2),.IN2(A[29:29]),.Q(DIFF[29:29]));
  XOR2X1 U88(.IN1(n1),.IN2(A[28:28]),.Q(DIFF[28:28]));
  XOR2X1 U89(.IN1(n37),.IN2(A[27:27]),.Q(DIFF[27:27]));
  XOR2X1 U90(.IN1(n22),.IN2(A[50:50]),.Q(DIFF[50:50]));
  XOR2X1 U91(.IN1(n21),.IN2(A[49:49]),.Q(DIFF[49:49]));
  XOR2X1 U92(.IN1(n20),.IN2(A[48:48]),.Q(DIFF[48:48]));
  XOR2X1 U93(.IN1(n19),.IN2(A[47:47]),.Q(DIFF[47:47]));
  XOR2X1 U94(.IN1(n18),.IN2(A[46:46]),.Q(DIFF[46:46]));
  INVX1 U95(.INP(A[46:46]),.ZN(n42));
  XOR2X1 U96(.IN1(n17),.IN2(A[45:45]),.Q(DIFF[45:45]));
  XOR2X1 U97(.IN1(n16),.IN2(A[44:44]),.Q(DIFF[44:44]));
  XOR2X1 U98(.IN1(n15),.IN2(A[43:43]),.Q(DIFF[43:43]));
  XOR2X1 U99(.IN1(n14),.IN2(A[42:42]),.Q(DIFF[42:42]));
  XOR2X1 U100(.IN1(n13),.IN2(A[41:41]),.Q(DIFF[41:41]));
  XOR2X1 U101(.IN1(n12),.IN2(A[40:40]),.Q(DIFF[40:40]));
  XOR2X1 U102(.IN1(n11),.IN2(A[39:39]),.Q(DIFF[39:39]));
assign DIFF[0:0]=\A[0] ;
assign \A[0] =A[0:0];
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_inc_0_inj (A,SUM);
input [51:0] A ;
output [51:0] SUM ;
wire [51:2] carry ;
// instances
  HADDX1 U1_1_50(.A0(A[50:50]),.B0(carry[50:50]),.C1(carry[51:51]),.SO(SUM[50:50]));
  HADDX1 U1_1_49(.A0(A[49:49]),.B0(carry[49:49]),.C1(carry[50:50]),.SO(SUM[49:49]));
  HADDX1 U1_1_48(.A0(A[48:48]),.B0(carry[48:48]),.C1(carry[49:49]),.SO(SUM[48:48]));
  HADDX1 U1_1_47(.A0(A[47:47]),.B0(carry[47:47]),.C1(carry[48:48]),.SO(SUM[47:47]));
  HADDX1 U1_1_46(.A0(A[46:46]),.B0(carry[46:46]),.C1(carry[47:47]),.SO(SUM[46:46]));
  HADDX1 U1_1_45(.A0(A[45:45]),.B0(carry[45:45]),.C1(carry[46:46]),.SO(SUM[45:45]));
  HADDX1 U1_1_44(.A0(A[44:44]),.B0(carry[44:44]),.C1(carry[45:45]),.SO(SUM[44:44]));
  HADDX1 U1_1_43(.A0(A[43:43]),.B0(carry[43:43]),.C1(carry[44:44]),.SO(SUM[43:43]));
  HADDX1 U1_1_42(.A0(A[42:42]),.B0(carry[42:42]),.C1(carry[43:43]),.SO(SUM[42:42]));
  HADDX1 U1_1_41(.A0(A[41:41]),.B0(carry[41:41]),.C1(carry[42:42]),.SO(SUM[41:41]));
  HADDX1 U1_1_40(.A0(A[40:40]),.B0(carry[40:40]),.C1(carry[41:41]),.SO(SUM[40:40]));
  HADDX1 U1_1_39(.A0(A[39:39]),.B0(carry[39:39]),.C1(carry[40:40]),.SO(SUM[39:39]));
  HADDX1 U1_1_38(.A0(A[38:38]),.B0(carry[38:38]),.C1(carry[39:39]),.SO(SUM[38:38]));
  HADDX1 U1_1_37(.A0(A[37:37]),.B0(carry[37:37]),.C1(carry[38:38]),.SO(SUM[37:37]));
  HADDX1 U1_1_36(.A0(A[36:36]),.B0(carry[36:36]),.C1(carry[37:37]),.SO(SUM[36:36]));
  HADDX1 U1_1_35(.A0(A[35:35]),.B0(carry[35:35]),.C1(carry[36:36]),.SO(SUM[35:35]));
  HADDX1 U1_1_34(.A0(A[34:34]),.B0(carry[34:34]),.C1(carry[35:35]),.SO(SUM[34:34]));
  HADDX1 U1_1_33(.A0(A[33:33]),.B0(carry[33:33]),.C1(carry[34:34]),.SO(SUM[33:33]));
  HADDX1 U1_1_32(.A0(A[32:32]),.B0(carry[32:32]),.C1(carry[33:33]),.SO(SUM[32:32]));
  HADDX1 U1_1_31(.A0(A[31:31]),.B0(carry[31:31]),.C1(carry[32:32]),.SO(SUM[31:31]));
  HADDX1 U1_1_30(.A0(A[30:30]),.B0(carry[30:30]),.C1(carry[31:31]),.SO(SUM[30:30]));
  HADDX1 U1_1_29(.A0(A[29:29]),.B0(carry[29:29]),.C1(carry[30:30]),.SO(SUM[29:29]));
  HADDX1 U1_1_28(.A0(A[28:28]),.B0(carry[28:28]),.C1(carry[29:29]),.SO(SUM[28:28]));
  HADDX1 U1_1_27(.A0(A[27:27]),.B0(carry[27:27]),.C1(carry[28:28]),.SO(SUM[27:27]));
  HADDX1 U1_1_26(.A0(A[26:26]),.B0(carry[26:26]),.C1(carry[27:27]),.SO(SUM[26:26]));
  HADDX1 U1_1_25(.A0(A[25:25]),.B0(carry[25:25]),.C1(carry[26:26]),.SO(SUM[25:25]));
  HADDX1 U1_1_24(.A0(A[24:24]),.B0(carry[24:24]),.C1(carry[25:25]),.SO(SUM[24:24]));
  HADDX1 U1_1_23(.A0(A[23:23]),.B0(carry[23:23]),.C1(carry[24:24]),.SO(SUM[23:23]));
  HADDX1 U1_1_22(.A0(A[22:22]),.B0(carry[22:22]),.C1(carry[23:23]),.SO(SUM[22:22]));
  HADDX1 U1_1_21(.A0(A[21:21]),.B0(carry[21:21]),.C1(carry[22:22]),.SO(SUM[21:21]));
  HADDX1 U1_1_20(.A0(A[20:20]),.B0(carry[20:20]),.C1(carry[21:21]),.SO(SUM[20:20]));
  HADDX1 U1_1_19(.A0(A[19:19]),.B0(carry[19:19]),.C1(carry[20:20]),.SO(SUM[19:19]));
  HADDX1 U1_1_18(.A0(A[18:18]),.B0(carry[18:18]),.C1(carry[19:19]),.SO(SUM[18:18]));
  HADDX1 U1_1_17(.A0(A[17:17]),.B0(carry[17:17]),.C1(carry[18:18]),.SO(SUM[17:17]));
  HADDX1 U1_1_16(.A0(A[16:16]),.B0(carry[16:16]),.C1(carry[17:17]),.SO(SUM[16:16]));
  HADDX1 U1_1_15(.A0(A[15:15]),.B0(carry[15:15]),.C1(carry[16:16]),.SO(SUM[15:15]));
  HADDX1 U1_1_14(.A0(A[14:14]),.B0(carry[14:14]),.C1(carry[15:15]),.SO(SUM[14:14]));
  HADDX1 U1_1_13(.A0(A[13:13]),.B0(carry[13:13]),.C1(carry[14:14]),.SO(SUM[13:13]));
  HADDX1 U1_1_12(.A0(A[12:12]),.B0(carry[12:12]),.C1(carry[13:13]),.SO(SUM[12:12]));
  HADDX1 U1_1_11(.A0(A[11:11]),.B0(carry[11:11]),.C1(carry[12:12]),.SO(SUM[11:11]));
  HADDX1 U1_1_10(.A0(A[10:10]),.B0(carry[10:10]),.C1(carry[11:11]),.SO(SUM[10:10]));
  HADDX1 U1_1_9(.A0(A[9:9]),.B0(carry[9:9]),.C1(carry[10:10]),.SO(SUM[9:9]));
  HADDX1 U1_1_8(.A0(A[8:8]),.B0(carry[8:8]),.C1(carry[9:9]),.SO(SUM[8:8]));
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[51:51]),.IN2(A[51:51]),.Q(SUM[51:51]));
endmodule
module sqrt_RD_WIDTH52_SQ_WIDTH26_inj (clk_i,rad_i,start_i,ready_o,sqr_o,ine_o);
input [51:0] rad_i ;
output [25:0] sqr_o ;
input clk_i ;
input start_i ;
output ready_o ;
output ine_o ;
wire s_ine_o ;
wire s_ready_o ;
wire s_state ;
wire \s_count[4]  ;
wire \s_count[3]  ;
wire \s_count[2]  ;
wire \s_count[1]  ;
wire \s_count[0]  ;
wire N11 ;
wire N12 ;
wire N13 ;
wire N14 ;
wire N31 ;
wire N32 ;
wire N33 ;
wire N34 ;
wire N35 ;
wire N36 ;
wire N37 ;
wire N38 ;
wire N39 ;
wire N40 ;
wire N41 ;
wire N42 ;
wire N43 ;
wire N44 ;
wire N45 ;
wire N46 ;
wire N47 ;
wire N48 ;
wire N49 ;
wire N50 ;
wire N51 ;
wire N52 ;
wire N53 ;
wire N54 ;
wire N55 ;
wire N56 ;
wire N57 ;
wire N58 ;
wire N59 ;
wire N86 ;
wire N88 ;
wire N90 ;
wire N92 ;
wire N94 ;
wire N96 ;
wire N98 ;
wire N100 ;
wire N102 ;
wire N104 ;
wire N106 ;
wire N108 ;
wire N110 ;
wire N112 ;
wire N114 ;
wire N116 ;
wire N118 ;
wire N120 ;
wire N122 ;
wire N124 ;
wire N126 ;
wire N128 ;
wire N130 ;
wire N132 ;
wire N134 ;
wire N136 ;
wire N137 ;
wire N138 ;
wire N139 ;
wire N140 ;
wire N142 ;
wire N306 ;
wire N309 ;
wire N310 ;
wire N311 ;
wire N312 ;
wire N313 ;
wire N314 ;
wire N315 ;
wire N316 ;
wire N317 ;
wire N318 ;
wire N319 ;
wire N320 ;
wire N321 ;
wire N322 ;
wire N323 ;
wire N324 ;
wire N325 ;
wire N326 ;
wire N327 ;
wire N328 ;
wire N329 ;
wire N330 ;
wire N331 ;
wire N332 ;
wire N333 ;
wire N334 ;
wire N414 ;
wire N415 ;
wire N416 ;
wire N417 ;
wire N418 ;
wire N419 ;
wire N420 ;
wire N421 ;
wire N422 ;
wire N423 ;
wire N424 ;
wire N425 ;
wire N426 ;
wire N427 ;
wire N428 ;
wire N429 ;
wire N430 ;
wire N431 ;
wire N432 ;
wire N433 ;
wire N434 ;
wire N435 ;
wire N436 ;
wire N437 ;
wire N438 ;
wire N439 ;
wire N440 ;
wire N441 ;
wire N442 ;
wire N443 ;
wire N444 ;
wire N445 ;
wire N446 ;
wire N447 ;
wire N448 ;
wire N449 ;
wire N450 ;
wire N451 ;
wire N452 ;
wire N453 ;
wire N454 ;
wire N455 ;
wire N456 ;
wire N457 ;
wire N458 ;
wire N459 ;
wire N460 ;
wire N461 ;
wire N462 ;
wire N463 ;
wire N464 ;
wire N465 ;
wire N466 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n49 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n90 ;
wire n91 ;
wire n92 ;
wire n93 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n128 ;
wire n129 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire n277 ;
wire n278 ;
wire n279 ;
wire n280 ;
wire n281 ;
wire n282 ;
wire n283 ;
wire n284 ;
wire n285 ;
wire n286 ;
wire n287 ;
wire n288 ;
wire n289 ;
wire n290 ;
wire n291 ;
wire n292 ;
wire n293 ;
wire n294 ;
wire n295 ;
wire n296 ;
wire n297 ;
wire n298 ;
wire n299 ;
wire n300 ;
wire n301 ;
wire n302 ;
wire n303 ;
wire n304 ;
wire n305 ;
wire n306 ;
wire n307 ;
wire n308 ;
wire n309 ;
wire n310 ;
wire n311 ;
wire n312 ;
wire n313 ;
wire n314 ;
wire n315 ;
wire n316 ;
wire n317 ;
wire n318 ;
wire n319 ;
wire n320 ;
wire n321 ;
wire n322 ;
wire n323 ;
wire n324 ;
wire n325 ;
wire n326 ;
wire n327 ;
wire n328 ;
wire n329 ;
wire n330 ;
wire n331 ;
wire n332 ;
wire n333 ;
wire n334 ;
wire n335 ;
wire n336 ;
wire n337 ;
wire n338 ;
wire n339 ;
wire n340 ;
wire n341 ;
wire n342 ;
wire n343 ;
wire n344 ;
wire n345 ;
wire n346 ;
wire n347 ;
wire n348 ;
wire n349 ;
wire n350 ;
wire n351 ;
wire n352 ;
wire n353 ;
wire n354 ;
wire n355 ;
wire n356 ;
wire n357 ;
wire n358 ;
wire n359 ;
wire n360 ;
wire n361 ;
wire n362 ;
wire n363 ;
wire n364 ;
wire n365 ;
wire n366 ;
wire n367 ;
wire n368 ;
wire n369 ;
wire n370 ;
wire n371 ;
wire n372 ;
wire n373 ;
wire n374 ;
wire n375 ;
wire n376 ;
wire n377 ;
wire n378 ;
wire n379 ;
wire n380 ;
wire n381 ;
wire n382 ;
wire n383 ;
wire n384 ;
wire n385 ;
wire n386 ;
wire n387 ;
wire n388 ;
wire n389 ;
wire n390 ;
wire n391 ;
wire n392 ;
wire n393 ;
wire n394 ;
wire n395 ;
wire n396 ;
wire n397 ;
wire n398 ;
wire n399 ;
wire n400 ;
wire N413 ;
wire N412 ;
wire N411 ;
wire N410 ;
wire N409 ;
wire N408 ;
wire N407 ;
wire N406 ;
wire N405 ;
wire N404 ;
wire N403 ;
wire N402 ;
wire N401 ;
wire N400 ;
wire N399 ;
wire N398 ;
wire N397 ;
wire N396 ;
wire N395 ;
wire N394 ;
wire N393 ;
wire N392 ;
wire N391 ;
wire N390 ;
wire N389 ;
wire N388 ;
wire N387 ;
wire N386 ;
wire N385 ;
wire N384 ;
wire N383 ;
wire N382 ;
wire N381 ;
wire N380 ;
wire N379 ;
wire N378 ;
wire N377 ;
wire N376 ;
wire N375 ;
wire N374 ;
wire N373 ;
wire N372 ;
wire N371 ;
wire N370 ;
wire N369 ;
wire N368 ;
wire N367 ;
wire N366 ;
wire N365 ;
wire N364 ;
wire N363 ;
wire N362 ;
wire n1 ;
wire n2 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n117 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n130 ;
wire n401 ;
wire n402 ;
wire n403 ;
wire n404 ;
wire n405 ;
wire n406 ;
wire n407 ;
wire n408 ;
wire n409 ;
wire n410 ;
wire n411 ;
wire n412 ;
wire n413 ;
wire n414 ;
wire n415 ;
wire n416 ;
wire n417 ;
wire n418 ;
wire n419 ;
wire n420 ;
wire n421 ;
wire n422 ;
wire n423 ;
wire n424 ;
wire n425 ;
wire n426 ;
wire n427 ;
wire n428 ;
wire n429 ;
wire n430 ;
wire n431 ;
wire n432 ;
wire n433 ;
wire n434 ;
wire n435 ;
wire n436 ;
wire n437 ;
wire n438 ;
wire n439 ;
wire n440 ;
wire n441 ;
wire n442 ;
wire n443 ;
wire n444 ;
wire n445 ;
wire n446 ;
wire n447 ;
wire n448 ;
wire n449 ;
wire n450 ;
wire n451 ;
wire n452 ;
wire n453 ;
wire n454 ;
wire n455 ;
wire n456 ;
wire n457 ;
wire n458 ;
wire n459 ;
wire n460 ;
wire n461 ;
wire n462 ;
wire n463 ;
wire n464 ;
wire n465 ;
wire n466 ;
wire n467 ;
wire n468 ;
wire n469 ;
wire n470 ;
wire n471 ;
wire n472 ;
wire n473 ;
wire n474 ;
wire n475 ;
wire n478 ;
wire n479 ;
wire n480 ;
wire n481 ;
wire n482 ;
wire n483 ;
wire n484 ;
wire n485 ;
wire n486 ;
wire n487 ;
wire n488 ;
wire n489 ;
wire n490 ;
wire n491 ;
wire n492 ;
wire n493 ;
wire n494 ;
wire n495 ;
wire n496 ;
wire n497 ;
wire n498 ;
wire n499 ;
wire n500 ;
wire n501 ;
wire n502 ;
wire n503 ;
wire n504 ;
wire n505 ;
wire n506 ;
wire n507 ;
wire n508 ;
wire n509 ;
wire n510 ;
wire n511 ;
wire n512 ;
wire n513 ;
wire n514 ;
wire n515 ;
wire n516 ;
wire n517 ;
wire n518 ;
wire n519 ;
wire n520 ;
wire n521 ;
wire n522 ;
wire n523 ;
wire n524 ;
wire n525 ;
wire n526 ;
wire n527 ;
wire n528 ;
wire n529 ;
wire n530 ;
wire n531 ;
wire n532 ;
wire n533 ;
wire n534 ;
wire n535 ;
wire n536 ;
wire n537 ;
wire n538 ;
wire n539 ;
wire n540 ;
wire n541 ;
wire n542 ;
wire n543 ;
wire n544 ;
wire n545 ;
wire n546 ;
wire n547 ;
wire n548 ;
wire n549 ;
wire n550 ;
wire n551 ;
wire n552 ;
wire n553 ;
wire n554 ;
wire n555 ;
wire n556 ;
wire n557 ;
wire n558 ;
wire n559 ;
wire n560 ;
wire n561 ;
wire n562 ;
wire n563 ;
wire n564 ;
wire n565 ;
wire n566 ;
wire n567 ;
wire n568 ;
wire n569 ;
wire n570 ;
wire n571 ;
wire n572 ;
wire n573 ;
wire n574 ;
wire n575 ;
wire n576 ;
wire n577 ;
wire n578 ;
wire n579 ;
wire n580 ;
wire n581 ;
wire n582 ;
wire n583 ;
wire n584 ;
wire n585 ;
wire n586 ;
wire n587 ;
wire n588 ;
wire n589 ;
wire n590 ;
wire n591 ;
wire n592 ;
wire n593 ;
wire n594 ;
wire n595 ;
wire n596 ;
wire n597 ;
wire n598 ;
wire n599 ;
wire n600 ;
wire n601 ;
wire n602 ;
wire n603 ;
wire n604 ;
wire n605 ;
wire n606 ;
wire n607 ;
wire n608 ;
wire n609 ;
wire n610 ;
wire n611 ;
wire n612 ;
wire n613 ;
wire n614 ;
wire n615 ;
wire n616 ;
wire n617 ;
wire [51:0] s_rad_i ;
wire [25:0] s_sqr_o ;
wire [51:0] b ;
wire [51:0] b_2 ;
wire [4:0] c ;
wire [51:0] r0_2 ;
wire [51:0] s_op1 ;
wire [51:0] r0 ;
wire [51:0] s_op2 ;
wire [25:0] s_sum1a ;
wire [25:0] s_sum2a ;
wire [51:0] s_sum1b ;
wire [51:0] s_sum2b ;
wire [50:0] r1 ;
wire [51:0] r1_2 ;
// instances
  DFFX1 desc1955(.D(rad_i[51:51]),.CLK(clk_i),.Q(s_rad_i[51:51]));
  DFFX1 desc1956(.D(rad_i[50:50]),.CLK(clk_i),.Q(s_rad_i[50:50]));
  DFFX1 desc1957(.D(rad_i[49:49]),.CLK(clk_i),.Q(s_rad_i[49:49]));
  DFFX1 desc1958(.D(rad_i[48:48]),.CLK(clk_i),.Q(s_rad_i[48:48]));
  DFFX1 desc1959(.D(rad_i[47:47]),.CLK(clk_i),.Q(s_rad_i[47:47]),.QN(n168));
  DFFX1 desc1960(.D(rad_i[46:46]),.CLK(clk_i),.Q(s_rad_i[46:46]));
  DFFX1 desc1961(.D(rad_i[45:45]),.CLK(clk_i),.Q(s_rad_i[45:45]));
  DFFX1 desc1962(.D(rad_i[44:44]),.CLK(clk_i),.Q(s_rad_i[44:44]));
  DFFX1 desc1963(.D(rad_i[43:43]),.CLK(clk_i),.Q(s_rad_i[43:43]));
  DFFX1 desc1964(.D(rad_i[42:42]),.CLK(clk_i),.Q(s_rad_i[42:42]),.QN(n169));
  DFFX1 desc1965(.D(rad_i[41:41]),.CLK(clk_i),.Q(s_rad_i[41:41]));
  DFFX1 desc1966(.D(rad_i[40:40]),.CLK(clk_i),.Q(s_rad_i[40:40]));
  DFFX1 desc1967(.D(rad_i[39:39]),.CLK(clk_i),.Q(s_rad_i[39:39]),.QN(n163));
  DFFX1 desc1968(.D(rad_i[38:38]),.CLK(clk_i),.Q(s_rad_i[38:38]),.QN(n179));
  DFFX1 desc1969(.D(rad_i[37:37]),.CLK(clk_i),.Q(s_rad_i[37:37]),.QN(n177));
  DFFX1 desc1970(.D(rad_i[36:36]),.CLK(clk_i),.Q(s_rad_i[36:36]),.QN(n178));
  DFFX1 desc1971(.D(rad_i[35:35]),.CLK(clk_i),.Q(s_rad_i[35:35]),.QN(n164));
  DFFX1 desc1972(.D(rad_i[34:34]),.CLK(clk_i),.Q(s_rad_i[34:34]));
  DFFX1 desc1973(.D(rad_i[33:33]),.CLK(clk_i),.Q(s_rad_i[33:33]),.QN(n165));
  DFFX1 desc1974(.D(rad_i[32:32]),.CLK(clk_i),.Q(s_rad_i[32:32]),.QN(n180));
  DFFX1 desc1975(.D(rad_i[31:31]),.CLK(clk_i),.Q(s_rad_i[31:31]),.QN(n182));
  DFFX1 desc1976(.D(rad_i[30:30]),.CLK(clk_i),.Q(s_rad_i[30:30]),.QN(n181));
  DFFX1 desc1977(.D(rad_i[29:29]),.CLK(clk_i),.Q(s_rad_i[29:29]),.QN(n166));
  DFFX1 desc1978(.D(rad_i[28:28]),.CLK(clk_i),.Q(s_rad_i[28:28]),.QN(n167));
  DFFX1 desc1979(.D(rad_i[27:27]),.CLK(clk_i),.Q(s_rad_i[27:27]),.QN(n190));
  DFFX1 desc1980(.D(rad_i[26:26]),.CLK(clk_i),.Q(s_rad_i[26:26]),.QN(n189));
  DFFX1 desc1981(.D(rad_i[25:25]),.CLK(clk_i),.Q(s_rad_i[25:25]));
  DFFX1 desc1982(.D(rad_i[24:24]),.CLK(clk_i),.Q(s_rad_i[24:24]));
  DFFX1 desc1983(.D(rad_i[23:23]),.CLK(clk_i),.Q(s_rad_i[23:23]));
  DFFX1 desc1984(.D(rad_i[22:22]),.CLK(clk_i),.Q(s_rad_i[22:22]));
  DFFX1 desc1985(.D(rad_i[21:21]),.CLK(clk_i),.Q(s_rad_i[21:21]));
  DFFX1 desc1986(.D(rad_i[20:20]),.CLK(clk_i),.Q(s_rad_i[20:20]),.QN(n175));
  DFFX1 desc1987(.D(rad_i[19:19]),.CLK(clk_i),.Q(s_rad_i[19:19]));
  DFFX1 desc1988(.D(rad_i[18:18]),.CLK(clk_i),.Q(s_rad_i[18:18]));
  DFFX1 desc1989(.D(rad_i[17:17]),.CLK(clk_i),.Q(s_rad_i[17:17]),.QN(n184));
  DFFX1 desc1990(.D(rad_i[16:16]),.CLK(clk_i),.Q(s_rad_i[16:16]));
  DFFX1 desc1991(.D(rad_i[15:15]),.CLK(clk_i),.Q(s_rad_i[15:15]),.QN(n176));
  DFFX1 desc1992(.D(rad_i[14:14]),.CLK(clk_i),.Q(s_rad_i[14:14]));
  DFFX1 desc1993(.D(rad_i[13:13]),.CLK(clk_i),.Q(s_rad_i[13:13]));
  DFFX1 desc1994(.D(rad_i[12:12]),.CLK(clk_i),.Q(s_rad_i[12:12]),.QN(n185));
  DFFX1 desc1995(.D(rad_i[11:11]),.CLK(clk_i),.Q(s_rad_i[11:11]));
  DFFX1 desc1996(.D(rad_i[10:10]),.CLK(clk_i),.Q(s_rad_i[10:10]),.QN(n188));
  DFFX1 desc1997(.D(rad_i[9:9]),.CLK(clk_i),.Q(s_rad_i[9:9]),.QN(n172));
  DFFX1 desc1998(.D(rad_i[8:8]),.CLK(clk_i),.Q(s_rad_i[8:8]),.QN(n171));
  DFFX1 desc1999(.D(rad_i[7:7]),.CLK(clk_i),.Q(s_rad_i[7:7]),.QN(n170));
  DFFX1 desc2000(.D(rad_i[6:6]),.CLK(clk_i),.Q(s_rad_i[6:6]),.QN(n187));
  DFFX1 desc2001(.D(rad_i[5:5]),.CLK(clk_i),.Q(s_rad_i[5:5]),.QN(n186));
  DFFX1 desc2002(.D(rad_i[4:4]),.CLK(clk_i),.Q(s_rad_i[4:4]),.QN(n183));
  DFFX1 desc2003(.D(rad_i[3:3]),.CLK(clk_i),.Q(s_rad_i[3:3]));
  DFFX1 desc2004(.D(rad_i[2:2]),.CLK(clk_i),.Q(s_rad_i[2:2]),.QN(n173));
  DFFX1 desc2005(.D(rad_i[1:1]),.CLK(clk_i),.Q(s_rad_i[1:1]),.QN(n174));
  DFFX1 desc2006(.D(rad_i[0:0]),.CLK(clk_i),.Q(s_rad_i[0:0]));
  DFFX1 s_start_i_reg(.D(start_i),.CLK(clk_i),.QN(n1));
  DFFX1 desc2007(.D(n400),.CLK(clk_i),.Q(\s_count[0] ),.QN(n16));
  DFFX1 s_state_reg(.D(n398),.CLK(clk_i),.Q(s_state));
  DFFX1 s_ready_o_reg(.D(n397),.CLK(clk_i),.Q(s_ready_o));
  DFFX1 ready_o_reg(.D(s_ready_o),.CLK(clk_i),.Q(ready_o));
  DFFX1 desc2008(.D(n399),.CLK(clk_i),.Q(\s_count[4] ));
  DFFX1 desc2009(.D(n396),.CLK(clk_i),.Q(\s_count[1] ));
  DFFX1 desc2010(.D(n395),.CLK(clk_i),.Q(\s_count[2] ));
  DFFX1 desc2011(.D(n394),.CLK(clk_i),.Q(\s_count[3] ));
  DFFX1 desc2012(.D(N136),.CLK(clk_i),.Q(c[0:0]),.QN(n17));
  DFFX1 desc2013(.D(N137),.CLK(clk_i),.Q(c[1:1]),.QN(n2));
  DFFX1 desc2014(.D(N138),.CLK(clk_i),.Q(c[2:2]),.QN(n13));
  DFFX1 desc2015(.D(n424),.CLK(clk_i),.Q(b[25:25]),.QN(n203));
  DFFX1 desc2016(.D(N59),.CLK(clk_i),.Q(b[24:24]),.QN(n202));
  DFFX1 desc2017(.D(N58),.CLK(clk_i),.Q(b[23:23]),.QN(n201));
  DFFX1 desc2018(.D(N57),.CLK(clk_i),.Q(b[22:22]),.QN(n200));
  DFFX1 desc2019(.D(N56),.CLK(clk_i),.Q(b[21:21]),.QN(n199));
  DFFX1 desc2020(.D(N55),.CLK(clk_i),.Q(b[20:20]),.QN(n198));
  DFFX1 desc2021(.D(N54),.CLK(clk_i),.Q(b[19:19]),.QN(n197));
  DFFX1 desc2022(.D(N53),.CLK(clk_i),.Q(b[18:18]),.QN(n196));
  DFFX1 desc2023(.D(N52),.CLK(clk_i),.Q(b[17:17]),.QN(n195));
  DFFX1 desc2024(.D(N51),.CLK(clk_i),.Q(b[16:16]),.QN(n194));
  DFFX1 desc2025(.D(N50),.CLK(clk_i),.Q(b[15:15]),.QN(n193));
  DFFX1 desc2026(.D(N49),.CLK(clk_i),.Q(b[14:14]),.QN(n192));
  DFFX1 desc2027(.D(N48),.CLK(clk_i),.Q(b[13:13]),.QN(n191));
  DFFX1 desc2028(.D(N47),.CLK(clk_i),.Q(b[12:12]),.QN(n162));
  DFFX1 desc2029(.D(N46),.CLK(clk_i),.Q(b[11:11]),.QN(n161));
  DFFX1 desc2030(.D(N45),.CLK(clk_i),.Q(b[10:10]),.QN(n160));
  DFFX1 desc2031(.D(N44),.CLK(clk_i),.Q(b[9:9]),.QN(n159));
  DFFX1 desc2032(.D(N43),.CLK(clk_i),.Q(b[8:8]),.QN(n158));
  DFFX1 desc2033(.D(N42),.CLK(clk_i),.Q(b[7:7]),.QN(n157));
  DFFX1 desc2034(.D(N41),.CLK(clk_i),.Q(b[6:6]),.QN(n156));
  DFFX1 desc2035(.D(N40),.CLK(clk_i),.Q(b[5:5]),.QN(n155));
  DFFX1 desc2036(.D(N39),.CLK(clk_i),.Q(b[4:4]),.QN(n154));
  DFFX1 desc2037(.D(N38),.CLK(clk_i),.Q(b[3:3]),.QN(n153));
  DFFX1 desc2038(.D(N37),.CLK(clk_i),.Q(b[2:2]),.QN(n152));
  DFFX1 desc2039(.D(N36),.CLK(clk_i),.Q(b[1:1]),.QN(n151));
  DFFX1 desc2040(.D(N35),.CLK(clk_i),.Q(b[0:0]));
  DFFX1 desc2041(.D(n423),.CLK(clk_i),.Q(b_2[50:50]),.QN(n150));
  DFFX1 desc2042(.D(N134),.CLK(clk_i),.Q(b_2[48:48]),.QN(n149));
  DFFX1 desc2043(.D(N132),.CLK(clk_i),.Q(b_2[46:46]),.QN(n148));
  DFFX1 desc2044(.D(N130),.CLK(clk_i),.Q(b_2[44:44]),.QN(n147));
  DFFX1 desc2045(.D(N128),.CLK(clk_i),.Q(b_2[42:42]),.QN(n146));
  DFFX1 desc2046(.D(N126),.CLK(clk_i),.Q(b_2[40:40]),.QN(n145));
  DFFX1 desc2047(.D(N124),.CLK(clk_i),.Q(b_2[38:38]),.QN(n144));
  DFFX1 desc2048(.D(N122),.CLK(clk_i),.Q(b_2[36:36]),.QN(n143));
  DFFX1 desc2049(.D(N120),.CLK(clk_i),.Q(b_2[34:34]),.QN(n142));
  DFFX1 desc2050(.D(N118),.CLK(clk_i),.Q(b_2[32:32]),.QN(n141));
  DFFX1 desc2051(.D(N116),.CLK(clk_i),.Q(b_2[30:30]),.QN(n140));
  DFFX1 desc2052(.D(N114),.CLK(clk_i),.Q(b_2[28:28]),.QN(n139));
  DFFX1 desc2053(.D(N112),.CLK(clk_i),.Q(b_2[26:26]),.QN(n138));
  DFFX1 desc2054(.D(N110),.CLK(clk_i),.Q(b_2[24:24]),.QN(n137));
  DFFX1 desc2055(.D(N108),.CLK(clk_i),.Q(b_2[22:22]),.QN(n136));
  DFFX1 desc2056(.D(N106),.CLK(clk_i),.Q(b_2[20:20]),.QN(n135));
  DFFX1 desc2057(.D(N104),.CLK(clk_i),.Q(b_2[18:18]),.QN(n134));
  DFFX1 desc2058(.D(N102),.CLK(clk_i),.Q(b_2[16:16]),.QN(n133));
  DFFX1 desc2059(.D(N100),.CLK(clk_i),.Q(b_2[14:14]),.QN(n210));
  DFFX1 desc2060(.D(N98),.CLK(clk_i),.Q(b_2[12:12]),.QN(n209));
  DFFX1 desc2061(.D(N96),.CLK(clk_i),.Q(b_2[10:10]),.QN(n208));
  DFFX1 desc2062(.D(N94),.CLK(clk_i),.Q(b_2[8:8]),.QN(n207));
  DFFX1 desc2063(.D(N92),.CLK(clk_i),.Q(b_2[6:6]),.QN(n206));
  DFFX1 desc2064(.D(N90),.CLK(clk_i),.Q(b_2[4:4]),.QN(n205));
  DFFX1 desc2065(.D(N88),.CLK(clk_i),.Q(b_2[2:2]),.QN(n204));
  DFFX1 desc2066(.D(N86),.CLK(clk_i),.Q(b_2[0:0]));
  DFFX1 desc2067(.D(n393),.CLK(clk_i),.Q(r0_2[0:0]));
  DFFX1 desc2068(.D(n366),.CLK(clk_i),.Q(r0[0:0]));
  DFFX1 desc2069(.D(n341),.CLK(clk_i),.Q(r0[25:25]));
  DFFX1 desc2070(.D(n365),.CLK(clk_i),.Q(r0[1:1]));
  DFFX1 desc2071(.D(n364),.CLK(clk_i),.Q(r0[2:2]));
  DFFX1 desc2072(.D(n363),.CLK(clk_i),.Q(r0[3:3]));
  DFFX1 desc2073(.D(n362),.CLK(clk_i),.Q(r0[4:4]));
  DFFX1 desc2074(.D(n361),.CLK(clk_i),.Q(r0[5:5]));
  DFFX1 desc2075(.D(n360),.CLK(clk_i),.Q(r0[6:6]));
  DFFX1 desc2076(.D(n359),.CLK(clk_i),.Q(r0[7:7]));
  DFFX1 desc2077(.D(n358),.CLK(clk_i),.Q(r0[8:8]));
  DFFX1 desc2078(.D(n357),.CLK(clk_i),.Q(r0[9:9]));
  DFFX1 desc2079(.D(n356),.CLK(clk_i),.Q(r0[10:10]));
  DFFX1 desc2080(.D(n355),.CLK(clk_i),.Q(r0[11:11]));
  DFFX1 desc2081(.D(n354),.CLK(clk_i),.Q(r0[12:12]));
  DFFX1 desc2082(.D(n353),.CLK(clk_i),.Q(r0[13:13]));
  DFFX1 desc2083(.D(n352),.CLK(clk_i),.Q(r0[14:14]));
  DFFX1 desc2084(.D(n351),.CLK(clk_i),.Q(r0[15:15]));
  DFFX1 desc2085(.D(n350),.CLK(clk_i),.Q(r0[16:16]));
  DFFX1 desc2086(.D(n349),.CLK(clk_i),.Q(r0[17:17]));
  DFFX1 desc2087(.D(n348),.CLK(clk_i),.Q(r0[18:18]));
  DFFX1 desc2088(.D(n347),.CLK(clk_i),.Q(r0[19:19]));
  DFFX1 desc2089(.D(n346),.CLK(clk_i),.Q(r0[20:20]));
  DFFX1 desc2090(.D(n345),.CLK(clk_i),.Q(r0[21:21]));
  DFFX1 desc2091(.D(n344),.CLK(clk_i),.Q(r0[22:22]));
  DFFX1 desc2092(.D(n343),.CLK(clk_i),.Q(r0[23:23]));
  DFFX1 desc2093(.D(n342),.CLK(clk_i),.Q(r0[24:24]));
  DFFX1 desc2094(.D(n290),.CLK(clk_i),.Q(r0_2[51:51]));
  DFFX1 desc2095(.D(n340),.CLK(clk_i),.Q(r0_2[1:1]));
  DFFX1 desc2096(.D(n339),.CLK(clk_i),.Q(r0_2[2:2]));
  DFFX1 desc2097(.D(n338),.CLK(clk_i),.Q(r0_2[3:3]));
  DFFX1 desc2098(.D(n337),.CLK(clk_i),.Q(r0_2[4:4]));
  DFFX1 desc2099(.D(n336),.CLK(clk_i),.Q(r0_2[5:5]));
  DFFX1 desc2100(.D(n335),.CLK(clk_i),.Q(r0_2[6:6]));
  DFFX1 desc2101(.D(n334),.CLK(clk_i),.Q(r0_2[7:7]));
  DFFX1 desc2102(.D(n333),.CLK(clk_i),.Q(r0_2[8:8]));
  DFFX1 desc2103(.D(n332),.CLK(clk_i),.Q(r0_2[9:9]));
  DFFX1 desc2104(.D(n331),.CLK(clk_i),.Q(r0_2[10:10]));
  DFFX1 desc2105(.D(n330),.CLK(clk_i),.Q(r0_2[11:11]));
  DFFX1 desc2106(.D(n329),.CLK(clk_i),.Q(r0_2[12:12]));
  DFFX1 desc2107(.D(n328),.CLK(clk_i),.Q(r0_2[13:13]));
  DFFX1 desc2108(.D(n327),.CLK(clk_i),.Q(r0_2[14:14]));
  DFFX1 desc2109(.D(n326),.CLK(clk_i),.Q(r0_2[15:15]));
  DFFX1 desc2110(.D(n325),.CLK(clk_i),.Q(r0_2[16:16]));
  DFFX1 desc2111(.D(n324),.CLK(clk_i),.Q(r0_2[17:17]));
  DFFX1 desc2112(.D(n323),.CLK(clk_i),.Q(r0_2[18:18]));
  DFFX1 desc2113(.D(n322),.CLK(clk_i),.Q(r0_2[19:19]));
  DFFX1 desc2114(.D(n321),.CLK(clk_i),.Q(r0_2[20:20]));
  DFFX1 desc2115(.D(n320),.CLK(clk_i),.Q(r0_2[21:21]));
  DFFX1 desc2116(.D(n319),.CLK(clk_i),.Q(r0_2[22:22]));
  DFFX1 desc2117(.D(n318),.CLK(clk_i),.Q(r0_2[23:23]));
  DFFX1 desc2118(.D(n317),.CLK(clk_i),.Q(r0_2[24:24]));
  DFFX1 desc2119(.D(n316),.CLK(clk_i),.Q(r0_2[25:25]));
  DFFX1 desc2120(.D(n315),.CLK(clk_i),.Q(r0_2[26:26]));
  DFFX1 desc2121(.D(n314),.CLK(clk_i),.Q(r0_2[27:27]));
  DFFX1 desc2122(.D(n313),.CLK(clk_i),.Q(r0_2[28:28]));
  DFFX1 desc2123(.D(n312),.CLK(clk_i),.Q(r0_2[29:29]));
  DFFX1 desc2124(.D(n311),.CLK(clk_i),.Q(r0_2[30:30]));
  DFFX1 desc2125(.D(n310),.CLK(clk_i),.Q(r0_2[31:31]));
  DFFX1 desc2126(.D(n309),.CLK(clk_i),.Q(r0_2[32:32]));
  DFFX1 desc2127(.D(n308),.CLK(clk_i),.Q(r0_2[33:33]));
  DFFX1 desc2128(.D(n307),.CLK(clk_i),.Q(r0_2[34:34]));
  DFFX1 desc2129(.D(n306),.CLK(clk_i),.Q(r0_2[35:35]));
  DFFX1 desc2130(.D(n305),.CLK(clk_i),.Q(r0_2[36:36]));
  DFFX1 desc2131(.D(n304),.CLK(clk_i),.Q(r0_2[37:37]));
  DFFX1 desc2132(.D(n303),.CLK(clk_i),.Q(r0_2[38:38]));
  DFFX1 desc2133(.D(n302),.CLK(clk_i),.Q(r0_2[39:39]));
  DFFX1 desc2134(.D(n301),.CLK(clk_i),.Q(r0_2[40:40]));
  DFFX1 desc2135(.D(n300),.CLK(clk_i),.Q(r0_2[41:41]));
  DFFX1 desc2136(.D(n299),.CLK(clk_i),.Q(r0_2[42:42]));
  DFFX1 desc2137(.D(n298),.CLK(clk_i),.Q(r0_2[43:43]));
  DFFX1 desc2138(.D(n297),.CLK(clk_i),.Q(r0_2[44:44]));
  DFFX1 desc2139(.D(n296),.CLK(clk_i),.Q(r0_2[45:45]));
  DFFX1 desc2140(.D(n295),.CLK(clk_i),.Q(r0_2[46:46]));
  DFFX1 desc2141(.D(n294),.CLK(clk_i),.Q(r0_2[47:47]));
  DFFX1 desc2142(.D(n293),.CLK(clk_i),.Q(r0_2[48:48]));
  DFFX1 desc2143(.D(n292),.CLK(clk_i),.Q(r0_2[49:49]));
  DFFX1 desc2144(.D(n291),.CLK(clk_i),.Q(r0_2[50:50]));
  DFFX1 desc2145(.D(n367),.CLK(clk_i),.Q(r1[25:25]));
  DFFX1 desc2146(.D(n368),.CLK(clk_i),.Q(r1[24:24]));
  DFFX1 desc2147(.D(n369),.CLK(clk_i),.Q(r1[23:23]));
  DFFX1 desc2148(.D(n370),.CLK(clk_i),.Q(r1[22:22]));
  DFFX1 desc2149(.D(n371),.CLK(clk_i),.Q(r1[21:21]));
  DFFX1 desc2150(.D(n372),.CLK(clk_i),.Q(r1[20:20]));
  DFFX1 desc2151(.D(n373),.CLK(clk_i),.Q(r1[19:19]));
  DFFX1 desc2152(.D(n374),.CLK(clk_i),.Q(r1[18:18]));
  DFFX1 desc2153(.D(n375),.CLK(clk_i),.Q(r1[17:17]));
  DFFX1 desc2154(.D(n376),.CLK(clk_i),.Q(r1[16:16]));
  DFFX1 desc2155(.D(n377),.CLK(clk_i),.Q(r1[15:15]));
  DFFX1 desc2156(.D(n378),.CLK(clk_i),.Q(r1[14:14]));
  DFFX1 desc2157(.D(n379),.CLK(clk_i),.Q(r1[13:13]));
  DFFX1 desc2158(.D(n380),.CLK(clk_i),.Q(r1[12:12]));
  DFFX1 desc2159(.D(n381),.CLK(clk_i),.Q(r1[11:11]));
  DFFX1 desc2160(.D(n382),.CLK(clk_i),.Q(r1[10:10]));
  DFFX1 desc2161(.D(n383),.CLK(clk_i),.Q(r1[9:9]));
  DFFX1 desc2162(.D(n384),.CLK(clk_i),.Q(r1[8:8]));
  DFFX1 desc2163(.D(n385),.CLK(clk_i),.Q(r1[7:7]));
  DFFX1 desc2164(.D(n386),.CLK(clk_i),.Q(r1[6:6]));
  DFFX1 desc2165(.D(n387),.CLK(clk_i),.Q(r1[5:5]));
  DFFX1 desc2166(.D(n388),.CLK(clk_i),.Q(r1[4:4]));
  DFFX1 desc2167(.D(n389),.CLK(clk_i),.Q(r1[3:3]));
  DFFX1 desc2168(.D(n390),.CLK(clk_i),.Q(r1[2:2]));
  DFFX1 desc2169(.D(n391),.CLK(clk_i),.Q(r1[1:1]));
  DFFX1 desc2170(.D(n392),.CLK(clk_i),.Q(r1[0:0]));
  DFFX1 desc2171(.D(n289),.CLK(clk_i),.Q(r1_2[51:51]));
  DFFX1 desc2172(.D(n288),.CLK(clk_i),.Q(r1_2[50:50]));
  DFFX1 desc2173(.D(n287),.CLK(clk_i),.Q(r1_2[49:49]));
  DFFX1 desc2174(.D(n286),.CLK(clk_i),.Q(r1_2[48:48]));
  DFFX1 desc2175(.D(n285),.CLK(clk_i),.Q(r1_2[47:47]));
  DFFX1 desc2176(.D(n284),.CLK(clk_i),.Q(r1_2[46:46]));
  DFFX1 desc2177(.D(n283),.CLK(clk_i),.Q(r1_2[45:45]));
  DFFX1 desc2178(.D(n282),.CLK(clk_i),.Q(r1_2[44:44]));
  DFFX1 desc2179(.D(n281),.CLK(clk_i),.Q(r1_2[43:43]));
  DFFX1 desc2180(.D(n280),.CLK(clk_i),.Q(r1_2[42:42]));
  DFFX1 desc2181(.D(n279),.CLK(clk_i),.Q(r1_2[41:41]));
  DFFX1 desc2182(.D(n278),.CLK(clk_i),.Q(r1_2[40:40]));
  DFFX1 desc2183(.D(n277),.CLK(clk_i),.Q(r1_2[39:39]));
  DFFX1 desc2184(.D(n276),.CLK(clk_i),.Q(r1_2[38:38]));
  DFFX1 desc2185(.D(n275),.CLK(clk_i),.Q(r1_2[37:37]));
  DFFX1 desc2186(.D(n274),.CLK(clk_i),.Q(r1_2[36:36]));
  DFFX1 desc2187(.D(n273),.CLK(clk_i),.Q(r1_2[35:35]));
  DFFX1 desc2188(.D(n272),.CLK(clk_i),.Q(r1_2[34:34]));
  DFFX1 desc2189(.D(n271),.CLK(clk_i),.Q(r1_2[33:33]));
  DFFX1 desc2190(.D(n270),.CLK(clk_i),.Q(r1_2[32:32]));
  DFFX1 desc2191(.D(n269),.CLK(clk_i),.Q(r1_2[31:31]));
  DFFX1 desc2192(.D(n268),.CLK(clk_i),.Q(r1_2[30:30]));
  DFFX1 desc2193(.D(n267),.CLK(clk_i),.Q(r1_2[29:29]));
  DFFX1 desc2194(.D(n266),.CLK(clk_i),.Q(r1_2[28:28]));
  DFFX1 desc2195(.D(n265),.CLK(clk_i),.Q(r1_2[27:27]));
  DFFX1 desc2196(.D(n264),.CLK(clk_i),.Q(r1_2[26:26]));
  DFFX1 desc2197(.D(n263),.CLK(clk_i),.Q(r1_2[25:25]));
  DFFX1 desc2198(.D(n262),.CLK(clk_i),.Q(r1_2[24:24]));
  DFFX1 desc2199(.D(n261),.CLK(clk_i),.Q(r1_2[23:23]));
  DFFX1 desc2200(.D(n260),.CLK(clk_i),.Q(r1_2[22:22]));
  DFFX1 desc2201(.D(n259),.CLK(clk_i),.Q(r1_2[21:21]));
  DFFX1 desc2202(.D(n258),.CLK(clk_i),.Q(r1_2[20:20]));
  DFFX1 desc2203(.D(n257),.CLK(clk_i),.Q(r1_2[19:19]));
  DFFX1 desc2204(.D(n256),.CLK(clk_i),.Q(r1_2[18:18]));
  DFFX1 desc2205(.D(n255),.CLK(clk_i),.Q(r1_2[17:17]));
  DFFX1 desc2206(.D(n254),.CLK(clk_i),.Q(r1_2[16:16]));
  DFFX1 desc2207(.D(n253),.CLK(clk_i),.Q(r1_2[15:15]));
  DFFX1 desc2208(.D(n252),.CLK(clk_i),.Q(r1_2[14:14]));
  DFFX1 desc2209(.D(n251),.CLK(clk_i),.Q(r1_2[13:13]));
  DFFX1 desc2210(.D(n250),.CLK(clk_i),.Q(r1_2[12:12]));
  DFFX1 desc2211(.D(n249),.CLK(clk_i),.Q(r1_2[11:11]));
  DFFX1 desc2212(.D(n248),.CLK(clk_i),.Q(r1_2[10:10]));
  DFFX1 desc2213(.D(n247),.CLK(clk_i),.Q(r1_2[9:9]));
  DFFX1 desc2214(.D(n246),.CLK(clk_i),.Q(r1_2[8:8]));
  DFFX1 desc2215(.D(n245),.CLK(clk_i),.Q(r1_2[7:7]));
  DFFX1 desc2216(.D(n244),.CLK(clk_i),.Q(r1_2[6:6]));
  DFFX1 desc2217(.D(n243),.CLK(clk_i),.Q(r1_2[5:5]));
  DFFX1 desc2218(.D(n242),.CLK(clk_i),.Q(r1_2[4:4]));
  DFFX1 desc2219(.D(n241),.CLK(clk_i),.Q(r1_2[3:3]));
  DFFX1 desc2220(.D(n240),.CLK(clk_i),.Q(r1_2[2:2]));
  DFFX1 desc2221(.D(n239),.CLK(clk_i),.Q(r1_2[1:1]));
  DFFX1 desc2222(.D(n238),.CLK(clk_i),.Q(r1_2[0:0]));
  DFFX1 desc2223(.D(n237),.CLK(clk_i),.Q(s_sqr_o[25:25]));
  DFFX1 desc2224(.D(s_sqr_o[25:25]),.CLK(clk_i),.Q(sqr_o[25:25]));
  DFFX1 desc2225(.D(n236),.CLK(clk_i),.Q(s_sqr_o[24:24]));
  DFFX1 desc2226(.D(s_sqr_o[24:24]),.CLK(clk_i),.Q(sqr_o[24:24]));
  DFFX1 desc2227(.D(n235),.CLK(clk_i),.Q(s_sqr_o[23:23]));
  DFFX1 desc2228(.D(s_sqr_o[23:23]),.CLK(clk_i),.Q(sqr_o[23:23]));
  DFFX1 desc2229(.D(n234),.CLK(clk_i),.Q(s_sqr_o[22:22]));
  DFFX1 desc2230(.D(s_sqr_o[22:22]),.CLK(clk_i),.Q(sqr_o[22:22]));
  DFFX1 desc2231(.D(n233),.CLK(clk_i),.Q(s_sqr_o[21:21]));
  DFFX1 desc2232(.D(s_sqr_o[21:21]),.CLK(clk_i),.Q(sqr_o[21:21]));
  DFFX1 desc2233(.D(n232),.CLK(clk_i),.Q(s_sqr_o[20:20]));
  DFFX1 desc2234(.D(s_sqr_o[20:20]),.CLK(clk_i),.Q(sqr_o[20:20]));
  DFFX1 desc2235(.D(n231),.CLK(clk_i),.Q(s_sqr_o[19:19]));
  DFFX1 desc2236(.D(s_sqr_o[19:19]),.CLK(clk_i),.Q(sqr_o[19:19]));
  DFFX1 desc2237(.D(n230),.CLK(clk_i),.Q(s_sqr_o[18:18]));
  DFFX1 desc2238(.D(s_sqr_o[18:18]),.CLK(clk_i),.Q(sqr_o[18:18]));
  DFFX1 desc2239(.D(n229),.CLK(clk_i),.Q(s_sqr_o[17:17]));
  DFFX1 desc2240(.D(s_sqr_o[17:17]),.CLK(clk_i),.Q(sqr_o[17:17]));
  DFFX1 desc2241(.D(n228),.CLK(clk_i),.Q(s_sqr_o[16:16]));
  DFFX1 desc2242(.D(s_sqr_o[16:16]),.CLK(clk_i),.Q(sqr_o[16:16]));
  DFFX1 desc2243(.D(n227),.CLK(clk_i),.Q(s_sqr_o[15:15]));
  DFFX1 desc2244(.D(s_sqr_o[15:15]),.CLK(clk_i),.Q(sqr_o[15:15]));
  DFFX1 desc2245(.D(n226),.CLK(clk_i),.Q(s_sqr_o[14:14]));
  DFFX1 desc2246(.D(s_sqr_o[14:14]),.CLK(clk_i),.Q(sqr_o[14:14]));
  DFFX1 desc2247(.D(n225),.CLK(clk_i),.Q(s_sqr_o[13:13]));
  DFFX1 desc2248(.D(s_sqr_o[13:13]),.CLK(clk_i),.Q(sqr_o[13:13]));
  DFFX1 desc2249(.D(n224),.CLK(clk_i),.Q(s_sqr_o[12:12]));
  DFFX1 desc2250(.D(s_sqr_o[12:12]),.CLK(clk_i),.Q(sqr_o[12:12]));
  DFFX1 desc2251(.D(n223),.CLK(clk_i),.Q(s_sqr_o[11:11]));
  DFFX1 desc2252(.D(s_sqr_o[11:11]),.CLK(clk_i),.Q(sqr_o[11:11]));
  DFFX1 desc2253(.D(n222),.CLK(clk_i),.Q(s_sqr_o[10:10]));
  DFFX1 desc2254(.D(s_sqr_o[10:10]),.CLK(clk_i),.Q(sqr_o[10:10]));
  DFFX1 desc2255(.D(n221),.CLK(clk_i),.Q(s_sqr_o[9:9]));
  DFFX1 desc2256(.D(s_sqr_o[9:9]),.CLK(clk_i),.Q(sqr_o[9:9]));
  DFFX1 desc2257(.D(n220),.CLK(clk_i),.Q(s_sqr_o[8:8]));
  DFFX1 desc2258(.D(s_sqr_o[8:8]),.CLK(clk_i),.Q(sqr_o[8:8]));
  DFFX1 desc2259(.D(n219),.CLK(clk_i),.Q(s_sqr_o[7:7]));
  DFFX1 desc2260(.D(s_sqr_o[7:7]),.CLK(clk_i),.Q(sqr_o[7:7]));
  DFFX1 desc2261(.D(n218),.CLK(clk_i),.Q(s_sqr_o[6:6]));
  DFFX1 desc2262(.D(s_sqr_o[6:6]),.CLK(clk_i),.Q(sqr_o[6:6]));
  DFFX1 desc2263(.D(n217),.CLK(clk_i),.Q(s_sqr_o[5:5]));
  DFFX1 desc2264(.D(s_sqr_o[5:5]),.CLK(clk_i),.Q(sqr_o[5:5]));
  DFFX1 desc2265(.D(n216),.CLK(clk_i),.Q(s_sqr_o[4:4]));
  DFFX1 desc2266(.D(s_sqr_o[4:4]),.CLK(clk_i),.Q(sqr_o[4:4]));
  DFFX1 desc2267(.D(n215),.CLK(clk_i),.Q(s_sqr_o[3:3]));
  DFFX1 desc2268(.D(s_sqr_o[3:3]),.CLK(clk_i),.Q(sqr_o[3:3]));
  DFFX1 desc2269(.D(n214),.CLK(clk_i),.Q(s_sqr_o[2:2]));
  DFFX1 desc2270(.D(s_sqr_o[2:2]),.CLK(clk_i),.Q(sqr_o[2:2]));
  DFFX1 desc2271(.D(n213),.CLK(clk_i),.Q(s_sqr_o[1:1]));
  DFFX1 desc2272(.D(s_sqr_o[1:1]),.CLK(clk_i),.Q(sqr_o[1:1]));
  DFFX1 desc2273(.D(n212),.CLK(clk_i),.Q(s_sqr_o[0:0]));
  DFFX1 desc2274(.D(s_sqr_o[0:0]),.CLK(clk_i),.Q(sqr_o[0:0]));
  DFFX1 s_ine_o_reg(.D(n211),.CLK(clk_i),.Q(s_ine_o));
  DFFX1 ine_o_reg(.D(s_ine_o),.CLK(clk_i),.Q(ine_o));
  AO22X1 U3(.IN1(s_ine_o),.IN2(n437),.IN3(n44),.IN4(n45),.Q(n211));
  NAND4X0 U6(.IN1(n49),.IN2(n50),.IN3(n51),.IN4(n52),.QN(n48));
  NOR4X0 U7(.IN1(n53),.IN2(n54),.IN3(n55),.IN4(n56),.QN(n52));
  XOR2X1 U8(.IN1(s_rad_i[34:34]),.IN2(N448),.Q(n56));
  XOR2X1 U9(.IN1(s_rad_i[40:40]),.IN2(N454),.Q(n55));
  XOR2X1 U10(.IN1(s_rad_i[41:41]),.IN2(N455),.Q(n54));
  NAND4X0 U20(.IN1(n57),.IN2(n58),.IN3(n59),.IN4(n60),.QN(n53));
  XOR2X1 U21(.IN1(n189),.IN2(N440),.Q(n60));
  XOR2X1 U22(.IN1(n190),.IN2(N441),.Q(n59));
  XOR2X1 U23(.IN1(n166),.IN2(N443),.Q(n58));
  XOR2X1 U24(.IN1(n167),.IN2(N442),.Q(n57));
  NOR4X0 U25(.IN1(n61),.IN2(n62),.IN3(n63),.IN4(n64),.QN(n51));
  XOR2X1 U26(.IN1(s_rad_i[3:3]),.IN2(N417),.Q(n64));
  XOR2X1 U27(.IN1(s_rad_i[13:13]),.IN2(N427),.Q(n63));
  XOR2X1 U28(.IN1(s_rad_i[14:14]),.IN2(N428),.Q(n62));
  NAND3X0 U29(.IN1(n65),.IN2(n66),.IN3(n67),.QN(n61));
  XOR2X1 U30(.IN1(n173),.IN2(N416),.Q(n67));
  XOR2X1 U31(.IN1(n174),.IN2(N415),.Q(n66));
  XOR2X1 U32(.IN1(n169),.IN2(N456),.Q(n65));
  NOR4X0 U33(.IN1(n68),.IN2(n69),.IN3(n70),.IN4(n71),.QN(n50));
  XOR2X1 U34(.IN1(s_rad_i[45:45]),.IN2(N459),.Q(n71));
  XOR2X1 U35(.IN1(s_rad_i[44:44]),.IN2(N458),.Q(n70));
  XOR2X1 U36(.IN1(s_rad_i[43:43]),.IN2(N457),.Q(n69));
  NAND4X0 U37(.IN1(n72),.IN2(n73),.IN3(n74),.IN4(n75),.QN(n68));
  XOR2X1 U38(.IN1(n176),.IN2(N429),.Q(n75));
  XOR2X1 U39(.IN1(n180),.IN2(N446),.Q(n74));
  XOR2X1 U40(.IN1(n181),.IN2(N444),.Q(n73));
  XOR2X1 U41(.IN1(n182),.IN2(N445),.Q(n72));
  NOR4X0 U42(.IN1(n76),.IN2(n77),.IN3(n78),.IN4(n79),.QN(n49));
  XOR2X1 U43(.IN1(s_rad_i[18:18]),.IN2(N432),.Q(n79));
  XOR2X1 U44(.IN1(s_rad_i[23:23]),.IN2(N437),.Q(n78));
  XOR2X1 U45(.IN1(s_rad_i[19:19]),.IN2(N433),.Q(n77));
  NAND3X0 U46(.IN1(n80),.IN2(n81),.IN3(n82),.QN(n76));
  XOR2X1 U47(.IN1(n187),.IN2(N420),.Q(n82));
  XOR2X1 U48(.IN1(n188),.IN2(N424),.Q(n81));
  XOR2X1 U49(.IN1(n186),.IN2(N419),.Q(n80));
  NAND4X0 U50(.IN1(n83),.IN2(n84),.IN3(n85),.IN4(n86),.QN(n47));
  NOR4X0 U51(.IN1(n87),.IN2(n88),.IN3(n89),.IN4(n90),.QN(n86));
  XOR2X1 U52(.IN1(s_rad_i[48:48]),.IN2(N462),.Q(n90));
  XOR2X1 U53(.IN1(s_rad_i[0:0]),.IN2(N414),.Q(n89));
  XOR2X1 U54(.IN1(s_rad_i[46:46]),.IN2(N460),.Q(n88));
  NAND4X0 U55(.IN1(n91),.IN2(n92),.IN3(n93),.IN4(n94),.QN(n87));
  XOR2X1 U56(.IN1(n163),.IN2(N453),.Q(n94));
  XOR2X1 U57(.IN1(n164),.IN2(N449),.Q(n93));
  XOR2X1 U58(.IN1(n165),.IN2(N447),.Q(n92));
  XOR2X1 U59(.IN1(n168),.IN2(N461),.Q(n91));
  NOR4X0 U60(.IN1(n95),.IN2(n96),.IN3(n97),.IN4(n98),.QN(n85));
  XOR2X1 U61(.IN1(s_rad_i[16:16]),.IN2(N430),.Q(n98));
  XOR2X1 U62(.IN1(s_rad_i[22:22]),.IN2(N436),.Q(n97));
  XOR2X1 U63(.IN1(s_rad_i[21:21]),.IN2(N435),.Q(n96));
  NAND3X0 U64(.IN1(n99),.IN2(n100),.IN3(n101),.QN(n95));
  XOR2X1 U65(.IN1(n171),.IN2(N422),.Q(n101));
  XOR2X1 U66(.IN1(n172),.IN2(N423),.Q(n100));
  XOR2X1 U67(.IN1(n170),.IN2(N421),.Q(n99));
  NOR4X0 U68(.IN1(n102),.IN2(n103),.IN3(n104),.IN4(n105),.QN(n84));
  XOR2X1 U69(.IN1(s_rad_i[49:49]),.IN2(N463),.Q(n105));
  XOR2X1 U70(.IN1(s_rad_i[50:50]),.IN2(N464),.Q(n104));
  XOR2X1 U71(.IN1(s_rad_i[51:51]),.IN2(N465),.Q(n103));
  NAND4X0 U72(.IN1(n106),.IN2(n107),.IN3(n108),.IN4(n109),.QN(n102));
  XOR2X1 U73(.IN1(n175),.IN2(N434),.Q(n109));
  XOR2X1 U74(.IN1(n177),.IN2(N451),.Q(n108));
  XOR2X1 U75(.IN1(n178),.IN2(N450),.Q(n107));
  XOR2X1 U76(.IN1(n179),.IN2(N452),.Q(n106));
  NOR4X0 U77(.IN1(n110),.IN2(n111),.IN3(n112),.IN4(n113),.QN(n83));
  XOR2X1 U78(.IN1(s_rad_i[11:11]),.IN2(N425),.Q(n113));
  XOR2X1 U79(.IN1(s_rad_i[24:24]),.IN2(N438),.Q(n112));
  XOR2X1 U80(.IN1(s_rad_i[25:25]),.IN2(N439),.Q(n111));
  NAND3X0 U81(.IN1(n114),.IN2(n115),.IN3(n116),.QN(n110));
  XOR2X1 U82(.IN1(n184),.IN2(N431),.Q(n116));
  XOR2X1 U83(.IN1(n185),.IN2(N426),.Q(n115));
  XOR2X1 U84(.IN1(n183),.IN2(N418),.Q(n114));
  AO22X1 U86(.IN1(s_sqr_o[0:0]),.IN2(n15),.IN3(N309),.IN4(n419),.Q(n212));
  AO22X1 U87(.IN1(s_sqr_o[1:1]),.IN2(n15),.IN3(N310),.IN4(n419),.Q(n213));
  AO22X1 U88(.IN1(s_sqr_o[2:2]),.IN2(n15),.IN3(N311),.IN4(n419),.Q(n214));
  AO22X1 U89(.IN1(s_sqr_o[3:3]),.IN2(n15),.IN3(N312),.IN4(n419),.Q(n215));
  AO22X1 U90(.IN1(s_sqr_o[4:4]),.IN2(n15),.IN3(N313),.IN4(n419),.Q(n216));
  AO22X1 U91(.IN1(s_sqr_o[5:5]),.IN2(n15),.IN3(N314),.IN4(n419),.Q(n217));
  AO22X1 U92(.IN1(s_sqr_o[6:6]),.IN2(n15),.IN3(N315),.IN4(n419),.Q(n218));
  AO22X1 U93(.IN1(s_sqr_o[7:7]),.IN2(n15),.IN3(N316),.IN4(n419),.Q(n219));
  AO22X1 U94(.IN1(s_sqr_o[8:8]),.IN2(n15),.IN3(N317),.IN4(n419),.Q(n220));
  AO22X1 U95(.IN1(s_sqr_o[9:9]),.IN2(n15),.IN3(N318),.IN4(n419),.Q(n221));
  AO22X1 U96(.IN1(s_sqr_o[10:10]),.IN2(n15),.IN3(N319),.IN4(n419),.Q(n222));
  AO22X1 U97(.IN1(s_sqr_o[11:11]),.IN2(n15),.IN3(N320),.IN4(n419),.Q(n223));
  AO22X1 U98(.IN1(s_sqr_o[12:12]),.IN2(n15),.IN3(N321),.IN4(n420),.Q(n224));
  AO22X1 U99(.IN1(s_sqr_o[13:13]),.IN2(n15),.IN3(N322),.IN4(n420),.Q(n225));
  AO22X1 U100(.IN1(s_sqr_o[14:14]),.IN2(n15),.IN3(N323),.IN4(n420),.Q(n226));
  AO22X1 U101(.IN1(s_sqr_o[15:15]),.IN2(n15),.IN3(N324),.IN4(n420),.Q(n227));
  AO22X1 U102(.IN1(s_sqr_o[16:16]),.IN2(n15),.IN3(N325),.IN4(n420),.Q(n228));
  AO22X1 U103(.IN1(s_sqr_o[17:17]),.IN2(n15),.IN3(N326),.IN4(n420),.Q(n229));
  AO22X1 U104(.IN1(s_sqr_o[18:18]),.IN2(n15),.IN3(N327),.IN4(n420),.Q(n230));
  AO22X1 U105(.IN1(s_sqr_o[19:19]),.IN2(n15),.IN3(N328),.IN4(n420),.Q(n231));
  AO22X1 U106(.IN1(s_sqr_o[20:20]),.IN2(n15),.IN3(N329),.IN4(n420),.Q(n232));
  AO22X1 U107(.IN1(s_sqr_o[21:21]),.IN2(n15),.IN3(N330),.IN4(n420),.Q(n233));
  AO22X1 U108(.IN1(s_sqr_o[22:22]),.IN2(n15),.IN3(N331),.IN4(n420),.Q(n234));
  AO22X1 U109(.IN1(s_sqr_o[23:23]),.IN2(n15),.IN3(N332),.IN4(n420),.Q(n235));
  AO22X1 U110(.IN1(s_sqr_o[24:24]),.IN2(n15),.IN3(N333),.IN4(n421),.Q(n236));
  AO22X1 U111(.IN1(s_sqr_o[25:25]),.IN2(n15),.IN3(N334),.IN4(n421),.Q(n237));
  AO222X1 U114(.IN1(s_sum1b[0:0]),.IN2(n412),.IN3(s_sum2b[0:0]),.IN4(n405),.IN5(r1_2[0:0]),.IN6(n22),.Q(n238));
  AO222X1 U115(.IN1(s_sum1b[1:1]),.IN2(n412),.IN3(s_sum2b[1:1]),.IN4(n405),.IN5(r1_2[1:1]),.IN6(n404),.Q(n239));
  AO222X1 U116(.IN1(s_sum1b[2:2]),.IN2(n412),.IN3(s_sum2b[2:2]),.IN4(n405),.IN5(r1_2[2:2]),.IN6(n404),.Q(n240));
  AO222X1 U117(.IN1(s_sum1b[3:3]),.IN2(n412),.IN3(s_sum2b[3:3]),.IN4(n405),.IN5(r1_2[3:3]),.IN6(n404),.Q(n241));
  AO222X1 U118(.IN1(s_sum1b[4:4]),.IN2(n412),.IN3(s_sum2b[4:4]),.IN4(n405),.IN5(r1_2[4:4]),.IN6(n404),.Q(n242));
  AO222X1 U119(.IN1(s_sum1b[5:5]),.IN2(n412),.IN3(s_sum2b[5:5]),.IN4(n405),.IN5(r1_2[5:5]),.IN6(n404),.Q(n243));
  AO222X1 U120(.IN1(s_sum1b[6:6]),.IN2(n412),.IN3(s_sum2b[6:6]),.IN4(n405),.IN5(r1_2[6:6]),.IN6(n404),.Q(n244));
  AO222X1 U121(.IN1(s_sum1b[7:7]),.IN2(n412),.IN3(s_sum2b[7:7]),.IN4(n405),.IN5(r1_2[7:7]),.IN6(n404),.Q(n245));
  AO222X1 U122(.IN1(s_sum1b[8:8]),.IN2(n412),.IN3(s_sum2b[8:8]),.IN4(n405),.IN5(r1_2[8:8]),.IN6(n404),.Q(n246));
  AO222X1 U123(.IN1(s_sum1b[9:9]),.IN2(n412),.IN3(s_sum2b[9:9]),.IN4(n405),.IN5(r1_2[9:9]),.IN6(n404),.Q(n247));
  AO222X1 U124(.IN1(s_sum1b[10:10]),.IN2(n412),.IN3(s_sum2b[10:10]),.IN4(n405),.IN5(r1_2[10:10]),.IN6(n404),.Q(n248));
  AO222X1 U125(.IN1(s_sum1b[11:11]),.IN2(n412),.IN3(s_sum2b[11:11]),.IN4(n405),.IN5(r1_2[11:11]),.IN6(n404),.Q(n249));
  AO222X1 U126(.IN1(s_sum1b[12:12]),.IN2(n413),.IN3(s_sum2b[12:12]),.IN4(n406),.IN5(r1_2[12:12]),.IN6(n404),.Q(n250));
  AO222X1 U127(.IN1(s_sum1b[13:13]),.IN2(n413),.IN3(s_sum2b[13:13]),.IN4(n406),.IN5(r1_2[13:13]),.IN6(n403),.Q(n251));
  AO222X1 U128(.IN1(s_sum1b[14:14]),.IN2(n413),.IN3(s_sum2b[14:14]),.IN4(n406),.IN5(r1_2[14:14]),.IN6(n403),.Q(n252));
  AO222X1 U129(.IN1(s_sum1b[15:15]),.IN2(n413),.IN3(s_sum2b[15:15]),.IN4(n406),.IN5(r1_2[15:15]),.IN6(n403),.Q(n253));
  AO222X1 U130(.IN1(s_sum1b[16:16]),.IN2(n413),.IN3(s_sum2b[16:16]),.IN4(n406),.IN5(r1_2[16:16]),.IN6(n403),.Q(n254));
  AO222X1 U131(.IN1(s_sum1b[17:17]),.IN2(n413),.IN3(s_sum2b[17:17]),.IN4(n406),.IN5(r1_2[17:17]),.IN6(n403),.Q(n255));
  AO222X1 U132(.IN1(s_sum1b[18:18]),.IN2(n413),.IN3(s_sum2b[18:18]),.IN4(n406),.IN5(r1_2[18:18]),.IN6(n403),.Q(n256));
  AO222X1 U133(.IN1(s_sum1b[19:19]),.IN2(n413),.IN3(s_sum2b[19:19]),.IN4(n406),.IN5(r1_2[19:19]),.IN6(n403),.Q(n257));
  AO222X1 U134(.IN1(s_sum1b[20:20]),.IN2(n413),.IN3(s_sum2b[20:20]),.IN4(n406),.IN5(r1_2[20:20]),.IN6(n403),.Q(n258));
  AO222X1 U135(.IN1(s_sum1b[21:21]),.IN2(n413),.IN3(s_sum2b[21:21]),.IN4(n406),.IN5(r1_2[21:21]),.IN6(n403),.Q(n259));
  AO222X1 U136(.IN1(s_sum1b[22:22]),.IN2(n413),.IN3(s_sum2b[22:22]),.IN4(n406),.IN5(r1_2[22:22]),.IN6(n403),.Q(n260));
  AO222X1 U137(.IN1(s_sum1b[23:23]),.IN2(n413),.IN3(s_sum2b[23:23]),.IN4(n406),.IN5(r1_2[23:23]),.IN6(n403),.Q(n261));
  AO222X1 U138(.IN1(s_sum1b[24:24]),.IN2(n414),.IN3(s_sum2b[24:24]),.IN4(n407),.IN5(r1_2[24:24]),.IN6(n403),.Q(n262));
  AO222X1 U139(.IN1(s_sum1b[25:25]),.IN2(n414),.IN3(s_sum2b[25:25]),.IN4(n407),.IN5(r1_2[25:25]),.IN6(n403),.Q(n263));
  AO222X1 U140(.IN1(s_sum1b[26:26]),.IN2(n414),.IN3(s_sum2b[26:26]),.IN4(n407),.IN5(r1_2[26:26]),.IN6(n403),.Q(n264));
  AO222X1 U141(.IN1(s_sum1b[27:27]),.IN2(n414),.IN3(s_sum2b[27:27]),.IN4(n407),.IN5(r1_2[27:27]),.IN6(n403),.Q(n265));
  AO222X1 U142(.IN1(s_sum1b[28:28]),.IN2(n414),.IN3(s_sum2b[28:28]),.IN4(n407),.IN5(r1_2[28:28]),.IN6(n403),.Q(n266));
  AO222X1 U143(.IN1(s_sum1b[29:29]),.IN2(n414),.IN3(s_sum2b[29:29]),.IN4(n407),.IN5(r1_2[29:29]),.IN6(n403),.Q(n267));
  AO222X1 U144(.IN1(s_sum1b[30:30]),.IN2(n414),.IN3(s_sum2b[30:30]),.IN4(n407),.IN5(r1_2[30:30]),.IN6(n403),.Q(n268));
  AO222X1 U145(.IN1(s_sum1b[31:31]),.IN2(n414),.IN3(s_sum2b[31:31]),.IN4(n407),.IN5(r1_2[31:31]),.IN6(n403),.Q(n269));
  AO222X1 U146(.IN1(s_sum1b[32:32]),.IN2(n414),.IN3(s_sum2b[32:32]),.IN4(n407),.IN5(r1_2[32:32]),.IN6(n403),.Q(n270));
  AO222X1 U147(.IN1(s_sum1b[33:33]),.IN2(n414),.IN3(s_sum2b[33:33]),.IN4(n407),.IN5(r1_2[33:33]),.IN6(n403),.Q(n271));
  AO222X1 U148(.IN1(s_sum1b[34:34]),.IN2(n414),.IN3(s_sum2b[34:34]),.IN4(n407),.IN5(r1_2[34:34]),.IN6(n403),.Q(n272));
  AO222X1 U149(.IN1(s_sum1b[35:35]),.IN2(n414),.IN3(s_sum2b[35:35]),.IN4(n407),.IN5(r1_2[35:35]),.IN6(n403),.Q(n273));
  AO222X1 U150(.IN1(s_sum1b[36:36]),.IN2(n415),.IN3(s_sum2b[36:36]),.IN4(n408),.IN5(r1_2[36:36]),.IN6(n403),.Q(n274));
  AO222X1 U151(.IN1(s_sum1b[37:37]),.IN2(n415),.IN3(s_sum2b[37:37]),.IN4(n408),.IN5(r1_2[37:37]),.IN6(n403),.Q(n275));
  AO222X1 U152(.IN1(s_sum1b[38:38]),.IN2(n415),.IN3(s_sum2b[38:38]),.IN4(n408),.IN5(r1_2[38:38]),.IN6(n403),.Q(n276));
  AO222X1 U153(.IN1(s_sum1b[39:39]),.IN2(n415),.IN3(s_sum2b[39:39]),.IN4(n408),.IN5(r1_2[39:39]),.IN6(n403),.Q(n277));
  AO222X1 U154(.IN1(s_sum1b[40:40]),.IN2(n415),.IN3(s_sum2b[40:40]),.IN4(n408),.IN5(r1_2[40:40]),.IN6(n403),.Q(n278));
  AO222X1 U155(.IN1(s_sum1b[41:41]),.IN2(n415),.IN3(s_sum2b[41:41]),.IN4(n408),.IN5(r1_2[41:41]),.IN6(n403),.Q(n279));
  AO222X1 U156(.IN1(s_sum1b[42:42]),.IN2(n415),.IN3(s_sum2b[42:42]),.IN4(n408),.IN5(r1_2[42:42]),.IN6(n403),.Q(n280));
  AO222X1 U157(.IN1(s_sum1b[43:43]),.IN2(n415),.IN3(s_sum2b[43:43]),.IN4(n408),.IN5(r1_2[43:43]),.IN6(n403),.Q(n281));
  AO222X1 U158(.IN1(s_sum1b[44:44]),.IN2(n415),.IN3(s_sum2b[44:44]),.IN4(n408),.IN5(r1_2[44:44]),.IN6(n403),.Q(n282));
  AO222X1 U159(.IN1(s_sum1b[45:45]),.IN2(n415),.IN3(s_sum2b[45:45]),.IN4(n408),.IN5(r1_2[45:45]),.IN6(n403),.Q(n283));
  AO222X1 U160(.IN1(s_sum1b[46:46]),.IN2(n415),.IN3(s_sum2b[46:46]),.IN4(n408),.IN5(r1_2[46:46]),.IN6(n403),.Q(n284));
  AO222X1 U161(.IN1(s_sum1b[47:47]),.IN2(n415),.IN3(s_sum2b[47:47]),.IN4(n408),.IN5(r1_2[47:47]),.IN6(n403),.Q(n285));
  AO222X1 U162(.IN1(s_sum1b[48:48]),.IN2(n416),.IN3(s_sum2b[48:48]),.IN4(n409),.IN5(r1_2[48:48]),.IN6(n23),.Q(n286));
  AO222X1 U163(.IN1(s_sum1b[49:49]),.IN2(n416),.IN3(s_sum2b[49:49]),.IN4(n409),.IN5(r1_2[49:49]),.IN6(n22),.Q(n287));
  AO222X1 U164(.IN1(s_sum1b[50:50]),.IN2(n416),.IN3(s_sum2b[50:50]),.IN4(n409),.IN5(r1_2[50:50]),.IN6(n23),.Q(n288));
  AO222X1 U165(.IN1(s_sum1b[51:51]),.IN2(n416),.IN3(s_sum2b[51:51]),.IN4(n409),.IN5(r1_2[51:51]),.IN6(n22),.Q(n289));
  AO222X1 U166(.IN1(n125),.IN2(s_sum1b[51:51]),.IN3(n38),.IN4(s_sum2b[51:51]),.IN5(r0_2[51:51]),.IN6(n124),.Q(n290));
  AO222X1 U167(.IN1(n127),.IN2(s_sum1b[50:50]),.IN3(n40),.IN4(s_sum2b[50:50]),.IN5(r0_2[50:50]),.IN6(n19),.Q(n291));
  AO222X1 U168(.IN1(n127),.IN2(s_sum1b[49:49]),.IN3(n40),.IN4(s_sum2b[49:49]),.IN5(r0_2[49:49]),.IN6(n20),.Q(n292));
  AO222X1 U169(.IN1(n127),.IN2(s_sum1b[48:48]),.IN3(n40),.IN4(s_sum2b[48:48]),.IN5(r0_2[48:48]),.IN6(n19),.Q(n293));
  AO222X1 U170(.IN1(n127),.IN2(s_sum1b[47:47]),.IN3(n40),.IN4(s_sum2b[47:47]),.IN5(r0_2[47:47]),.IN6(n20),.Q(n294));
  AO222X1 U171(.IN1(n126),.IN2(s_sum1b[46:46]),.IN3(n39),.IN4(s_sum2b[46:46]),.IN5(r0_2[46:46]),.IN6(n19),.Q(n295));
  AO222X1 U172(.IN1(n126),.IN2(s_sum1b[45:45]),.IN3(n39),.IN4(s_sum2b[45:45]),.IN5(r0_2[45:45]),.IN6(n20),.Q(n296));
  AO222X1 U173(.IN1(n126),.IN2(s_sum1b[44:44]),.IN3(n39),.IN4(s_sum2b[44:44]),.IN5(r0_2[44:44]),.IN6(n19),.Q(n297));
  AO222X1 U174(.IN1(n126),.IN2(s_sum1b[43:43]),.IN3(n39),.IN4(s_sum2b[43:43]),.IN5(r0_2[43:43]),.IN6(n20),.Q(n298));
  AO222X1 U175(.IN1(n126),.IN2(s_sum1b[42:42]),.IN3(n39),.IN4(s_sum2b[42:42]),.IN5(r0_2[42:42]),.IN6(n19),.Q(n299));
  AO222X1 U176(.IN1(n126),.IN2(s_sum1b[41:41]),.IN3(n39),.IN4(s_sum2b[41:41]),.IN5(r0_2[41:41]),.IN6(n20),.Q(n300));
  AO222X1 U177(.IN1(n126),.IN2(s_sum1b[40:40]),.IN3(n39),.IN4(s_sum2b[40:40]),.IN5(r0_2[40:40]),.IN6(n19),.Q(n301));
  AO222X1 U178(.IN1(n126),.IN2(s_sum1b[39:39]),.IN3(n39),.IN4(s_sum2b[39:39]),.IN5(r0_2[39:39]),.IN6(n20),.Q(n302));
  AO222X1 U179(.IN1(n126),.IN2(s_sum1b[38:38]),.IN3(n39),.IN4(s_sum2b[38:38]),.IN5(r0_2[38:38]),.IN6(n19),.Q(n303));
  AO222X1 U180(.IN1(n126),.IN2(s_sum1b[37:37]),.IN3(n39),.IN4(s_sum2b[37:37]),.IN5(r0_2[37:37]),.IN6(n20),.Q(n304));
  AO222X1 U181(.IN1(n126),.IN2(s_sum1b[36:36]),.IN3(n39),.IN4(s_sum2b[36:36]),.IN5(r0_2[36:36]),.IN6(n19),.Q(n305));
  AO222X1 U182(.IN1(n126),.IN2(s_sum1b[35:35]),.IN3(n39),.IN4(s_sum2b[35:35]),.IN5(r0_2[35:35]),.IN6(n20),.Q(n306));
  AO222X1 U183(.IN1(n125),.IN2(s_sum1b[34:34]),.IN3(n38),.IN4(s_sum2b[34:34]),.IN5(r0_2[34:34]),.IN6(n19),.Q(n307));
  AO222X1 U184(.IN1(n125),.IN2(s_sum1b[33:33]),.IN3(n38),.IN4(s_sum2b[33:33]),.IN5(r0_2[33:33]),.IN6(n20),.Q(n308));
  AO222X1 U185(.IN1(n125),.IN2(s_sum1b[32:32]),.IN3(n38),.IN4(s_sum2b[32:32]),.IN5(r0_2[32:32]),.IN6(n19),.Q(n309));
  AO222X1 U186(.IN1(n125),.IN2(s_sum1b[31:31]),.IN3(n38),.IN4(s_sum2b[31:31]),.IN5(r0_2[31:31]),.IN6(n20),.Q(n310));
  AO222X1 U187(.IN1(n125),.IN2(s_sum1b[30:30]),.IN3(n38),.IN4(s_sum2b[30:30]),.IN5(r0_2[30:30]),.IN6(n19),.Q(n311));
  AO222X1 U188(.IN1(n125),.IN2(s_sum1b[29:29]),.IN3(n38),.IN4(s_sum2b[29:29]),.IN5(r0_2[29:29]),.IN6(n20),.Q(n312));
  AO222X1 U189(.IN1(n125),.IN2(s_sum1b[28:28]),.IN3(n38),.IN4(s_sum2b[28:28]),.IN5(r0_2[28:28]),.IN6(n19),.Q(n313));
  AO222X1 U190(.IN1(n125),.IN2(s_sum1b[27:27]),.IN3(n38),.IN4(s_sum2b[27:27]),.IN5(r0_2[27:27]),.IN6(n20),.Q(n314));
  AO222X1 U191(.IN1(n125),.IN2(s_sum1b[26:26]),.IN3(n38),.IN4(s_sum2b[26:26]),.IN5(r0_2[26:26]),.IN6(n19),.Q(n315));
  AO222X1 U192(.IN1(n125),.IN2(s_sum1b[25:25]),.IN3(n38),.IN4(s_sum2b[25:25]),.IN5(r0_2[25:25]),.IN6(n20),.Q(n316));
  AO222X1 U193(.IN1(n125),.IN2(s_sum1b[24:24]),.IN3(n38),.IN4(s_sum2b[24:24]),.IN5(r0_2[24:24]),.IN6(n19),.Q(n317));
  AO222X1 U194(.IN1(n117),.IN2(s_sum1b[23:23]),.IN3(n37),.IN4(s_sum2b[23:23]),.IN5(r0_2[23:23]),.IN6(n20),.Q(n318));
  AO222X1 U195(.IN1(n117),.IN2(s_sum1b[22:22]),.IN3(n37),.IN4(s_sum2b[22:22]),.IN5(r0_2[22:22]),.IN6(n124),.Q(n319));
  AO222X1 U196(.IN1(n117),.IN2(s_sum1b[21:21]),.IN3(n37),.IN4(s_sum2b[21:21]),.IN5(r0_2[21:21]),.IN6(n19),.Q(n320));
  AO222X1 U197(.IN1(n117),.IN2(s_sum1b[20:20]),.IN3(n37),.IN4(s_sum2b[20:20]),.IN5(r0_2[20:20]),.IN6(n124),.Q(n321));
  AO222X1 U198(.IN1(n117),.IN2(s_sum1b[19:19]),.IN3(n37),.IN4(s_sum2b[19:19]),.IN5(r0_2[19:19]),.IN6(n18),.Q(n322));
  AO222X1 U199(.IN1(n117),.IN2(s_sum1b[18:18]),.IN3(n37),.IN4(s_sum2b[18:18]),.IN5(r0_2[18:18]),.IN6(n124),.Q(n323));
  AO222X1 U200(.IN1(n117),.IN2(s_sum1b[17:17]),.IN3(n37),.IN4(s_sum2b[17:17]),.IN5(r0_2[17:17]),.IN6(n20),.Q(n324));
  AO222X1 U201(.IN1(n117),.IN2(s_sum1b[16:16]),.IN3(n37),.IN4(s_sum2b[16:16]),.IN5(r0_2[16:16]),.IN6(n124),.Q(n325));
  AO222X1 U202(.IN1(n117),.IN2(s_sum1b[15:15]),.IN3(n37),.IN4(s_sum2b[15:15]),.IN5(r0_2[15:15]),.IN6(n19),.Q(n326));
  AO222X1 U203(.IN1(n117),.IN2(s_sum1b[14:14]),.IN3(n37),.IN4(s_sum2b[14:14]),.IN5(r0_2[14:14]),.IN6(n124),.Q(n327));
  AO222X1 U204(.IN1(n117),.IN2(s_sum1b[13:13]),.IN3(n37),.IN4(s_sum2b[13:13]),.IN5(r0_2[13:13]),.IN6(n18),.Q(n328));
  AO222X1 U205(.IN1(n117),.IN2(s_sum1b[12:12]),.IN3(n37),.IN4(s_sum2b[12:12]),.IN5(r0_2[12:12]),.IN6(n18),.Q(n329));
  AO222X1 U206(.IN1(n43),.IN2(s_sum1b[11:11]),.IN3(n36),.IN4(s_sum2b[11:11]),.IN5(r0_2[11:11]),.IN6(n20),.Q(n330));
  AO222X1 U207(.IN1(n43),.IN2(s_sum1b[10:10]),.IN3(n36),.IN4(s_sum2b[10:10]),.IN5(r0_2[10:10]),.IN6(n18),.Q(n331));
  AO222X1 U208(.IN1(n43),.IN2(s_sum1b[9:9]),.IN3(n36),.IN4(s_sum2b[9:9]),.IN5(r0_2[9:9]),.IN6(n19),.Q(n332));
  AO222X1 U209(.IN1(n43),.IN2(s_sum1b[8:8]),.IN3(n36),.IN4(s_sum2b[8:8]),.IN5(r0_2[8:8]),.IN6(n18),.Q(n333));
  AO222X1 U210(.IN1(n43),.IN2(s_sum1b[7:7]),.IN3(n36),.IN4(s_sum2b[7:7]),.IN5(r0_2[7:7]),.IN6(n18),.Q(n334));
  AO222X1 U211(.IN1(n43),.IN2(s_sum1b[6:6]),.IN3(n36),.IN4(s_sum2b[6:6]),.IN5(r0_2[6:6]),.IN6(n18),.Q(n335));
  AO222X1 U212(.IN1(n43),.IN2(s_sum1b[5:5]),.IN3(n36),.IN4(s_sum2b[5:5]),.IN5(r0_2[5:5]),.IN6(n20),.Q(n336));
  AO222X1 U213(.IN1(n43),.IN2(s_sum1b[4:4]),.IN3(n36),.IN4(s_sum2b[4:4]),.IN5(r0_2[4:4]),.IN6(n18),.Q(n337));
  AO222X1 U214(.IN1(n43),.IN2(s_sum1b[3:3]),.IN3(n36),.IN4(s_sum2b[3:3]),.IN5(r0_2[3:3]),.IN6(n19),.Q(n338));
  AO222X1 U215(.IN1(n43),.IN2(s_sum1b[2:2]),.IN3(n36),.IN4(s_sum2b[2:2]),.IN5(r0_2[2:2]),.IN6(n18),.Q(n339));
  AO222X1 U216(.IN1(n43),.IN2(s_sum1b[1:1]),.IN3(n36),.IN4(s_sum2b[1:1]),.IN5(r0_2[1:1]),.IN6(n18),.Q(n340));
  AO222X1 U217(.IN1(s_sum1a[25:25]),.IN2(n127),.IN3(s_sum2a[25:25]),.IN4(n40),.IN5(r0[25:25]),.IN6(n124),.Q(n341));
  AO222X1 U218(.IN1(s_sum1a[24:24]),.IN2(n127),.IN3(s_sum2a[24:24]),.IN4(n40),.IN5(r0[24:24]),.IN6(n124),.Q(n342));
  AO222X1 U219(.IN1(s_sum1a[23:23]),.IN2(n127),.IN3(s_sum2a[23:23]),.IN4(n40),.IN5(r0[23:23]),.IN6(n124),.Q(n343));
  AO222X1 U220(.IN1(s_sum1a[22:22]),.IN2(n401),.IN3(s_sum2a[22:22]),.IN4(n42),.IN5(r0[22:22]),.IN6(n124),.Q(n344));
  AO222X1 U221(.IN1(s_sum1a[21:21]),.IN2(n127),.IN3(s_sum2a[21:21]),.IN4(n40),.IN5(r0[21:21]),.IN6(n124),.Q(n345));
  AO222X1 U222(.IN1(s_sum1a[20:20]),.IN2(n127),.IN3(s_sum2a[20:20]),.IN4(n40),.IN5(r0[20:20]),.IN6(n124),.Q(n346));
  AO222X1 U223(.IN1(s_sum1a[19:19]),.IN2(n127),.IN3(s_sum2a[19:19]),.IN4(n40),.IN5(r0[19:19]),.IN6(n124),.Q(n347));
  AO222X1 U224(.IN1(s_sum1a[18:18]),.IN2(n127),.IN3(s_sum2a[18:18]),.IN4(n40),.IN5(r0[18:18]),.IN6(n124),.Q(n348));
  AO222X1 U225(.IN1(s_sum1a[17:17]),.IN2(n127),.IN3(s_sum2a[17:17]),.IN4(n40),.IN5(r0[17:17]),.IN6(n124),.Q(n349));
  AO222X1 U226(.IN1(s_sum1a[16:16]),.IN2(n127),.IN3(s_sum2a[16:16]),.IN4(n40),.IN5(r0[16:16]),.IN6(n18),.Q(n350));
  AO222X1 U227(.IN1(s_sum1a[15:15]),.IN2(n130),.IN3(s_sum2a[15:15]),.IN4(n41),.IN5(r0[15:15]),.IN6(n19),.Q(n351));
  AO222X1 U228(.IN1(s_sum1a[14:14]),.IN2(n130),.IN3(s_sum2a[14:14]),.IN4(n41),.IN5(r0[14:14]),.IN6(n20),.Q(n352));
  AO222X1 U229(.IN1(s_sum1a[13:13]),.IN2(n130),.IN3(s_sum2a[13:13]),.IN4(n41),.IN5(r0[13:13]),.IN6(n18),.Q(n353));
  AO222X1 U230(.IN1(s_sum1a[12:12]),.IN2(n130),.IN3(s_sum2a[12:12]),.IN4(n41),.IN5(r0[12:12]),.IN6(n19),.Q(n354));
  AO222X1 U231(.IN1(s_sum1a[11:11]),.IN2(n130),.IN3(s_sum2a[11:11]),.IN4(n41),.IN5(r0[11:11]),.IN6(n20),.Q(n355));
  AO222X1 U232(.IN1(s_sum1a[10:10]),.IN2(n130),.IN3(s_sum2a[10:10]),.IN4(n41),.IN5(r0[10:10]),.IN6(n18),.Q(n356));
  AO222X1 U233(.IN1(s_sum1a[9:9]),.IN2(n130),.IN3(s_sum2a[9:9]),.IN4(n41),.IN5(r0[9:9]),.IN6(n19),.Q(n357));
  AO222X1 U234(.IN1(s_sum1a[8:8]),.IN2(n130),.IN3(s_sum2a[8:8]),.IN4(n41),.IN5(r0[8:8]),.IN6(n20),.Q(n358));
  AO222X1 U235(.IN1(s_sum1a[7:7]),.IN2(n130),.IN3(s_sum2a[7:7]),.IN4(n41),.IN5(r0[7:7]),.IN6(n18),.Q(n359));
  AO222X1 U236(.IN1(s_sum1a[6:6]),.IN2(n130),.IN3(s_sum2a[6:6]),.IN4(n41),.IN5(r0[6:6]),.IN6(n19),.Q(n360));
  AO222X1 U237(.IN1(s_sum1a[5:5]),.IN2(n130),.IN3(s_sum2a[5:5]),.IN4(n41),.IN5(r0[5:5]),.IN6(n20),.Q(n361));
  AO222X1 U238(.IN1(s_sum1a[4:4]),.IN2(n130),.IN3(s_sum2a[4:4]),.IN4(n41),.IN5(r0[4:4]),.IN6(n18),.Q(n362));
  AO222X1 U239(.IN1(s_sum1a[3:3]),.IN2(n130),.IN3(s_sum2a[3:3]),.IN4(n41),.IN5(r0[3:3]),.IN6(n20),.Q(n363));
  AO222X1 U240(.IN1(s_sum1a[2:2]),.IN2(n401),.IN3(s_sum2a[2:2]),.IN4(n42),.IN5(r0[2:2]),.IN6(n18),.Q(n364));
  AO222X1 U241(.IN1(s_sum1a[1:1]),.IN2(n401),.IN3(s_sum2a[1:1]),.IN4(n42),.IN5(r0[1:1]),.IN6(n18),.Q(n365));
  AO222X1 U242(.IN1(s_sum1a[0:0]),.IN2(n401),.IN3(s_sum2a[0:0]),.IN4(n42),.IN5(r0[0:0]),.IN6(n18),.Q(n366));
  AO222X1 U243(.IN1(s_sum1a[25:25]),.IN2(n416),.IN3(s_sum2a[25:25]),.IN4(n409),.IN5(r1[25:25]),.IN6(n23),.Q(n367));
  AO222X1 U244(.IN1(s_sum1a[24:24]),.IN2(n416),.IN3(s_sum2a[24:24]),.IN4(n409),.IN5(r1[24:24]),.IN6(n22),.Q(n368));
  AO222X1 U245(.IN1(s_sum1a[23:23]),.IN2(n416),.IN3(s_sum2a[23:23]),.IN4(n409),.IN5(r1[23:23]),.IN6(n23),.Q(n369));
  AO222X1 U246(.IN1(s_sum1a[22:22]),.IN2(n416),.IN3(s_sum2a[22:22]),.IN4(n409),.IN5(r1[22:22]),.IN6(n22),.Q(n370));
  AO222X1 U247(.IN1(s_sum1a[21:21]),.IN2(n416),.IN3(s_sum2a[21:21]),.IN4(n409),.IN5(r1[21:21]),.IN6(n23),.Q(n371));
  AO222X1 U248(.IN1(s_sum1a[20:20]),.IN2(n416),.IN3(s_sum2a[20:20]),.IN4(n409),.IN5(r1[20:20]),.IN6(n22),.Q(n372));
  AO222X1 U249(.IN1(s_sum1a[19:19]),.IN2(n416),.IN3(s_sum2a[19:19]),.IN4(n409),.IN5(r1[19:19]),.IN6(n23),.Q(n373));
  AO222X1 U250(.IN1(s_sum1a[18:18]),.IN2(n416),.IN3(s_sum2a[18:18]),.IN4(n409),.IN5(r1[18:18]),.IN6(n403),.Q(n374));
  AO222X1 U251(.IN1(s_sum1a[17:17]),.IN2(n417),.IN3(s_sum2a[17:17]),.IN4(n410),.IN5(r1[17:17]),.IN6(n22),.Q(n375));
  AO222X1 U252(.IN1(s_sum1a[16:16]),.IN2(n417),.IN3(s_sum2a[16:16]),.IN4(n410),.IN5(r1[16:16]),.IN6(n23),.Q(n376));
  AO222X1 U253(.IN1(s_sum1a[15:15]),.IN2(n417),.IN3(s_sum2a[15:15]),.IN4(n410),.IN5(r1[15:15]),.IN6(n22),.Q(n377));
  AO222X1 U254(.IN1(s_sum1a[14:14]),.IN2(n417),.IN3(s_sum2a[14:14]),.IN4(n410),.IN5(r1[14:14]),.IN6(n23),.Q(n378));
  AO222X1 U255(.IN1(s_sum1a[13:13]),.IN2(n417),.IN3(s_sum2a[13:13]),.IN4(n410),.IN5(r1[13:13]),.IN6(n22),.Q(n379));
  AO222X1 U256(.IN1(s_sum1a[12:12]),.IN2(n417),.IN3(s_sum2a[12:12]),.IN4(n410),.IN5(r1[12:12]),.IN6(n23),.Q(n380));
  AO222X1 U257(.IN1(s_sum1a[11:11]),.IN2(n417),.IN3(s_sum2a[11:11]),.IN4(n410),.IN5(r1[11:11]),.IN6(n22),.Q(n381));
  AO222X1 U258(.IN1(s_sum1a[10:10]),.IN2(n417),.IN3(s_sum2a[10:10]),.IN4(n410),.IN5(r1[10:10]),.IN6(n23),.Q(n382));
  AO222X1 U259(.IN1(s_sum1a[9:9]),.IN2(n417),.IN3(s_sum2a[9:9]),.IN4(n410),.IN5(r1[9:9]),.IN6(n22),.Q(n383));
  AO222X1 U260(.IN1(s_sum1a[8:8]),.IN2(n417),.IN3(s_sum2a[8:8]),.IN4(n410),.IN5(r1[8:8]),.IN6(n23),.Q(n384));
  AO222X1 U261(.IN1(s_sum1a[7:7]),.IN2(n417),.IN3(s_sum2a[7:7]),.IN4(n410),.IN5(r1[7:7]),.IN6(n22),.Q(n385));
  AO222X1 U262(.IN1(s_sum1a[6:6]),.IN2(n417),.IN3(s_sum2a[6:6]),.IN4(n410),.IN5(r1[6:6]),.IN6(n23),.Q(n386));
  AO222X1 U263(.IN1(s_sum1a[5:5]),.IN2(n418),.IN3(s_sum2a[5:5]),.IN4(n411),.IN5(r1[5:5]),.IN6(n22),.Q(n387));
  AO222X1 U264(.IN1(s_sum1a[4:4]),.IN2(n418),.IN3(s_sum2a[4:4]),.IN4(n411),.IN5(r1[4:4]),.IN6(n23),.Q(n388));
  AO222X1 U265(.IN1(s_sum1a[3:3]),.IN2(n418),.IN3(s_sum2a[3:3]),.IN4(n411),.IN5(r1[3:3]),.IN6(n22),.Q(n389));
  AO222X1 U266(.IN1(s_sum1a[2:2]),.IN2(n418),.IN3(s_sum2a[2:2]),.IN4(n411),.IN5(r1[2:2]),.IN6(n23),.Q(n390));
  AO222X1 U267(.IN1(s_sum1a[1:1]),.IN2(n418),.IN3(s_sum2a[1:1]),.IN4(n411),.IN5(r1[1:1]),.IN6(n22),.Q(n391));
  AO222X1 U268(.IN1(s_sum1a[0:0]),.IN2(n418),.IN3(s_sum2a[0:0]),.IN4(n411),.IN5(r1[0:0]),.IN6(n23),.Q(n392));
  AO222X1 U272(.IN1(n43),.IN2(s_sum1b[0:0]),.IN3(n36),.IN4(s_sum2b[0:0]),.IN5(r0_2[0:0]),.IN6(n18),.Q(n393));
  AND3X1 U273(.IN1(n436),.IN2(n1),.IN3(n35),.Q(n123));
  AND3X1 U275(.IN1(n35),.IN2(n1),.IN3(N142),.Q(n122));
  AO221X1 U276(.IN1(N13),.IN2(n35),.IN3(\s_count[3] ),.IN4(n18),.IN5(n128),.Q(n394));
  AO22X1 U277(.IN1(\s_count[2] ),.IN2(n18),.IN3(n129),.IN4(N12),.Q(n395));
  AO221X1 U278(.IN1(N11),.IN2(n35),.IN3(\s_count[1] ),.IN4(n19),.IN5(n128),.Q(n396));
  AO22X1 U279(.IN1(s_ready_o),.IN2(n35),.IN3(n438),.IN4(n1),.Q(n397));
  AO21X1 U281(.IN1(s_state),.IN2(n131),.IN3(n423),.Q(n398));
  AO221X1 U282(.IN1(N14),.IN2(n35),.IN3(\s_count[4] ),.IN4(n20),.IN5(n128),.Q(n399));
  AO22X1 U284(.IN1(\s_count[0] ),.IN2(n18),.IN3(n129),.IN4(n16),.Q(n400));
  NOR4X0 U288(.IN1(\s_count[0] ),.IN2(\s_count[1] ),.IN3(n132),.IN4(\s_count[2] ),.QN(n45));
  OR2X1 U289(.IN1(\s_count[4] ),.IN2(\s_count[3] ),.Q(n132));
  OR2X1 U323(.IN1(N34),.IN2(n425),.Q(N140));
  OR2X1 U324(.IN1(N33),.IN2(n425),.Q(N139));
  AND2X1 U325(.IN1(N32),.IN2(n1),.Q(N138));
  OR2X1 U326(.IN1(N31),.IN2(n425),.Q(N137));
  AND2X1 U327(.IN1(n17),.IN2(n1),.Q(N136));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_0_inj sub_185_aco(.A(r1[25:0]),.B({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,N306}),.CI(1'b0),.DIFF({N334,N333,N332,N331,N330,N329,N328,N327,N326,N325,N324,N323,N322,N321,N320,N319,N318,N317,N316,N315,N314,N313,N312,N311,N310,N309}));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW_cmp_0_inj lt_gt_163(.A(s_rad_i),.B(r0_2),.TC(1'b0),.GE_LT(1'b1),.GE_GT_EQ(1'b0),.GE_LT_GT_LE(N142));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_0_inj add_151(.A(s_op1),.B({s_op2[51:33],n444,n455,n443,n457,n441,n454,n442,n458,n440,s_op2[23:17],n439,s_op2[15:0]}),.CI(1'b0),.SUM(s_sum2b));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_1_inj sub_150(.A(s_op1),.B({s_op2[51:33],n444,n455,n443,n457,n441,n454,n442,n458,n440,s_op2[23:17],n439,s_op2[15:0]}),.CI(1'b0),.DIFF(s_sum1b));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_1_inj add_149(.A(r0[25:0]),.B(b[25:0]),.CI(1'b0),.SUM(s_sum2a));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_2_inj sub_148(.A(r0[25:0]),.B(b[25:0]),.CI(1'b0),.DIFF(s_sum1a));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_add_2_inj add_146(.A(r0_2),.B({1'b0,b_2[50:50],1'b0,b_2[48:48],1'b0,b_2[46:46],1'b0,b_2[44:44],1'b0,b_2[42:42],1'b0,b_2[40:40],1'b0,b_2[38:38],1'b0,b_2[36:36],1'b0,b_2[34:34],1'b0,b_2[32:32],1'b0,b_2[30:30],1'b0,b_2[28:28],1'b0,b_2[26:26],1'b0,b_2[24:24],1'b0,b_2[22:22],1'b0,b_2[20:20],1'b0,b_2[18:18],1'b0,b_2[16:16],1'b0,b_2[14:14],1'b0,b_2[12:12],1'b0,b_2[10:10],1'b0,b_2[8:8],1'b0,b_2[6:6],1'b0,b_2[4:4],1'b0,b_2[2:2],1'b0,b_2[0:0]}),.CI(1'b0),.SUM(s_op1));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_cmp6_0_inj r375(.A(s_rad_i),.B(r1_2),.TC(1'b0),.LT(N306),.EQ(N466));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_sub_3_inj sub_1_root_add_199(.A(r1_2),.B({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,r1[25:0],1'b0}),.CI(1'b0),.DIFF({N413,N412,N411,N410,N409,N408,N407,N406,N405,N404,N403,N402,N401,N400,N399,N398,N397,N396,N395,N394,N393,N392,N391,N390,N389,N388,N387,N386,N385,N384,N383,N382,N381,N380,N379,N378,N377,N376,N375,N374,N373,N372,N371,N370,N369,N368,N367,N366,N365,N364,N363,N362}));
  sqrt_RD_WIDTH52_SQ_WIDTH26_DW01_inc_0_inj add_0_root_add_199(.A({N413,N412,N411,N410,N409,N408,N407,N406,N405,N404,N403,N402,N401,N400,N399,N398,N397,N396,N395,N394,N393,N392,N391,N390,N389,N388,N387,N386,N385,N384,N383,N382,N381,N380,N379,N378,N377,N376,N375,N374,N373,N372,N371,N370,N369,N368,N367,N366,N365,N364,N363,N362}),.SUM({N465,N464,N463,N462,N461,N460,N459,N458,N457,N456,N455,N454,N453,N452,N451,N450,N449,N448,N447,N446,N445,N444,N443,N442,N441,N440,N439,N438,N437,N436,N435,N434,N433,N432,N431,N430,N429,N428,N427,N426,N425,N424,N423,N422,N421,N420,N419,N418,N417,N416,N415,N414}));
  DFFX1 desc2275(.D(N139),.CLK(clk_i),.Q(c[3:3]),.QN(n14));
  DFFX1 desc2276(.D(N140),.CLK(clk_i),.Q(c[4:4]),.QN(n12));
  NOR2X0 U4(.IN1(n45),.IN2(n422),.QN(n15));
  NBUFFX2 U5(.INP(n119),.Z(n418));
  NBUFFX2 U85(.INP(n119),.Z(n412));
  NBUFFX2 U112(.INP(n119),.Z(n413));
  NBUFFX2 U113(.INP(n119),.Z(n414));
  NBUFFX2 U269(.INP(n119),.Z(n415));
  NBUFFX2 U270(.INP(n119),.Z(n417));
  NBUFFX2 U271(.INP(n119),.Z(n416));
  NBUFFX2 U274(.INP(n120),.Z(n411));
  NBUFFX2 U280(.INP(n120),.Z(n405));
  NBUFFX2 U283(.INP(n120),.Z(n406));
  NBUFFX2 U285(.INP(n120),.Z(n407));
  NBUFFX2 U286(.INP(n120),.Z(n408));
  NBUFFX2 U287(.INP(n120),.Z(n410));
  NBUFFX2 U290(.INP(n120),.Z(n409));
  NBUFFX2 U291(.INP(n124),.Z(n18));
  NOR2X0 U292(.IN1(n436),.IN2(n21),.QN(n119));
  NBUFFX2 U293(.INP(n118),.Z(n419));
  NBUFFX2 U294(.INP(n118),.Z(n420));
  NBUFFX2 U295(.INP(n118),.Z(n421));
  NBUFFX2 U296(.INP(n124),.Z(n19));
  NBUFFX2 U297(.INP(n124),.Z(n20));
  NAND2X0 U298(.IN1(n497),.IN2(n28),.QN(n517));
  INVX0 U299(.INP(n511),.ZN(n459));
  INVX0 U300(.INP(n520),.ZN(n461));
  INVX0 U301(.INP(n530),.ZN(n462));
  INVX0 U302(.INP(n500),.ZN(n456));
  INVX0 U303(.INP(n516),.ZN(n446));
  INVX0 U304(.INP(n556),.ZN(n442));
  INVX0 U305(.INP(n545),.ZN(n440));
  INVX0 U306(.INP(n552),.ZN(n458));
  INVX0 U307(.INP(n551),.ZN(n463));
  INVX0 U308(.INP(n526),.ZN(n448));
  INVX0 U309(.INP(n535),.ZN(n450));
  INVX0 U310(.INP(n561),.ZN(n454));
  INVX0 U311(.INP(n566),.ZN(n441));
  INVX0 U312(.INP(n570),.ZN(n457));
  INVX0 U313(.INP(n557),.ZN(n465));
  INVX0 U314(.INP(n579),.ZN(n475));
  INVX0 U315(.INP(n575),.ZN(n443));
  INVX0 U316(.INP(n578),.ZN(n455));
  INVX0 U317(.INP(n582),.ZN(n444));
  INVX0 U318(.INP(n576),.ZN(n469));
  NOR2X0 U319(.IN1(n588),.IN2(n30),.QN(n589));
  NOR2X0 U320(.IN1(n30),.IN2(n585),.QN(n611));
  NOR2X0 U321(.IN1(n30),.IN2(n586),.QN(n612));
  NOR2X0 U322(.IN1(n30),.IN2(n593),.QN(n594));
  NOR2X0 U328(.IN1(n463),.IN2(n32),.QN(s_op2[41:41]));
  NOR2X0 U329(.IN1(n602),.IN2(n32),.QN(s_op2[42:42]));
  NOR2X0 U330(.IN1(n603),.IN2(n32),.QN(s_op2[43:43]));
  NOR2X0 U331(.IN1(n604),.IN2(n32),.QN(s_op2[44:44]));
  NOR2X0 U332(.IN1(n605),.IN2(n32),.QN(s_op2[45:45]));
  NOR2X0 U333(.IN1(n606),.IN2(n32),.QN(s_op2[46:46]));
  NOR2X0 U334(.IN1(n607),.IN2(n32),.QN(s_op2[47:47]));
  NOR2X0 U335(.IN1(n608),.IN2(n32),.QN(s_op2[48:48]));
  NBUFFX2 U336(.INP(n123),.Z(n42));
  NBUFFX2 U337(.INP(n122),.Z(n401));
  NOR2X0 U338(.IN1(n15),.IN2(n422),.QN(n118));
  NBUFFX2 U339(.INP(n123),.Z(n40));
  NBUFFX2 U340(.INP(n123),.Z(n41));
  NOR2X0 U341(.IN1(n21),.IN2(N142),.QN(n120));
  NBUFFX2 U342(.INP(n123),.Z(n39));
  NBUFFX2 U343(.INP(n123),.Z(n37));
  NBUFFX2 U344(.INP(n123),.Z(n38));
  NBUFFX2 U345(.INP(n123),.Z(n36));
  NBUFFX2 U346(.INP(n122),.Z(n127));
  NBUFFX2 U347(.INP(n122),.Z(n130));
  NBUFFX2 U348(.INP(n122),.Z(n126));
  NBUFFX2 U349(.INP(n122),.Z(n117));
  NBUFFX2 U350(.INP(n122),.Z(n125));
  NBUFFX2 U351(.INP(n122),.Z(n43));
  NBUFFX2 U352(.INP(n402),.Z(n21));
  INVX0 U353(.INP(N142),.ZN(n436));
  NOR2X0 U354(.IN1(n18),.IN2(n128),.QN(n129));
  NBUFFX2 U355(.INP(n402),.Z(n22));
  NBUFFX2 U356(.INP(n402),.Z(n23));
  NBUFFX2 U357(.INP(n17),.Z(n25));
  NBUFFX2 U358(.INP(n2),.Z(n27));
  NAND2X0 U359(.IN1(n486),.IN2(n26),.QN(n507));
  NBUFFX2 U360(.INP(n12),.Z(n34));
  NBUFFX2 U361(.INP(n13),.Z(n29));
  NOR2X0 U362(.IN1(n47),.IN2(n48),.QN(n46));
  NBUFFX2 U363(.INP(n14),.Z(n31));
  INVX0 U364(.INP(n546),.ZN(n460));
  INVX0 U365(.INP(n506),.ZN(n439));
  NOR2X0 U366(.IN1(n562),.IN2(n26),.QN(n579));
  INVX0 U367(.INP(n567),.ZN(n467));
  INVX0 U368(.INP(n558),.ZN(n472));
  NOR2X0 U369(.IN1(n30),.IN2(n590),.QN(n591));
  NOR2X0 U370(.IN1(n30),.IN2(n595),.QN(n596));
  NOR2X0 U371(.IN1(n30),.IN2(n600),.QN(n601));
  INVX0 U372(.INP(n599),.ZN(n452));
  INVX0 U424(.INP(n1),.ZN(n422));
  NAND2X1 U425(.IN1(n1),.IN2(n131),.QN(n128));
  INVX0 U426(.INP(n432),.ZN(n435));
  INVX0 U427(.INP(n427),.ZN(n430));
  INVX0 U428(.INP(n431),.ZN(n434));
  INVX0 U429(.INP(n426),.ZN(n429));
  INVX0 U430(.INP(n1),.ZN(n423));
  INVX0 U431(.INP(n1),.ZN(n424));
  INVX0 U432(.INP(n1),.ZN(n425));
  NBUFFX2 U433(.INP(n121),.Z(n404));
  NOR2X0 U434(.IN1(c[4:4]),.IN2(n505),.QN(s_op2[0:0]));
  NOR2X0 U435(.IN1(n547),.IN2(c[3:3]),.QN(n521));
  NOR2X0 U436(.IN1(n512),.IN2(c[3:3]),.QN(n571));
  NAND2X0 U437(.IN1(r0[0:0]),.IN2(n24),.QN(n479));
  INVX0 U438(.INP(n478),.ZN(n445));
  NOR2X0 U439(.IN1(n517),.IN2(c[3:3]),.QN(n598));
  NOR2X0 U440(.IN1(n522),.IN2(c[3:3]),.QN(n610));
  NOR2X0 U441(.IN1(n527),.IN2(c[3:3]),.QN(n613));
  NOR2X0 U442(.IN1(n531),.IN2(c[3:3]),.QN(n614));
  INVX0 U443(.INP(n45),.ZN(n437));
  NOR2X0 U444(.IN1(N466),.IN2(n46),.QN(n44));
  INVX0 U445(.INP(n480),.ZN(n447));
  INVX0 U446(.INP(n481),.ZN(n449));
  NOR2X0 U447(.IN1(c[4:4]),.IN2(n616),.QN(s_op2[8:8]));
  NOR2X0 U448(.IN1(c[4:4]),.IN2(n617),.QN(s_op2[9:9]));
  NOR2X0 U449(.IN1(c[4:4]),.IN2(n555),.QN(s_op2[10:10]));
  INVX0 U450(.INP(n482),.ZN(n451));
  INVX0 U451(.INP(n483),.ZN(n453));
  NOR2X0 U452(.IN1(c[4:4]),.IN2(n560),.QN(s_op2[11:11]));
  NOR2X0 U453(.IN1(c[4:4]),.IN2(n565),.QN(s_op2[12:12]));
  NOR2X0 U454(.IN1(c[4:4]),.IN2(n569),.QN(s_op2[13:13]));
  NOR2X0 U455(.IN1(c[4:4]),.IN2(n574),.QN(s_op2[14:14]));
  INVX0 U456(.INP(n494),.ZN(n466));
  INVX0 U457(.INP(n485),.ZN(n464));
  NOR2X0 U458(.IN1(c[4:4]),.IN2(n456),.QN(s_op2[15:15]));
  INVX0 U459(.INP(n503),.ZN(n468));
  INVX0 U460(.INP(n513),.ZN(n470));
  INVX0 U461(.INP(n542),.ZN(n474));
  INVX0 U462(.INP(n523),.ZN(n471));
  INVX0 U463(.INP(n532),.ZN(n473));
  NAND2X0 U464(.IN1(r0[25:25]),.IN2(c[0:0]),.QN(n562));
  NAND2X0 U465(.IN1(c[2:2]),.IN2(n568),.QN(n590));
  NAND2X0 U466(.IN1(c[1:1]),.IN2(n559),.QN(n577));
  NAND2X0 U467(.IN1(n579),.IN2(c[2:2]),.QN(n600));
  NOR2X0 U468(.IN1(n422),.IN2(s_state),.QN(n124));
  NAND2X1 U469(.IN1(s_state),.IN2(n1),.QN(n121));
  NAND2X1 U470(.IN1(s_state),.IN2(n45),.QN(n131));
  INVX0 U471(.INP(n131),.ZN(n438));
  NOR2X0 U472(.IN1(n423),.IN2(n144),.QN(N122));
  NOR2X0 U473(.IN1(n423),.IN2(n145),.QN(N124));
  NOR2X0 U474(.IN1(n423),.IN2(n146),.QN(N126));
  NOR2X0 U475(.IN1(n423),.IN2(n147),.QN(N128));
  NOR2X0 U476(.IN1(n423),.IN2(n148),.QN(N130));
  NOR2X0 U477(.IN1(n423),.IN2(n149),.QN(N132));
  NOR2X0 U478(.IN1(n423),.IN2(n150),.QN(N134));
  NOR2X0 U479(.IN1(n423),.IN2(n151),.QN(N35));
  NOR2X0 U480(.IN1(n423),.IN2(n152),.QN(N36));
  NOR2X0 U481(.IN1(n423),.IN2(n153),.QN(N37));
  NOR2X0 U482(.IN1(n423),.IN2(n154),.QN(N38));
  NOR2X0 U483(.IN1(n423),.IN2(n155),.QN(N39));
  NOR2X0 U484(.IN1(n423),.IN2(n156),.QN(N40));
  NOR2X0 U485(.IN1(n423),.IN2(n157),.QN(N41));
  NOR2X0 U486(.IN1(n424),.IN2(n141),.QN(N116));
  NOR2X0 U487(.IN1(n424),.IN2(n158),.QN(N42));
  NOR2X0 U488(.IN1(n424),.IN2(n159),.QN(N43));
  NOR2X0 U489(.IN1(n424),.IN2(n160),.QN(N44));
  NOR2X0 U490(.IN1(n424),.IN2(n161),.QN(N45));
  NOR2X0 U491(.IN1(n424),.IN2(n162),.QN(N46));
  NOR2X0 U492(.IN1(n424),.IN2(n191),.QN(N47));
  NOR2X0 U493(.IN1(n424),.IN2(n192),.QN(N48));
  NOR2X0 U494(.IN1(n424),.IN2(n193),.QN(N49));
  NOR2X0 U495(.IN1(n424),.IN2(n194),.QN(N50));
  NOR2X0 U496(.IN1(n424),.IN2(n195),.QN(N51));
  NOR2X0 U497(.IN1(n424),.IN2(n196),.QN(N52));
  NOR2X0 U498(.IN1(n424),.IN2(n197),.QN(N53));
  NOR2X0 U499(.IN1(n424),.IN2(n198),.QN(N54));
  NOR2X0 U500(.IN1(n425),.IN2(n204),.QN(N86));
  NOR2X0 U501(.IN1(n425),.IN2(n205),.QN(N88));
  NOR2X0 U502(.IN1(n425),.IN2(n206),.QN(N90));
  NOR2X0 U503(.IN1(n425),.IN2(n207),.QN(N92));
  NOR2X0 U504(.IN1(n425),.IN2(n208),.QN(N94));
  NOR2X0 U505(.IN1(n425),.IN2(n209),.QN(N96));
  NOR2X0 U506(.IN1(n425),.IN2(n210),.QN(N98));
  NOR2X0 U507(.IN1(n425),.IN2(n199),.QN(N55));
  NOR2X0 U508(.IN1(n425),.IN2(n200),.QN(N56));
  NOR2X0 U509(.IN1(n425),.IN2(n201),.QN(N57));
  NOR2X0 U510(.IN1(n425),.IN2(n202),.QN(N58));
  NOR2X0 U511(.IN1(n425),.IN2(n203),.QN(N59));
  NOR2X0 U512(.IN1(n422),.IN2(n133),.QN(N100));
  NOR2X0 U513(.IN1(n422),.IN2(n134),.QN(N102));
  NOR2X0 U514(.IN1(n422),.IN2(n135),.QN(N104));
  NOR2X0 U515(.IN1(n422),.IN2(n136),.QN(N106));
  NOR2X0 U516(.IN1(n422),.IN2(n137),.QN(N108));
  NOR2X0 U517(.IN1(n422),.IN2(n138),.QN(N110));
  NOR2X0 U518(.IN1(n422),.IN2(n139),.QN(N112));
  NOR2X0 U519(.IN1(n422),.IN2(n140),.QN(N114));
  NOR2X0 U520(.IN1(n422),.IN2(n142),.QN(N118));
  NOR2X0 U521(.IN1(n422),.IN2(n143),.QN(N120));
  NBUFFX4 U522(.INP(n17),.Z(n24));
  NBUFFX4 U523(.INP(n2),.Z(n26));
  NBUFFX4 U524(.INP(n13),.Z(n28));
  NBUFFX4 U525(.INP(n14),.Z(n30));
  NBUFFX4 U526(.INP(n12),.Z(n32));
  NBUFFX4 U527(.INP(n12),.Z(n33));
  NBUFFX2 U528(.INP(n121),.Z(n402));
  NBUFFX4 U529(.INP(n121),.Z(n403));
  INVX0 U530(.INP(n124),.ZN(n35));
  NOR2X0 U531(.IN1(\s_count[1] ),.IN2(\s_count[0] ),.QN(n426));
  AO21X1 U532(.IN1(\s_count[1] ),.IN2(\s_count[0] ),.IN3(n426),.Q(N11));
  NOR2X0 U533(.IN1(n429),.IN2(\s_count[2] ),.QN(n427));
  AO21X1 U534(.IN1(\s_count[2] ),.IN2(n429),.IN3(n427),.Q(N12));
  XNOR2X1 U535(.IN1(\s_count[3] ),.IN2(n430),.Q(N13));
  NOR2X0 U536(.IN1(\s_count[3] ),.IN2(n430),.QN(n428));
  XOR2X1 U537(.IN1(\s_count[4] ),.IN2(n428),.Q(N14));
  NOR2X0 U538(.IN1(c[1:1]),.IN2(c[0:0]),.QN(n431));
  AO21X1 U539(.IN1(c[1:1]),.IN2(c[0:0]),.IN3(n431),.Q(N31));
  NOR2X0 U540(.IN1(n434),.IN2(c[2:2]),.QN(n432));
  AO21X1 U541(.IN1(c[2:2]),.IN2(n434),.IN3(n432),.Q(N32));
  XNOR2X1 U542(.IN1(c[3:3]),.IN2(n435),.Q(N33));
  NOR2X0 U543(.IN1(c[3:3]),.IN2(n435),.QN(n433));
  XOR2X1 U544(.IN1(c[4:4]),.IN2(n433),.Q(N34));
  OR2X1 U547(.IN1(n479),.IN2(c[1:1]),.Q(n484));
  OR2X1 U548(.IN1(n484),.IN2(c[2:2]),.Q(n541));
  OR2X1 U549(.IN1(n541),.IN2(c[3:3]),.Q(n505));
  MUX21X1 U550(.IN1(r0[1:1]),.IN2(r0[2:2]),.S(n25),.Q(n478));
  MUX21X1 U551(.IN1(n479),.IN2(n445),.S(n27),.Q(n493));
  OR2X1 U552(.IN1(n493),.IN2(c[2:2]),.Q(n512));
  MUX21X1 U553(.IN1(r0[3:3]),.IN2(r0[4:4]),.S(n25),.Q(n480));
  MUX21X1 U554(.IN1(r0[5:5]),.IN2(r0[6:6]),.S(n25),.Q(n481));
  MUX21X1 U555(.IN1(n447),.IN2(n449),.S(n27),.Q(n492));
  MUX21X1 U556(.IN1(r0[7:7]),.IN2(r0[8:8]),.S(n25),.Q(n482));
  MUX21X1 U557(.IN1(r0[9:9]),.IN2(r0[10:10]),.S(n25),.Q(n483));
  MUX21X1 U558(.IN1(n451),.IN2(n453),.S(n27),.Q(n495));
  MUX21X1 U559(.IN1(n492),.IN2(n495),.S(n28),.Q(n515));
  MUX21X1 U560(.IN1(n512),.IN2(n515),.S(n30),.Q(n555));
  MUX21X1 U561(.IN1(r0[0:0]),.IN2(r0[1:1]),.S(n25),.Q(n486));
  MUX21X1 U562(.IN1(r0[2:2]),.IN2(r0[3:3]),.S(n25),.Q(n488));
  MUX21X1 U563(.IN1(n486),.IN2(n488),.S(n27),.Q(n497));
  MUX21X1 U564(.IN1(r0[4:4]),.IN2(r0[5:5]),.S(n25),.Q(n487));
  MUX21X1 U565(.IN1(r0[6:6]),.IN2(r0[7:7]),.S(n25),.Q(n490));
  MUX21X1 U566(.IN1(n487),.IN2(n490),.S(n27),.Q(n496));
  MUX21X1 U567(.IN1(r0[8:8]),.IN2(r0[9:9]),.S(n24),.Q(n489));
  MUX21X1 U568(.IN1(r0[10:10]),.IN2(r0[11:11]),.S(n24),.Q(n491));
  MUX21X1 U569(.IN1(n489),.IN2(n491),.S(n27),.Q(n499));
  MUX21X1 U570(.IN1(n496),.IN2(n499),.S(n29),.Q(n520));
  MUX21X1 U571(.IN1(n517),.IN2(n461),.S(n30),.Q(n560));
  MUX21X1 U572(.IN1(n445),.IN2(n447),.S(n27),.Q(n502));
  MUX21X1 U573(.IN1(n484),.IN2(n502),.S(n29),.Q(n522));
  MUX21X1 U574(.IN1(n449),.IN2(n451),.S(n27),.Q(n501));
  MUX21X1 U575(.IN1(r0[11:11]),.IN2(r0[12:12]),.S(n24),.Q(n485));
  MUX21X1 U576(.IN1(n453),.IN2(n464),.S(n26),.Q(n504));
  MUX21X1 U577(.IN1(n501),.IN2(n504),.S(n29),.Q(n525));
  MUX21X1 U578(.IN1(n522),.IN2(n525),.S(n31),.Q(n565));
  MUX21X1 U579(.IN1(n488),.IN2(n487),.S(n26),.Q(n511));
  MUX21X1 U580(.IN1(n507),.IN2(n459),.S(n29),.Q(n527));
  MUX21X1 U581(.IN1(n490),.IN2(n489),.S(n26),.Q(n510));
  MUX21X1 U582(.IN1(r0[12:12]),.IN2(r0[13:13]),.S(n24),.Q(n498));
  MUX21X1 U583(.IN1(n491),.IN2(n498),.S(n26),.Q(n509));
  MUX21X1 U584(.IN1(n510),.IN2(n509),.S(n29),.Q(n530));
  MUX21X1 U585(.IN1(n527),.IN2(n462),.S(n31),.Q(n569));
  MUX21X1 U586(.IN1(n493),.IN2(n492),.S(n29),.Q(n531));
  MUX21X1 U587(.IN1(r0[13:13]),.IN2(r0[14:14]),.S(n24),.Q(n494));
  MUX21X1 U588(.IN1(n464),.IN2(n466),.S(n26),.Q(n514));
  MUX21X1 U589(.IN1(n495),.IN2(n514),.S(n29),.Q(n534));
  MUX21X1 U590(.IN1(n531),.IN2(n534),.S(n31),.Q(n574));
  MUX21X1 U591(.IN1(n497),.IN2(n496),.S(n29),.Q(n536));
  MUX21X1 U592(.IN1(r0[14:14]),.IN2(r0[15:15]),.S(n24),.Q(n508));
  MUX21X1 U593(.IN1(n498),.IN2(n508),.S(n26),.Q(n519));
  MUX21X1 U594(.IN1(n499),.IN2(n519),.S(n29),.Q(n539));
  MUX21X1 U595(.IN1(n536),.IN2(n539),.S(n31),.Q(n500));
  MUX21X1 U596(.IN1(n502),.IN2(n501),.S(n28),.Q(n540));
  MUX21X1 U597(.IN1(r0[15:15]),.IN2(r0[16:16]),.S(n24),.Q(n503));
  MUX21X1 U598(.IN1(n466),.IN2(n468),.S(n26),.Q(n524));
  MUX21X1 U599(.IN1(n504),.IN2(n524),.S(n28),.Q(n544));
  MUX21X1 U600(.IN1(n540),.IN2(n544),.S(n31),.Q(n581));
  MUX21X1 U601(.IN1(n505),.IN2(n581),.S(n33),.Q(n506));
  OR2X1 U602(.IN1(n507),.IN2(c[2:2]),.Q(n547));
  MUX21X1 U603(.IN1(r0[16:16]),.IN2(r0[17:17]),.S(n24),.Q(n518));
  MUX21X1 U604(.IN1(n508),.IN2(n518),.S(n26),.Q(n529));
  MUX21X1 U605(.IN1(n509),.IN2(n529),.S(n28),.Q(n550));
  MUX21X1 U606(.IN1(n511),.IN2(n510),.S(n28),.Q(n546));
  MUX21X1 U607(.IN1(n550),.IN2(n546),.S(c[3:3]),.Q(n584));
  MUX21X1 U608(.IN1(n521),.IN2(n584),.S(n32),.Q(s_op2[17:17]));
  MUX21X1 U609(.IN1(r0[17:17]),.IN2(r0[18:18]),.S(n24),.Q(n513));
  MUX21X1 U610(.IN1(n468),.IN2(n470),.S(n26),.Q(n533));
  MUX21X1 U611(.IN1(n514),.IN2(n533),.S(n28),.Q(n554));
  MUX21X1 U612(.IN1(n515),.IN2(n554),.S(n31),.Q(n516));
  MUX21X1 U613(.IN1(n571),.IN2(n446),.S(n33),.Q(s_op2[18:18]));
  MUX21X1 U614(.IN1(r0[18:18]),.IN2(r0[19:19]),.S(n24),.Q(n528));
  MUX21X1 U615(.IN1(n518),.IN2(n528),.S(n26),.Q(n538));
  MUX21X1 U616(.IN1(n519),.IN2(n538),.S(n28),.Q(n557));
  MUX21X1 U617(.IN1(n557),.IN2(n520),.S(c[3:3]),.Q(n587));
  MUX21X1 U618(.IN1(n598),.IN2(n587),.S(n33),.Q(s_op2[19:19]));
  AND2X1 U619(.IN1(n34),.IN2(n521),.Q(s_op2[1:1]));
  MUX21X1 U620(.IN1(r0[19:19]),.IN2(r0[20:20]),.S(n24),.Q(n523));
  MUX21X1 U621(.IN1(n470),.IN2(n471),.S(n26),.Q(n543));
  MUX21X1 U622(.IN1(n524),.IN2(n543),.S(n28),.Q(n564));
  MUX21X1 U623(.IN1(n525),.IN2(n564),.S(n31),.Q(n526));
  MUX21X1 U624(.IN1(n610),.IN2(n448),.S(n33),.Q(s_op2[20:20]));
  MUX21X1 U625(.IN1(r0[20:20]),.IN2(r0[21:21]),.S(n24),.Q(n537));
  MUX21X1 U626(.IN1(n528),.IN2(n537),.S(n26),.Q(n549));
  MUX21X1 U627(.IN1(n529),.IN2(n549),.S(n28),.Q(n567));
  MUX21X1 U628(.IN1(n567),.IN2(n530),.S(c[3:3]),.Q(n592));
  MUX21X1 U629(.IN1(n613),.IN2(n592),.S(n33),.Q(s_op2[21:21]));
  MUX21X1 U630(.IN1(r0[21:21]),.IN2(r0[22:22]),.S(n24),.Q(n532));
  MUX21X1 U631(.IN1(n471),.IN2(n473),.S(n26),.Q(n553));
  MUX21X1 U632(.IN1(n533),.IN2(n553),.S(n28),.Q(n573));
  MUX21X1 U633(.IN1(n534),.IN2(n573),.S(n31),.Q(n535));
  MUX21X1 U634(.IN1(n614),.IN2(n450),.S(n33),.Q(s_op2[22:22]));
  AND2X1 U635(.IN1(n536),.IN2(n31),.Q(n615));
  MUX21X1 U636(.IN1(r0[22:22]),.IN2(r0[23:23]),.S(n24),.Q(n548));
  MUX21X1 U637(.IN1(n537),.IN2(n548),.S(n26),.Q(n558));
  MUX21X1 U638(.IN1(n538),.IN2(n558),.S(n28),.Q(n576));
  MUX21X1 U639(.IN1(n576),.IN2(n539),.S(c[3:3]),.Q(n597));
  MUX21X1 U640(.IN1(n615),.IN2(n597),.S(n33),.Q(s_op2[23:23]));
  MUX21X1 U641(.IN1(n541),.IN2(n540),.S(n31),.Q(n616));
  MUX21X1 U642(.IN1(r0[23:23]),.IN2(r0[24:24]),.S(n24),.Q(n542));
  MUX21X1 U643(.IN1(n473),.IN2(n474),.S(n26),.Q(n563));
  MUX21X1 U644(.IN1(n543),.IN2(n563),.S(n28),.Q(n580));
  MUX21X1 U645(.IN1(n544),.IN2(n580),.S(n31),.Q(n599));
  MUX21X1 U646(.IN1(n616),.IN2(n599),.S(n33),.Q(n545));
  MUX21X1 U647(.IN1(n547),.IN2(n460),.S(n31),.Q(n617));
  MUX21X1 U648(.IN1(r0[24:24]),.IN2(r0[25:25]),.S(n24),.Q(n559));
  MUX21X1 U649(.IN1(n548),.IN2(n559),.S(n26),.Q(n568));
  MUX21X1 U650(.IN1(n549),.IN2(n568),.S(n28),.Q(n583));
  MUX21X1 U651(.IN1(n550),.IN2(n583),.S(n31),.Q(n551));
  MUX21X1 U652(.IN1(n617),.IN2(n463),.S(n33),.Q(n552));
  MUX21X1 U653(.IN1(n474),.IN2(n562),.S(n26),.Q(n572));
  MUX21X1 U654(.IN1(n553),.IN2(n572),.S(n28),.Q(n585));
  MUX21X1 U655(.IN1(n554),.IN2(n585),.S(n30),.Q(n602));
  MUX21X1 U656(.IN1(n555),.IN2(n602),.S(n33),.Q(n556));
  MUX21X1 U657(.IN1(n472),.IN2(n577),.S(n28),.Q(n586));
  MUX21X1 U658(.IN1(n465),.IN2(n586),.S(n30),.Q(n603));
  MUX21X1 U659(.IN1(n560),.IN2(n603),.S(n33),.Q(n561));
  MUX21X1 U660(.IN1(n563),.IN2(n475),.S(n28),.Q(n588));
  MUX21X1 U661(.IN1(n564),.IN2(n588),.S(n30),.Q(n604));
  MUX21X1 U662(.IN1(n565),.IN2(n604),.S(n33),.Q(n566));
  MUX21X1 U663(.IN1(n467),.IN2(n590),.S(n30),.Q(n605));
  MUX21X1 U664(.IN1(n569),.IN2(n605),.S(n33),.Q(n570));
  AND2X1 U665(.IN1(n34),.IN2(n571),.Q(s_op2[2:2]));
  OR2X1 U666(.IN1(n29),.IN2(n572),.Q(n593));
  MUX21X1 U667(.IN1(n573),.IN2(n593),.S(n30),.Q(n606));
  MUX21X1 U668(.IN1(n574),.IN2(n606),.S(n33),.Q(n575));
  OR2X1 U669(.IN1(n577),.IN2(n29),.Q(n595));
  MUX21X1 U670(.IN1(n469),.IN2(n595),.S(n30),.Q(n607));
  MUX21X1 U671(.IN1(n456),.IN2(n607),.S(n33),.Q(n578));
  MUX21X1 U672(.IN1(n580),.IN2(n600),.S(n30),.Q(n608));
  MUX21X1 U673(.IN1(n581),.IN2(n608),.S(n33),.Q(n582));
  AND2X1 U674(.IN1(c[3:3]),.IN2(n583),.Q(n609));
  MUX21X1 U675(.IN1(n584),.IN2(n609),.S(n33),.Q(s_op2[33:33]));
  MUX21X1 U676(.IN1(n446),.IN2(n611),.S(n33),.Q(s_op2[34:34]));
  MUX21X1 U677(.IN1(n587),.IN2(n612),.S(n32),.Q(s_op2[35:35]));
  MUX21X1 U678(.IN1(n448),.IN2(n589),.S(n32),.Q(s_op2[36:36]));
  MUX21X1 U679(.IN1(n592),.IN2(n591),.S(n32),.Q(s_op2[37:37]));
  MUX21X1 U680(.IN1(n450),.IN2(n594),.S(n32),.Q(s_op2[38:38]));
  MUX21X1 U681(.IN1(n597),.IN2(n596),.S(n32),.Q(s_op2[39:39]));
  AND2X1 U682(.IN1(n33),.IN2(n598),.Q(s_op2[3:3]));
  MUX21X1 U683(.IN1(n452),.IN2(n601),.S(n32),.Q(s_op2[40:40]));
  AND2X1 U684(.IN1(c[4:4]),.IN2(n609),.Q(s_op2[49:49]));
  AND2X1 U685(.IN1(n33),.IN2(n610),.Q(s_op2[4:4]));
  AND2X1 U686(.IN1(c[4:4]),.IN2(n611),.Q(s_op2[50:50]));
  AND2X1 U687(.IN1(n612),.IN2(c[4:4]),.Q(s_op2[51:51]));
  AND2X1 U688(.IN1(n33),.IN2(n613),.Q(s_op2[5:5]));
  AND2X1 U689(.IN1(n34),.IN2(n614),.Q(s_op2[6:6]));
  AND2X1 U690(.IN1(n34),.IN2(n615),.Q(s_op2[7:7]));
endmodule
module post_norm_sqrt_DW01_inc_0_inj (A,SUM);
input [22:0] A ;
output [22:0] SUM ;
wire [22:2] carry ;
// instances
  HADDX1 U1_1_21(.A0(A[21:21]),.B0(carry[21:21]),.C1(carry[22:22]),.SO(SUM[21:21]));
  HADDX1 U1_1_20(.A0(A[20:20]),.B0(carry[20:20]),.C1(carry[21:21]),.SO(SUM[20:20]));
  HADDX1 U1_1_19(.A0(A[19:19]),.B0(carry[19:19]),.C1(carry[20:20]),.SO(SUM[19:19]));
  HADDX1 U1_1_18(.A0(A[18:18]),.B0(carry[18:18]),.C1(carry[19:19]),.SO(SUM[18:18]));
  HADDX1 U1_1_17(.A0(A[17:17]),.B0(carry[17:17]),.C1(carry[18:18]),.SO(SUM[17:17]));
  HADDX1 U1_1_16(.A0(A[16:16]),.B0(carry[16:16]),.C1(carry[17:17]),.SO(SUM[16:16]));
  HADDX1 U1_1_15(.A0(A[15:15]),.B0(carry[15:15]),.C1(carry[16:16]),.SO(SUM[15:15]));
  HADDX1 U1_1_14(.A0(A[14:14]),.B0(carry[14:14]),.C1(carry[15:15]),.SO(SUM[14:14]));
  HADDX1 U1_1_13(.A0(A[13:13]),.B0(carry[13:13]),.C1(carry[14:14]),.SO(SUM[13:13]));
  HADDX1 U1_1_12(.A0(A[12:12]),.B0(carry[12:12]),.C1(carry[13:13]),.SO(SUM[12:12]));
  HADDX1 U1_1_11(.A0(A[11:11]),.B0(carry[11:11]),.C1(carry[12:12]),.SO(SUM[11:11]));
  HADDX1 U1_1_10(.A0(A[10:10]),.B0(carry[10:10]),.C1(carry[11:11]),.SO(SUM[10:10]));
  HADDX1 U1_1_9(.A0(A[9:9]),.B0(carry[9:9]),.C1(carry[10:10]),.SO(SUM[9:9]));
  HADDX1 U1_1_8(.A0(A[8:8]),.B0(carry[8:8]),.C1(carry[9:9]),.SO(SUM[8:8]));
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[22:22]),.IN2(A[22:22]),.Q(SUM[22:22]));
endmodule
module post_norm_sqrt_inj (clk_i,opa_i,fract_26_i,exp_i,ine_i,rmode_i,output_o,ine_o);
input [31:0] opa_i ;
input [25:0] fract_26_i ;
input [7:0] exp_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input clk_i ;
input ine_i ;
output ine_o ;
wire s_ine_i ;
wire \s_rmode_i[1]  ;
wire N25 ;
wire N26 ;
wire N27 ;
wire N28 ;
wire N29 ;
wire N30 ;
wire N31 ;
wire N32 ;
wire N33 ;
wire N34 ;
wire N35 ;
wire N36 ;
wire N37 ;
wire N38 ;
wire N39 ;
wire N40 ;
wire N41 ;
wire N42 ;
wire N43 ;
wire N44 ;
wire N45 ;
wire N46 ;
wire N47 ;
wire N48 ;
wire N49 ;
wire N50 ;
wire N51 ;
wire N52 ;
wire N53 ;
wire N54 ;
wire N55 ;
wire N56 ;
wire N57 ;
wire N58 ;
wire N59 ;
wire N60 ;
wire N61 ;
wire N62 ;
wire N63 ;
wire N64 ;
wire N65 ;
wire N66 ;
wire N67 ;
wire N68 ;
wire N69 ;
wire N70 ;
wire N134 ;
wire n10 ;
wire n11 ;
wire n12 ;
wire n13 ;
wire n14 ;
wire n15 ;
wire n16 ;
wire n17 ;
wire n22 ;
wire n23 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n31 ;
wire n32 ;
wire n33 ;
wire n34 ;
wire n35 ;
wire n36 ;
wire n37 ;
wire n38 ;
wire n39 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n46 ;
wire n47 ;
wire n48 ;
wire n1 ;
wire n18 ;
wire n19 ;
wire n20 ;
wire n21 ;
wire n49 ;
wire n50 ;
wire [30:0] s_opa_i ;
wire [7:0] s_expa ;
wire [24:0] s_fract_26_i ;
wire [31:0] s_output_o ;
wire [22:0] s_frac_rnd ;
// instances
  DFFX1 desc2277(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_opa_i[30:30]));
  DFFX1 desc2278(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_opa_i[29:29]));
  DFFX1 desc2279(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_opa_i[28:28]));
  DFFX1 desc2280(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_opa_i[27:27]));
  DFFX1 desc2281(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_opa_i[26:26]));
  DFFX1 desc2282(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_opa_i[25:25]));
  DFFX1 desc2283(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_opa_i[24:24]));
  DFFX1 desc2284(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_opa_i[23:23]));
  DFFX1 desc2285(.D(opa_i[22:22]),.CLK(clk_i),.Q(s_opa_i[22:22]));
  DFFX1 desc2286(.D(opa_i[21:21]),.CLK(clk_i),.Q(s_opa_i[21:21]));
  DFFX1 desc2287(.D(opa_i[20:20]),.CLK(clk_i),.Q(s_opa_i[20:20]));
  DFFX1 desc2288(.D(opa_i[19:19]),.CLK(clk_i),.Q(s_opa_i[19:19]));
  DFFX1 desc2289(.D(opa_i[18:18]),.CLK(clk_i),.Q(s_opa_i[18:18]));
  DFFX1 desc2290(.D(opa_i[17:17]),.CLK(clk_i),.Q(s_opa_i[17:17]));
  DFFX1 desc2291(.D(opa_i[16:16]),.CLK(clk_i),.Q(s_opa_i[16:16]));
  DFFX1 desc2292(.D(opa_i[15:15]),.CLK(clk_i),.Q(s_opa_i[15:15]));
  DFFX1 desc2293(.D(opa_i[14:14]),.CLK(clk_i),.Q(s_opa_i[14:14]));
  DFFX1 desc2294(.D(opa_i[13:13]),.CLK(clk_i),.Q(s_opa_i[13:13]));
  DFFX1 desc2295(.D(opa_i[12:12]),.CLK(clk_i),.Q(s_opa_i[12:12]));
  DFFX1 desc2296(.D(opa_i[11:11]),.CLK(clk_i),.Q(s_opa_i[11:11]));
  DFFX1 desc2297(.D(opa_i[10:10]),.CLK(clk_i),.Q(s_opa_i[10:10]));
  DFFX1 desc2298(.D(opa_i[9:9]),.CLK(clk_i),.Q(s_opa_i[9:9]));
  DFFX1 desc2299(.D(opa_i[8:8]),.CLK(clk_i),.Q(s_opa_i[8:8]));
  DFFX1 desc2300(.D(opa_i[7:7]),.CLK(clk_i),.Q(s_opa_i[7:7]));
  DFFX1 desc2301(.D(opa_i[6:6]),.CLK(clk_i),.Q(s_opa_i[6:6]));
  DFFX1 desc2302(.D(opa_i[5:5]),.CLK(clk_i),.Q(s_opa_i[5:5]));
  DFFX1 desc2303(.D(opa_i[4:4]),.CLK(clk_i),.Q(s_opa_i[4:4]));
  DFFX1 desc2304(.D(opa_i[3:3]),.CLK(clk_i),.Q(s_opa_i[3:3]));
  DFFX1 desc2305(.D(opa_i[2:2]),.CLK(clk_i),.Q(s_opa_i[2:2]));
  DFFX1 desc2306(.D(opa_i[1:1]),.CLK(clk_i),.Q(s_opa_i[1:1]));
  DFFX1 desc2307(.D(opa_i[0:0]),.CLK(clk_i),.Q(s_opa_i[0:0]));
  DFFX1 desc2308(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_expa[7:7]));
  DFFX1 desc2309(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_expa[6:6]));
  DFFX1 desc2310(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_expa[5:5]));
  DFFX1 desc2311(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_expa[4:4]));
  DFFX1 desc2312(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_expa[3:3]));
  DFFX1 desc2313(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_expa[2:2]));
  DFFX1 desc2314(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_expa[1:1]));
  DFFX1 desc2315(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_expa[0:0]));
  DFFX1 s_sign_i_reg(.D(opa_i[31:31]),.CLK(clk_i),.Q(s_output_o[31:31]));
  DFFX1 desc2316(.D(fract_26_i[24:24]),.CLK(clk_i),.Q(s_fract_26_i[24:24]));
  DFFX1 desc2317(.D(fract_26_i[23:23]),.CLK(clk_i),.Q(s_fract_26_i[23:23]));
  DFFX1 desc2318(.D(fract_26_i[22:22]),.CLK(clk_i),.Q(s_fract_26_i[22:22]));
  DFFX1 desc2319(.D(fract_26_i[21:21]),.CLK(clk_i),.Q(s_fract_26_i[21:21]));
  DFFX1 desc2320(.D(fract_26_i[20:20]),.CLK(clk_i),.Q(s_fract_26_i[20:20]));
  DFFX1 desc2321(.D(fract_26_i[19:19]),.CLK(clk_i),.Q(s_fract_26_i[19:19]));
  DFFX1 desc2322(.D(fract_26_i[18:18]),.CLK(clk_i),.Q(s_fract_26_i[18:18]));
  DFFX1 desc2323(.D(fract_26_i[17:17]),.CLK(clk_i),.Q(s_fract_26_i[17:17]));
  DFFX1 desc2324(.D(fract_26_i[16:16]),.CLK(clk_i),.Q(s_fract_26_i[16:16]));
  DFFX1 desc2325(.D(fract_26_i[15:15]),.CLK(clk_i),.Q(s_fract_26_i[15:15]));
  DFFX1 desc2326(.D(fract_26_i[14:14]),.CLK(clk_i),.Q(s_fract_26_i[14:14]));
  DFFX1 desc2327(.D(fract_26_i[13:13]),.CLK(clk_i),.Q(s_fract_26_i[13:13]));
  DFFX1 desc2328(.D(fract_26_i[12:12]),.CLK(clk_i),.Q(s_fract_26_i[12:12]));
  DFFX1 desc2329(.D(fract_26_i[11:11]),.CLK(clk_i),.Q(s_fract_26_i[11:11]));
  DFFX1 desc2330(.D(fract_26_i[10:10]),.CLK(clk_i),.Q(s_fract_26_i[10:10]));
  DFFX1 desc2331(.D(fract_26_i[9:9]),.CLK(clk_i),.Q(s_fract_26_i[9:9]));
  DFFX1 desc2332(.D(fract_26_i[8:8]),.CLK(clk_i),.Q(s_fract_26_i[8:8]));
  DFFX1 desc2333(.D(fract_26_i[7:7]),.CLK(clk_i),.Q(s_fract_26_i[7:7]));
  DFFX1 desc2334(.D(fract_26_i[6:6]),.CLK(clk_i),.Q(s_fract_26_i[6:6]));
  DFFX1 desc2335(.D(fract_26_i[5:5]),.CLK(clk_i),.Q(s_fract_26_i[5:5]));
  DFFX1 desc2336(.D(fract_26_i[4:4]),.CLK(clk_i),.Q(s_fract_26_i[4:4]));
  DFFX1 desc2337(.D(fract_26_i[3:3]),.CLK(clk_i),.Q(s_fract_26_i[3:3]));
  DFFX1 desc2338(.D(fract_26_i[2:2]),.CLK(clk_i),.Q(s_fract_26_i[2:2]));
  DFFX1 desc2339(.D(fract_26_i[1:1]),.CLK(clk_i),.Q(s_fract_26_i[1:1]));
  DFFX1 desc2340(.D(fract_26_i[0:0]),.CLK(clk_i),.Q(s_fract_26_i[0:0]));
  DFFX1 s_ine_i_reg(.D(ine_i),.CLK(clk_i),.Q(s_ine_i));
  DFFX1 desc2341(.D(exp_i[7:7]),.CLK(clk_i),.QN(n17));
  DFFX1 desc2342(.D(exp_i[6:6]),.CLK(clk_i),.QN(n16));
  DFFX1 desc2343(.D(exp_i[5:5]),.CLK(clk_i),.QN(n15));
  DFFX1 desc2344(.D(exp_i[4:4]),.CLK(clk_i),.QN(n14));
  DFFX1 desc2345(.D(exp_i[3:3]),.CLK(clk_i),.QN(n13));
  DFFX1 desc2346(.D(exp_i[2:2]),.CLK(clk_i),.QN(n12));
  DFFX1 desc2347(.D(exp_i[1:1]),.CLK(clk_i),.QN(n11));
  DFFX1 desc2348(.D(exp_i[0:0]),.CLK(clk_i),.QN(n10));
  DFFX1 desc2349(.D(rmode_i[1:1]),.CLK(clk_i),.Q(\s_rmode_i[1] ),.QN(n22));
  DFFX1 desc2350(.D(rmode_i[0:0]),.CLK(clk_i),.QN(n23));
  DFFX1 desc2351(.D(s_output_o[31:31]),.CLK(clk_i),.Q(output_o[31:31]));
  DFFSSRX1 desc2352(.D(n21),.RSTB(1'b1),.SETB(n17),.CLK(clk_i),.Q(output_o[30:30]));
  DFFSSRX1 desc2353(.D(n21),.RSTB(1'b1),.SETB(n16),.CLK(clk_i),.Q(output_o[29:29]));
  DFFSSRX1 desc2354(.D(n21),.RSTB(1'b1),.SETB(n15),.CLK(clk_i),.Q(output_o[28:28]));
  DFFSSRX1 desc2355(.D(n21),.RSTB(1'b1),.SETB(n14),.CLK(clk_i),.Q(output_o[27:27]));
  DFFSSRX1 desc2356(.D(n21),.RSTB(1'b1),.SETB(n13),.CLK(clk_i),.Q(output_o[26:26]));
  DFFSSRX1 desc2357(.D(n21),.RSTB(1'b1),.SETB(n12),.CLK(clk_i),.Q(output_o[25:25]));
  DFFSSRX1 desc2358(.D(n21),.RSTB(1'b1),.SETB(n11),.CLK(clk_i),.Q(output_o[24:24]));
  DFFSSRX1 desc2359(.D(n21),.RSTB(1'b1),.SETB(n10),.CLK(clk_i),.Q(output_o[23:23]));
  DFFX1 ine_o_reg(.D(N134),.CLK(clk_i),.Q(ine_o));
  DFFX1 desc2360(.D(N70),.CLK(clk_i),.Q(s_frac_rnd[22:22]));
  DFFSSRX1 desc2361(.D(s_frac_rnd[22:22]),.RSTB(n50),.SETB(n20),.CLK(clk_i),.Q(output_o[22:22]));
  DFFX1 desc2362(.D(N69),.CLK(clk_i),.Q(s_frac_rnd[21:21]));
  DFFX1 desc2363(.D(s_output_o[21:21]),.CLK(clk_i),.Q(output_o[21:21]));
  DFFX1 desc2364(.D(N68),.CLK(clk_i),.Q(s_frac_rnd[20:20]));
  DFFX1 desc2365(.D(s_output_o[20:20]),.CLK(clk_i),.Q(output_o[20:20]));
  DFFX1 desc2366(.D(N67),.CLK(clk_i),.Q(s_frac_rnd[19:19]));
  DFFX1 desc2367(.D(s_output_o[19:19]),.CLK(clk_i),.Q(output_o[19:19]));
  DFFX1 desc2368(.D(N66),.CLK(clk_i),.Q(s_frac_rnd[18:18]));
  DFFX1 desc2369(.D(s_output_o[18:18]),.CLK(clk_i),.Q(output_o[18:18]));
  DFFX1 desc2370(.D(N65),.CLK(clk_i),.Q(s_frac_rnd[17:17]));
  DFFX1 desc2371(.D(s_output_o[17:17]),.CLK(clk_i),.Q(output_o[17:17]));
  DFFX1 desc2372(.D(N64),.CLK(clk_i),.Q(s_frac_rnd[16:16]));
  DFFX1 desc2373(.D(s_output_o[16:16]),.CLK(clk_i),.Q(output_o[16:16]));
  DFFX1 desc2374(.D(N63),.CLK(clk_i),.Q(s_frac_rnd[15:15]));
  DFFX1 desc2375(.D(s_output_o[15:15]),.CLK(clk_i),.Q(output_o[15:15]));
  DFFX1 desc2376(.D(N62),.CLK(clk_i),.Q(s_frac_rnd[14:14]));
  DFFX1 desc2377(.D(s_output_o[14:14]),.CLK(clk_i),.Q(output_o[14:14]));
  DFFX1 desc2378(.D(N61),.CLK(clk_i),.Q(s_frac_rnd[13:13]));
  DFFX1 desc2379(.D(s_output_o[13:13]),.CLK(clk_i),.Q(output_o[13:13]));
  DFFX1 desc2380(.D(N60),.CLK(clk_i),.Q(s_frac_rnd[12:12]));
  DFFX1 desc2381(.D(s_output_o[12:12]),.CLK(clk_i),.Q(output_o[12:12]));
  DFFX1 desc2382(.D(N59),.CLK(clk_i),.Q(s_frac_rnd[11:11]));
  DFFX1 desc2383(.D(s_output_o[11:11]),.CLK(clk_i),.Q(output_o[11:11]));
  DFFX1 desc2384(.D(N58),.CLK(clk_i),.Q(s_frac_rnd[10:10]));
  DFFX1 desc2385(.D(s_output_o[10:10]),.CLK(clk_i),.Q(output_o[10:10]));
  DFFX1 desc2386(.D(N57),.CLK(clk_i),.Q(s_frac_rnd[9:9]));
  DFFX1 desc2387(.D(s_output_o[9:9]),.CLK(clk_i),.Q(output_o[9:9]));
  DFFX1 desc2388(.D(N56),.CLK(clk_i),.Q(s_frac_rnd[8:8]));
  DFFX1 desc2389(.D(s_output_o[8:8]),.CLK(clk_i),.Q(output_o[8:8]));
  DFFX1 desc2390(.D(N55),.CLK(clk_i),.Q(s_frac_rnd[7:7]));
  DFFX1 desc2391(.D(s_output_o[7:7]),.CLK(clk_i),.Q(output_o[7:7]));
  DFFX1 desc2392(.D(N54),.CLK(clk_i),.Q(s_frac_rnd[6:6]));
  DFFX1 desc2393(.D(s_output_o[6:6]),.CLK(clk_i),.Q(output_o[6:6]));
  DFFX1 desc2394(.D(N53),.CLK(clk_i),.Q(s_frac_rnd[5:5]));
  DFFX1 desc2395(.D(s_output_o[5:5]),.CLK(clk_i),.Q(output_o[5:5]));
  DFFX1 desc2396(.D(N52),.CLK(clk_i),.Q(s_frac_rnd[4:4]));
  DFFX1 desc2397(.D(s_output_o[4:4]),.CLK(clk_i),.Q(output_o[4:4]));
  DFFX1 desc2398(.D(N51),.CLK(clk_i),.Q(s_frac_rnd[3:3]));
  DFFX1 desc2399(.D(s_output_o[3:3]),.CLK(clk_i),.Q(output_o[3:3]));
  DFFX1 desc2400(.D(N50),.CLK(clk_i),.Q(s_frac_rnd[2:2]));
  DFFX1 desc2401(.D(s_output_o[2:2]),.CLK(clk_i),.Q(output_o[2:2]));
  DFFX1 desc2402(.D(N49),.CLK(clk_i),.Q(s_frac_rnd[1:1]));
  DFFX1 desc2403(.D(s_output_o[1:1]),.CLK(clk_i),.Q(output_o[1:1]));
  DFFX1 desc2404(.D(N48),.CLK(clk_i),.Q(s_frac_rnd[0:0]));
  DFFX1 desc2405(.D(s_output_o[0:0]),.CLK(clk_i),.Q(output_o[0:0]));
  AND2X1 U22(.IN1(s_frac_rnd[9:9]),.IN2(n18),.Q(s_output_o[9:9]));
  AND2X1 U23(.IN1(s_frac_rnd[8:8]),.IN2(n1),.Q(s_output_o[8:8]));
  AND2X1 U24(.IN1(s_frac_rnd[7:7]),.IN2(n24),.Q(s_output_o[7:7]));
  AND2X1 U25(.IN1(s_frac_rnd[6:6]),.IN2(n18),.Q(s_output_o[6:6]));
  AND2X1 U26(.IN1(s_frac_rnd[5:5]),.IN2(n1),.Q(s_output_o[5:5]));
  AND2X1 U27(.IN1(s_frac_rnd[4:4]),.IN2(n24),.Q(s_output_o[4:4]));
  AND2X1 U28(.IN1(s_frac_rnd[3:3]),.IN2(n18),.Q(s_output_o[3:3]));
  AND2X1 U29(.IN1(s_frac_rnd[2:2]),.IN2(n1),.Q(s_output_o[2:2]));
  AND2X1 U30(.IN1(s_frac_rnd[21:21]),.IN2(n24),.Q(s_output_o[21:21]));
  AND2X1 U31(.IN1(s_frac_rnd[20:20]),.IN2(n18),.Q(s_output_o[20:20]));
  AND2X1 U32(.IN1(s_frac_rnd[1:1]),.IN2(n1),.Q(s_output_o[1:1]));
  AND2X1 U33(.IN1(s_frac_rnd[19:19]),.IN2(n24),.Q(s_output_o[19:19]));
  AND2X1 U34(.IN1(s_frac_rnd[18:18]),.IN2(n18),.Q(s_output_o[18:18]));
  AND2X1 U35(.IN1(s_frac_rnd[17:17]),.IN2(n1),.Q(s_output_o[17:17]));
  AND2X1 U36(.IN1(s_frac_rnd[16:16]),.IN2(n24),.Q(s_output_o[16:16]));
  AND2X1 U37(.IN1(s_frac_rnd[15:15]),.IN2(n18),.Q(s_output_o[15:15]));
  AND2X1 U38(.IN1(s_frac_rnd[14:14]),.IN2(n1),.Q(s_output_o[14:14]));
  AND2X1 U39(.IN1(s_frac_rnd[13:13]),.IN2(n24),.Q(s_output_o[13:13]));
  AND2X1 U40(.IN1(s_frac_rnd[12:12]),.IN2(n18),.Q(s_output_o[12:12]));
  AND2X1 U41(.IN1(s_frac_rnd[11:11]),.IN2(n1),.Q(s_output_o[11:11]));
  AND2X1 U42(.IN1(s_frac_rnd[10:10]),.IN2(n18),.Q(s_output_o[10:10]));
  AND2X1 U43(.IN1(s_frac_rnd[0:0]),.IN2(n1),.Q(s_output_o[0:0]));
  AO21X1 U44(.IN1(n26),.IN2(n27),.IN3(n49),.Q(n25));
  AO22X1 U45(.IN1(N47),.IN2(n19),.IN3(s_fract_26_i[24:24]),.IN4(n29),.Q(N70));
  AO22X1 U46(.IN1(N46),.IN2(n19),.IN3(s_fract_26_i[23:23]),.IN4(n29),.Q(N69));
  AO22X1 U47(.IN1(N45),.IN2(n19),.IN3(s_fract_26_i[22:22]),.IN4(n29),.Q(N68));
  AO22X1 U48(.IN1(N44),.IN2(n19),.IN3(s_fract_26_i[21:21]),.IN4(n29),.Q(N67));
  AO22X1 U49(.IN1(N43),.IN2(n19),.IN3(s_fract_26_i[20:20]),.IN4(n29),.Q(N66));
  AO22X1 U50(.IN1(N42),.IN2(n19),.IN3(s_fract_26_i[19:19]),.IN4(n29),.Q(N65));
  AO22X1 U51(.IN1(N41),.IN2(n19),.IN3(s_fract_26_i[18:18]),.IN4(n29),.Q(N64));
  AO22X1 U52(.IN1(N40),.IN2(n19),.IN3(s_fract_26_i[17:17]),.IN4(n29),.Q(N63));
  AO22X1 U53(.IN1(N39),.IN2(n19),.IN3(s_fract_26_i[16:16]),.IN4(n29),.Q(N62));
  AO22X1 U54(.IN1(N38),.IN2(n19),.IN3(s_fract_26_i[15:15]),.IN4(n29),.Q(N61));
  AO22X1 U55(.IN1(N37),.IN2(n19),.IN3(s_fract_26_i[14:14]),.IN4(n29),.Q(N60));
  AO22X1 U56(.IN1(N36),.IN2(n19),.IN3(s_fract_26_i[13:13]),.IN4(n29),.Q(N59));
  AO22X1 U57(.IN1(N35),.IN2(n19),.IN3(s_fract_26_i[12:12]),.IN4(n29),.Q(N58));
  AO22X1 U58(.IN1(N34),.IN2(n19),.IN3(s_fract_26_i[11:11]),.IN4(n29),.Q(N57));
  AO22X1 U59(.IN1(N33),.IN2(n19),.IN3(s_fract_26_i[10:10]),.IN4(n29),.Q(N56));
  AO22X1 U60(.IN1(N32),.IN2(n19),.IN3(s_fract_26_i[9:9]),.IN4(n29),.Q(N55));
  AO22X1 U61(.IN1(N31),.IN2(n19),.IN3(s_fract_26_i[8:8]),.IN4(n29),.Q(N54));
  AO22X1 U62(.IN1(N30),.IN2(n19),.IN3(s_fract_26_i[7:7]),.IN4(n29),.Q(N53));
  AO22X1 U63(.IN1(N29),.IN2(n19),.IN3(s_fract_26_i[6:6]),.IN4(n29),.Q(N52));
  AO22X1 U64(.IN1(N28),.IN2(n19),.IN3(s_fract_26_i[5:5]),.IN4(n29),.Q(N51));
  AO22X1 U65(.IN1(N27),.IN2(n19),.IN3(s_fract_26_i[4:4]),.IN4(n29),.Q(N50));
  AO22X1 U66(.IN1(N26),.IN2(n19),.IN3(s_fract_26_i[3:3]),.IN4(n29),.Q(N49));
  AO22X1 U67(.IN1(N25),.IN2(n19),.IN3(s_fract_26_i[2:2]),.IN4(n29),.Q(N48));
  NAND4X0 U68(.IN1(s_fract_26_i[1:1]),.IN2(n33),.IN3(n23),.IN4(n22),.QN(n32));
  OR3X1 U69(.IN1(s_fract_26_i[3:3]),.IN2(s_ine_i),.IN3(s_fract_26_i[0:0]),.Q(n33));
  NAND3X0 U70(.IN1(s_output_o[31:31]),.IN2(n34),.IN3(\s_rmode_i[1] ),.QN(n35));
  NOR3X0 U71(.IN1(s_fract_26_i[0:0]),.IN2(s_ine_i),.IN3(s_fract_26_i[1:1]),.QN(n30));
  AND3X1 U72(.IN1(s_ine_i),.IN2(n50),.IN3(n28),.Q(N134));
  OR4X1 U73(.IN1(s_opa_i[27:27]),.IN2(s_opa_i[26:26]),.IN3(n37),.IN4(n38),.Q(n36));
  OR4X1 U74(.IN1(s_opa_i[23:23]),.IN2(n27),.IN3(s_opa_i[25:25]),.IN4(s_opa_i[24:24]),.Q(n38));
  NAND4X0 U75(.IN1(n39),.IN2(n40),.IN3(n41),.IN4(n42),.QN(n27));
  NOR4X0 U76(.IN1(n43),.IN2(s_opa_i[4:4]),.IN3(s_opa_i[6:6]),.IN4(s_opa_i[5:5]),.QN(n42));
  OR3X1 U77(.IN1(s_opa_i[9:9]),.IN2(s_opa_i[8:8]),.IN3(s_opa_i[7:7]),.Q(n43));
  NOR4X0 U78(.IN1(n44),.IN2(s_opa_i[1:1]),.IN3(s_opa_i[21:21]),.IN4(s_opa_i[20:20]),.QN(n41));
  OR3X1 U79(.IN1(s_opa_i[3:3]),.IN2(s_opa_i[2:2]),.IN3(s_opa_i[22:22]),.Q(n44));
  NOR4X0 U80(.IN1(n45),.IN2(s_opa_i[14:14]),.IN3(s_opa_i[16:16]),.IN4(s_opa_i[15:15]),.QN(n40));
  OR3X1 U81(.IN1(s_opa_i[19:19]),.IN2(s_opa_i[18:18]),.IN3(s_opa_i[17:17]),.Q(n45));
  NOR4X0 U82(.IN1(n46),.IN2(s_opa_i[11:11]),.IN3(s_opa_i[13:13]),.IN4(s_opa_i[12:12]),.QN(n39));
  OR2X1 U83(.IN1(s_opa_i[10:10]),.IN2(s_opa_i[0:0]),.Q(n46));
  OR3X1 U84(.IN1(s_opa_i[30:30]),.IN2(s_opa_i[29:29]),.IN3(s_opa_i[28:28]),.Q(n37));
  NAND4X0 U85(.IN1(s_expa[7:7]),.IN2(s_expa[6:6]),.IN3(s_expa[5:5]),.IN4(s_expa[4:4]),.QN(n48));
  NAND4X0 U86(.IN1(s_expa[3:3]),.IN2(s_expa[2:2]),.IN3(s_expa[1:1]),.IN4(s_expa[0:0]),.QN(n47));
  post_norm_sqrt_DW01_inc_0_inj add_136(.A(s_fract_26_i[24:2]),.SUM({N47,N46,N45,N44,N43,N42,N41,N40,N39,N38,N37,N36,N35,N34,N33,N32,N31,N30,N29,N28,N27,N26,N25}));
  INVX0 U3(.INP(n24),.ZN(n21));
  INVX0 U12(.INP(n25),.ZN(n20));
  INVX0 U13(.INP(n28),.ZN(n49));
  NOR2X0 U14(.IN1(n25),.IN2(n26),.QN(n24));
  NOR2X0 U15(.IN1(n25),.IN2(n26),.QN(n1));
  NOR2X0 U16(.IN1(n25),.IN2(n26),.QN(n18));
  INVX0 U17(.INP(n29),.ZN(n19));
  INVX0 U18(.INP(n26),.ZN(n50));
  NOR2X0 U19(.IN1(n47),.IN2(n48),.QN(n26));
  OA21X1 U20(.IN1(n30),.IN2(n31),.IN3(n32),.Q(n29));
  OA21X1 U21(.IN1(s_output_o[31:31]),.IN2(n34),.IN3(n35),.Q(n31));
  NAND2X1 U87(.IN1(\s_rmode_i[1] ),.IN2(n23),.QN(n34));
  NAND2X1 U88(.IN1(s_output_o[31:31]),.IN2(n36),.QN(n28));
endmodule
module fpu_DW01_inc_0_inj (A,SUM);
input [31:0] A ;
output [31:0] SUM ;
wire [31:2] carry ;
// instances
  HADDX1 U1_1_30(.A0(A[30:30]),.B0(carry[30:30]),.C1(carry[31:31]),.SO(SUM[30:30]));
  HADDX1 U1_1_29(.A0(A[29:29]),.B0(carry[29:29]),.C1(carry[30:30]),.SO(SUM[29:29]));
  HADDX1 U1_1_28(.A0(A[28:28]),.B0(carry[28:28]),.C1(carry[29:29]),.SO(SUM[28:28]));
  HADDX1 U1_1_27(.A0(A[27:27]),.B0(carry[27:27]),.C1(carry[28:28]),.SO(SUM[27:27]));
  HADDX1 U1_1_26(.A0(A[26:26]),.B0(carry[26:26]),.C1(carry[27:27]),.SO(SUM[26:26]));
  HADDX1 U1_1_25(.A0(A[25:25]),.B0(carry[25:25]),.C1(carry[26:26]),.SO(SUM[25:25]));
  HADDX1 U1_1_24(.A0(A[24:24]),.B0(carry[24:24]),.C1(carry[25:25]),.SO(SUM[24:24]));
  HADDX1 U1_1_23(.A0(A[23:23]),.B0(carry[23:23]),.C1(carry[24:24]),.SO(SUM[23:23]));
  HADDX1 U1_1_22(.A0(A[22:22]),.B0(carry[22:22]),.C1(carry[23:23]),.SO(SUM[22:22]));
  HADDX1 U1_1_21(.A0(A[21:21]),.B0(carry[21:21]),.C1(carry[22:22]),.SO(SUM[21:21]));
  HADDX1 U1_1_20(.A0(A[20:20]),.B0(carry[20:20]),.C1(carry[21:21]),.SO(SUM[20:20]));
  HADDX1 U1_1_19(.A0(A[19:19]),.B0(carry[19:19]),.C1(carry[20:20]),.SO(SUM[19:19]));
  HADDX1 U1_1_18(.A0(A[18:18]),.B0(carry[18:18]),.C1(carry[19:19]),.SO(SUM[18:18]));
  HADDX1 U1_1_17(.A0(A[17:17]),.B0(carry[17:17]),.C1(carry[18:18]),.SO(SUM[17:17]));
  HADDX1 U1_1_16(.A0(A[16:16]),.B0(carry[16:16]),.C1(carry[17:17]),.SO(SUM[16:16]));
  HADDX1 U1_1_15(.A0(A[15:15]),.B0(carry[15:15]),.C1(carry[16:16]),.SO(SUM[15:15]));
  HADDX1 U1_1_14(.A0(A[14:14]),.B0(carry[14:14]),.C1(carry[15:15]),.SO(SUM[14:14]));
  HADDX1 U1_1_13(.A0(A[13:13]),.B0(carry[13:13]),.C1(carry[14:14]),.SO(SUM[13:13]));
  HADDX1 U1_1_12(.A0(A[12:12]),.B0(carry[12:12]),.C1(carry[13:13]),.SO(SUM[12:12]));
  HADDX1 U1_1_11(.A0(A[11:11]),.B0(carry[11:11]),.C1(carry[12:12]),.SO(SUM[11:11]));
  HADDX1 U1_1_10(.A0(A[10:10]),.B0(carry[10:10]),.C1(carry[11:11]),.SO(SUM[10:10]));
  HADDX1 U1_1_9(.A0(A[9:9]),.B0(carry[9:9]),.C1(carry[10:10]),.SO(SUM[9:9]));
  HADDX1 U1_1_8(.A0(A[8:8]),.B0(carry[8:8]),.C1(carry[9:9]),.SO(SUM[8:8]));
  HADDX1 U1_1_7(.A0(A[7:7]),.B0(carry[7:7]),.C1(carry[8:8]),.SO(SUM[7:7]));
  HADDX1 U1_1_6(.A0(A[6:6]),.B0(carry[6:6]),.C1(carry[7:7]),.SO(SUM[6:6]));
  HADDX1 U1_1_5(.A0(A[5:5]),.B0(carry[5:5]),.C1(carry[6:6]),.SO(SUM[5:5]));
  HADDX1 U1_1_4(.A0(A[4:4]),.B0(carry[4:4]),.C1(carry[5:5]),.SO(SUM[4:4]));
  HADDX1 U1_1_3(.A0(A[3:3]),.B0(carry[3:3]),.C1(carry[4:4]),.SO(SUM[3:3]));
  HADDX1 U1_1_2(.A0(A[2:2]),.B0(carry[2:2]),.C1(carry[3:3]),.SO(SUM[2:2]));
  HADDX1 U1_1_1(.A0(A[1:1]),.B0(A[0:0]),.C1(carry[2:2]),.SO(SUM[1:1]));
  INVX0 U1(.INP(A[0:0]),.ZN(SUM[0:0]));
  XOR2X1 U2(.IN1(carry[31:31]),.IN2(A[31:31]),.Q(SUM[31:31]));
endmodule
module fpu_inj (clk_i,opa_i,opb_i,fpu_op_i,rmode_i,output_o,start_i,ready_o,ine_o,overflow_o,underflow_o,div_zero_o,inf_o,zero_o,qnan_o,snan_o,p_desc1176_p_O_DFFX1pre_norm_div_,p_desc1177_p_O_DFFX1pre_norm_div_,p_desc1178_p_O_DFFX1pre_norm_div_,p_desc1179_p_O_DFFX1pre_norm_div_,p_desc1180_p_O_DFFX1pre_norm_div_,p_desc1181_p_O_DFFX1pre_norm_div_,p_desc1182_p_O_DFFX1pre_norm_div_,p_desc1183_p_O_DFFX1pre_norm_div_,p_desc1184_p_O_DFFX1pre_norm_div_,p_desc1185_p_O_DFFX1pre_norm_div_,p_desc1186_p_O_DFFX1pre_norm_div_,p_desc1187_p_O_DFFX1pre_norm_div_,p_desc1188_p_O_DFFX1pre_norm_div_,p_desc1189_p_O_DFFX1pre_norm_div_,p_desc1190_p_O_DFFX1pre_norm_div_,p_desc1191_p_O_DFFX1pre_norm_div_,p_desc1192_p_O_DFFX1pre_norm_div_,p_desc1193_p_O_DFFX1pre_norm_div_,p_desc1194_p_O_DFFX1pre_norm_div_,p_desc1195_p_O_DFFX1pre_norm_div_,p_desc1196_p_O_DFFX1pre_norm_div_,p_desc1197_p_O_DFFX1pre_norm_div_,p_desc1198_p_O_DFFX1pre_norm_div_,p_desc1199_p_O_DFFX1pre_norm_div_,p_desc1200_p_O_DFFX1pre_norm_div_,p_desc1201_p_O_DFFX1pre_norm_div_,p_desc1202_p_O_DFFX1pre_norm_div_,p_desc1203_p_O_DFFX1pre_norm_div_,p_desc1204_p_O_DFFX1pre_norm_div_,p_desc1205_p_O_DFFX1pre_norm_div_,p_desc1206_p_O_DFFX1pre_norm_div_,p_desc1207_p_O_DFFX1pre_norm_div_,p_desc1208_p_O_DFFX1pre_norm_div_,p_desc1209_p_O_DFFX1pre_norm_div_,p_desc1210_p_O_DFFX1pre_norm_div_,p_desc1211_p_O_DFFX1pre_norm_div_,p_desc1212_p_O_DFFX1pre_norm_div_,p_desc1213_p_O_DFFX1pre_norm_div_,p_desc1368_p_O_DFFX1serial_div_,p_desc1369_p_O_DFFX1serial_div_,p_desc1370_p_O_DFFX1serial_div_,p_desc1371_p_O_DFFX1serial_div_,p_desc1372_p_O_DFFX1serial_div_,p_desc1373_p_O_DFFX1serial_div_,p_desc1374_p_O_DFFX1serial_div_,p_desc1375_p_O_DFFX1serial_div_,p_desc1376_p_O_DFFX1serial_div_,p_desc1377_p_O_DFFX1serial_div_,p_desc1378_p_O_DFFX1serial_div_,p_desc1379_p_O_DFFX1serial_div_,p_desc1380_p_O_DFFX1serial_div_,p_desc1381_p_O_DFFX1serial_div_,p_desc1382_p_O_DFFX1serial_div_,p_desc1383_p_O_DFFX1serial_div_,p_desc1384_p_O_DFFX1serial_div_,p_desc1385_p_O_DFFX1serial_div_,p_desc1386_p_O_DFFX1serial_div_,p_desc1387_p_O_DFFX1serial_div_,p_desc1388_p_O_DFFX1serial_div_,p_desc1389_p_O_DFFX1serial_div_,p_desc1390_p_O_DFFX1serial_div_,p_desc1391_p_O_DFFX1serial_div_,p_desc1392_p_O_DFFX1serial_div_,p_desc1393_p_O_DFFX1serial_div_,p_desc1394_p_O_DFFX1serial_div_,p_desc1395_p_O_DFFX1serial_div_,p_desc1396_p_O_DFFX1serial_div_,p_desc1397_p_O_DFFX1serial_div_,p_desc1398_p_O_DFFX1serial_div_,p_desc1399_p_O_DFFX1serial_div_,p_desc1400_p_O_DFFX1serial_div_,p_desc1401_p_O_DFFX1serial_div_,p_desc1402_p_O_DFFX1serial_div_,p_desc1403_p_O_DFFX1serial_div_,p_desc1404_p_O_DFFX1serial_div_,p_desc1405_p_O_DFFX1serial_div_,p_desc1406_p_O_DFFX1serial_div_,p_desc1407_p_O_DFFX1serial_div_,p_desc1408_p_O_DFFX1serial_div_,p_desc1409_p_O_DFFX1serial_div_,p_desc1410_p_O_DFFX1serial_div_,p_desc1411_p_O_DFFX1serial_div_,p_desc1412_p_O_DFFX1serial_div_,p_desc1413_p_O_DFFX1serial_div_,p_desc1414_p_O_DFFX1serial_div_,p_desc1415_p_O_DFFX1serial_div_,p_desc1416_p_O_DFFX1serial_div_,p_desc1417_p_O_DFFX1serial_div_,p_desc1418_p_O_DFFX1serial_div_,p_desc1419_p_O_DFFX1serial_div_,p_desc1420_p_O_DFFX1serial_div_,p_desc1421_p_O_DFFX1serial_div_,p_desc1422_p_O_DFFX1serial_div_,p_desc1423_p_O_DFFX1serial_div_,p_desc1424_p_O_DFFX1serial_div_,p_desc1425_p_O_DFFX1serial_div_,p_desc1426_p_O_DFFX1serial_div_,p_desc1427_p_O_DFFX1serial_div_,p_desc1428_p_O_DFFX1serial_div_,p_desc1429_p_O_DFFX1serial_div_,p_desc1430_p_O_DFFX1serial_div_,p_desc1431_p_O_DFFX1serial_div_,p_desc1432_p_O_DFFX1serial_div_,p_desc1433_p_O_DFFX1serial_div_,p_desc1434_p_O_DFFX1serial_div_,p_desc1435_p_O_DFFX1serial_div_,p_desc1436_p_O_DFFX1serial_div_,p_desc1437_p_O_DFFX1serial_div_,p_desc1438_p_O_DFFX1serial_div_,p_desc1439_p_O_DFFX1serial_div_,p_desc1440_p_O_DFFX1serial_div_,p_desc1441_p_O_DFFX1serial_div_,p_desc1442_p_O_DFFX1serial_div_,p_desc1443_p_O_DFFX1serial_div_,p_desc1444_p_O_DFFX1serial_div_,p_s_start_i_reg_p_O_DFFX1serial_div_,p_s_ready_o_reg_p_O_DFFX1serial_div_,p_desc1445_p_O_DFFX1serial_div_,p_desc1446_p_O_DFFX1serial_div_,p_desc1447_p_O_DFFX1serial_div_,p_desc1448_p_O_DFFX1serial_div_,p_desc1449_p_O_DFFX1serial_div_,p_desc1450_p_O_DFFX1serial_div_,p_desc1451_p_O_DFFX1serial_div_,p_desc1452_p_O_DFFX1serial_div_,p_desc1453_p_O_DFFX1serial_div_,p_desc1454_p_O_DFFX1serial_div_,p_desc1455_p_O_DFFX1serial_div_,p_desc1456_p_O_DFFX1serial_div_,p_desc1457_p_O_DFFX1serial_div_,p_desc1458_p_O_DFFX1serial_div_,p_desc1459_p_O_DFFX1serial_div_,p_desc1460_p_O_DFFX1serial_div_,p_desc1461_p_O_DFFX1serial_div_,p_desc1462_p_O_DFFX1serial_div_,p_desc1463_p_O_DFFX1serial_div_,p_desc1464_p_O_DFFX1serial_div_,p_desc1465_p_O_DFFX1serial_div_,p_desc1466_p_O_DFFX1serial_div_,p_desc1467_p_O_DFFX1serial_div_,p_desc1468_p_O_DFFX1serial_div_,p_desc1469_p_O_DFFX1serial_div_,p_desc1470_p_O_DFFX1serial_div_,p_desc1471_p_O_DFFX1serial_div_,p_desc1472_p_O_DFFX1serial_div_,p_desc1473_p_O_DFFX1serial_div_,p_desc1474_p_O_DFFX1serial_div_,p_desc1475_p_O_DFFX1serial_div_,p_desc1476_p_O_DFFX1serial_div_,p_desc1477_p_O_DFFX1serial_div_,p_desc1478_p_O_DFFX1serial_div_,p_desc1479_p_O_DFFX1serial_div_,p_desc1480_p_O_DFFX1serial_div_,p_desc1481_p_O_DFFX1serial_div_,p_desc1482_p_O_DFFX1serial_div_,p_desc1483_p_O_DFFX1serial_div_,p_desc1484_p_O_DFFX1serial_div_,p_desc1485_p_O_DFFX1serial_div_,p_desc1486_p_O_DFFX1serial_div_,p_desc1487_p_O_DFFX1serial_div_,p_desc1488_p_O_DFFX1serial_div_,p_desc1489_p_O_DFFX1serial_div_,p_desc1490_p_O_DFFX1serial_div_,p_desc1491_p_O_DFFX1serial_div_,p_desc1492_p_O_DFFX1serial_div_,p_desc1493_p_O_DFFX1serial_div_,p_desc1494_p_O_DFFX1serial_div_,p_desc1495_p_O_DFFX1serial_div_,p_desc1496_p_O_DFFX1serial_div_,p_desc1497_p_O_DFFX1serial_div_,p_desc1498_p_O_DFFX1serial_div_,p_desc1499_p_O_DFFX1serial_div_,p_desc1500_p_O_DFFX1serial_div_,p_desc1501_p_O_DFFX1serial_div_,p_desc1502_p_O_DFFX1serial_div_,p_desc1503_p_O_DFFX1serial_div_,p_desc1504_p_O_DFFX1serial_div_,p_desc1505_p_O_DFFX1serial_div_,p_desc1506_p_O_DFFX1serial_div_,p_desc1507_p_O_DFFX1serial_div_,p_desc1508_p_O_DFFX1serial_div_,p_desc1509_p_O_DFFX1serial_div_,p_desc1510_p_O_DFFX1serial_div_,p_desc1511_p_O_DFFX1serial_div_,p_desc1512_p_O_DFFX1serial_div_,p_desc1513_p_O_DFFX1serial_div_,p_desc1514_p_O_DFFX1serial_div_,p_desc1515_p_O_DFFX1serial_div_,p_desc1516_p_O_DFFX1serial_div_,p_desc1517_p_O_DFFX1serial_div_,p_desc1518_p_O_DFFX1serial_div_,p_desc1519_p_O_DFFX1serial_div_,p_desc1520_p_O_DFFX1serial_div_,p_desc1521_p_O_DFFX1serial_div_,p_desc1522_p_O_DFFX1serial_div_,p_desc1523_p_O_DFFX1serial_div_,p_desc1524_p_O_DFFX1serial_div_,p_desc1525_p_O_DFFX1serial_div_,p_desc1526_p_O_DFFX1serial_div_,p_desc1527_p_O_DFFX1serial_div_,p_desc1528_p_O_DFFX1serial_div_,p_s_state_reg_p_O_DFFX1serial_div_,p_desc1529_p_O_DFFX1serial_div_,p_desc1530_p_O_DFFX1post_norm_div_,p_desc1531_p_O_DFFX1post_norm_div_,p_desc1532_p_O_DFFX1post_norm_div_,p_desc1533_p_O_DFFX1post_norm_div_,p_desc1534_p_O_DFFX1post_norm_div_,p_desc1535_p_O_DFFX1post_norm_div_,p_desc1536_p_O_DFFX1post_norm_div_,p_desc1537_p_O_DFFX1post_norm_div_,p_desc1538_p_O_DFFX1post_norm_div_,p_desc1539_p_O_DFFX1post_norm_div_,p_desc1540_p_O_DFFX1post_norm_div_,p_desc1541_p_O_DFFX1post_norm_div_,p_desc1542_p_O_DFFX1post_norm_div_,p_desc1543_p_O_DFFX1post_norm_div_,p_desc1544_p_O_DFFX1post_norm_div_,p_desc1545_p_O_DFFX1post_norm_div_,p_desc1546_p_O_DFFX1post_norm_div_,p_desc1547_p_O_DFFX1post_norm_div_,p_desc1548_p_O_DFFX1post_norm_div_,p_desc1549_p_O_DFFX1post_norm_div_,p_desc1550_p_O_DFFX1post_norm_div_,p_desc1551_p_O_DFFX1post_norm_div_,p_desc1552_p_O_DFFX1post_norm_div_,p_desc1553_p_O_DFFX1post_norm_div_,p_desc1554_p_O_DFFX1post_norm_div_,p_desc1555_p_O_DFFX1post_norm_div_,p_desc1556_p_O_DFFX1post_norm_div_,p_desc1557_p_O_DFFX1post_norm_div_,p_desc1558_p_O_DFFX1post_norm_div_,p_desc1559_p_O_DFFX1post_norm_div_,p_desc1560_p_O_DFFX1post_norm_div_,p_desc1561_p_O_DFFX1post_norm_div_,p_desc1562_p_O_DFFX1post_norm_div_,p_desc1563_p_O_DFFX1post_norm_div_,p_desc1564_p_O_DFFX1post_norm_div_,p_desc1565_p_O_DFFX1post_norm_div_,p_desc1566_p_O_DFFX1post_norm_div_,p_desc1567_p_O_DFFX1post_norm_div_,p_desc1568_p_O_DFFX1post_norm_div_,p_desc1569_p_O_DFFX1post_norm_div_,p_desc1570_p_O_DFFX1post_norm_div_,p_desc1571_p_O_DFFX1post_norm_div_,p_desc1572_p_O_DFFX1post_norm_div_,p_desc1573_p_O_DFFX1post_norm_div_,p_desc1574_p_O_DFFX1post_norm_div_,p_desc1575_p_O_DFFX1post_norm_div_,p_desc1576_p_O_DFFX1post_norm_div_,p_desc1577_p_O_DFFX1post_norm_div_,p_desc1578_p_O_DFFX1post_norm_div_,p_desc1579_p_O_DFFX1post_norm_div_,p_desc1580_p_O_DFFX1post_norm_div_,p_desc1581_p_O_DFFX1post_norm_div_,p_desc1582_p_O_DFFX1post_norm_div_,p_desc1583_p_O_DFFX1post_norm_div_,p_desc1584_p_O_DFFX1post_norm_div_,p_desc1585_p_O_DFFX1post_norm_div_,p_desc1586_p_O_DFFX1post_norm_div_,p_desc1587_p_O_DFFX1post_norm_div_,p_desc1588_p_O_DFFX1post_norm_div_,p_desc1589_p_O_DFFX1post_norm_div_,p_desc1590_p_O_DFFX1post_norm_div_,p_desc1591_p_O_DFFX1post_norm_div_,p_desc1592_p_O_DFFX1post_norm_div_,p_desc1593_p_O_DFFX1post_norm_div_,p_desc1594_p_O_DFFX1post_norm_div_,p_desc1595_p_O_DFFX1post_norm_div_,p_desc1596_p_O_DFFX1post_norm_div_,p_desc1597_p_O_DFFX1post_norm_div_,p_desc1598_p_O_DFFX1post_norm_div_,p_desc1599_p_O_DFFX1post_norm_div_,p_desc1600_p_O_DFFX1post_norm_div_,p_desc1601_p_O_DFFX1post_norm_div_,p_desc1602_p_O_DFFX1post_norm_div_,p_desc1603_p_O_DFFX1post_norm_div_,p_desc1604_p_O_DFFX1post_norm_div_,p_desc1605_p_O_DFFX1post_norm_div_,p_desc1606_p_O_DFFX1post_norm_div_,p_desc1607_p_O_DFFX1post_norm_div_,p_desc1608_p_O_DFFX1post_norm_div_,p_desc1609_p_O_DFFX1post_norm_div_,p_desc1610_p_O_DFFX1post_norm_div_,p_desc1611_p_O_DFFX1post_norm_div_,p_desc1612_p_O_DFFX1post_norm_div_,p_desc1613_p_O_DFFX1post_norm_div_,p_desc1614_p_O_DFFX1post_norm_div_,p_desc1615_p_O_DFFX1post_norm_div_,p_desc1616_p_O_DFFX1post_norm_div_,p_desc1617_p_O_DFFX1post_norm_div_,p_desc1618_p_O_DFFX1post_norm_div_,p_desc1619_p_O_DFFX1post_norm_div_,p_desc1620_p_O_DFFX1post_norm_div_,p_desc1621_p_O_DFFX1post_norm_div_,p_desc1622_p_O_DFFX1post_norm_div_,p_desc1623_p_O_DFFX1post_norm_div_,p_desc1624_p_O_DFFX1post_norm_div_,p_desc1625_p_O_DFFX1post_norm_div_,p_desc1626_p_O_DFFX1post_norm_div_,p_desc1627_p_O_DFFX1post_norm_div_,p_desc1628_p_O_DFFX1post_norm_div_,p_desc1629_p_O_DFFX1post_norm_div_,p_desc1630_p_O_DFFX1post_norm_div_,p_desc1631_p_O_DFFX1post_norm_div_,p_desc1632_p_O_DFFX1post_norm_div_,p_desc1633_p_O_DFFX1post_norm_div_,p_desc1634_p_O_DFFX1post_norm_div_,p_desc1635_p_O_DFFX1post_norm_div_,p_desc1636_p_O_DFFX1post_norm_div_,p_desc1637_p_O_DFFX1post_norm_div_,p_desc1638_p_O_DFFX1post_norm_div_,p_desc1639_p_O_DFFX1post_norm_div_,p_desc1640_p_O_DFFX1post_norm_div_,p_desc1641_p_O_DFFX1post_norm_div_,p_desc1642_p_O_DFFX1post_norm_div_,p_desc1643_p_O_DFFX1post_norm_div_,p_desc1644_p_O_DFFX1post_norm_div_,p_desc1645_p_O_DFFX1post_norm_div_,p_desc1646_p_O_DFFX1post_norm_div_,p_desc1647_p_O_DFFX1post_norm_div_,p_desc1648_p_O_DFFX1post_norm_div_,p_desc1649_p_O_DFFX1post_norm_div_,p_desc1650_p_O_DFFX1post_norm_div_,p_desc1651_p_O_DFFX1post_norm_div_,p_s_sign_i_reg_p_O_DFFX1post_norm_div_,p_desc1652_p_O_DFFX1post_norm_div_,p_desc1653_p_O_DFFX1post_norm_div_,p_desc1654_p_O_DFFX1post_norm_div_,p_desc1658_p_O_DFFX1post_norm_div_,p_desc1659_p_O_DFFX1post_norm_div_,p_desc1663_p_O_DFFX1post_norm_div_,p_desc1664_p_O_DFFX1post_norm_div_,p_desc1665_p_O_DFFX1post_norm_div_,p_desc1666_p_O_DFFX1post_norm_div_,p_desc1667_p_O_DFFX1post_norm_div_,p_desc1668_p_O_DFFX1post_norm_div_,p_desc1669_p_O_DFFX1post_norm_div_,p_desc1670_p_O_DFFX1post_norm_div_,p_desc1671_p_O_DFFX1post_norm_div_,p_desc1672_p_O_DFFX1post_norm_div_,p_desc1673_p_O_DFFX1post_norm_div_,p_desc1674_p_O_DFFX1post_norm_div_,p_desc1675_p_O_DFFX1post_norm_div_,p_desc1676_p_O_DFFX1post_norm_div_,p_desc1677_p_O_DFFX1post_norm_div_,p_desc1678_p_O_DFFX1post_norm_div_,p_desc1679_p_O_DFFX1post_norm_div_,p_desc1680_p_O_DFFX1post_norm_div_,p_desc1681_p_O_DFFX1post_norm_div_,p_desc1682_p_O_DFFX1post_norm_div_,p_desc1683_p_O_DFFX1post_norm_div_,p_desc1684_p_O_DFFX1post_norm_div_,p_desc1685_p_O_DFFX1post_norm_div_,p_desc1686_p_O_DFFX1post_norm_div_,p_desc1687_p_O_DFFX1post_norm_div_,p_desc1688_p_O_DFFX1post_norm_div_,p_desc1689_p_O_DFFX1post_norm_div_,p_desc1690_p_O_DFFX1post_norm_div_,p_desc1691_p_O_DFFX1post_norm_div_,p_desc1692_p_O_DFFX1post_norm_div_,p_desc1693_p_O_DFFX1post_norm_div_,p_desc1694_p_O_DFFX1post_norm_div_,p_desc1695_p_O_DFFX1post_norm_div_,p_desc1696_p_O_DFFX1post_norm_div_,p_desc1697_p_O_DFFX1post_norm_div_,p_desc1698_p_O_DFFX1post_norm_div_,p_desc1699_p_O_DFFX1post_norm_div_,p_desc1700_p_O_DFFX1post_norm_div_,p_desc1701_p_O_DFFX1post_norm_div_,p_desc1702_p_O_DFFX1post_norm_div_,p_desc1703_p_O_DFFX1post_norm_div_,p_desc1704_p_O_DFFX1post_norm_div_,p_desc1705_p_O_DFFX1post_norm_div_,p_desc1706_p_O_DFFX1post_norm_div_,p_desc1707_p_O_DFFX1post_norm_div_,p_desc1708_p_O_DFFX1post_norm_div_,p_desc1709_p_O_DFFX1post_norm_div_,p_desc1710_p_O_DFFX1post_norm_div_,p_desc1711_p_O_DFFX1post_norm_div_,p_desc1712_p_O_DFFX1post_norm_div_,p_desc1713_p_O_DFFX1post_norm_div_,p_desc1714_p_O_DFFX1post_norm_div_,p_desc1715_p_O_DFFX1post_norm_div_,p_desc1716_p_O_DFFX1post_norm_div_,p_desc1717_p_O_DFFX1post_norm_div_,p_desc1718_p_O_DFFX1post_norm_div_,p_desc1719_p_O_DFFX1post_norm_div_,p_desc1720_p_O_DFFX1post_norm_div_,p_desc1721_p_O_DFFX1post_norm_div_,p_desc1722_p_O_DFFX1post_norm_div_,p_desc1723_p_O_DFFX1post_norm_div_,p_desc1724_p_O_DFFX1post_norm_div_,p_desc1725_p_O_DFFX1post_norm_div_,p_desc1726_p_O_DFFX1post_norm_div_,p_desc1727_p_O_DFFX1post_norm_div_,p_desc1728_p_O_DFFX1post_norm_div_,p_ine_o_reg_p_O_DFFX1post_norm_div_,p_desc1729_p_O_DFFX1post_norm_div_,p_desc1737_p_O_DFFX1post_norm_div_,p_desc1738_p_O_DFFX1post_norm_div_,p_desc1739_p_O_DFFX1post_norm_div_,p_desc1740_p_O_DFFX1post_norm_div_,p_desc1741_p_O_DFFX1post_norm_div_,p_desc1742_p_O_DFFX1post_norm_div_,p_desc1743_p_O_DFFX1post_norm_div_,p_desc1744_p_O_DFFX1post_norm_div_,p_desc1745_p_O_DFFX1post_norm_div_,p_desc1746_p_O_DFFX1post_norm_div_,p_desc1747_p_O_DFFX1post_norm_div_,p_desc1748_p_O_DFFX1post_norm_div_,p_desc1749_p_O_DFFX1post_norm_div_,p_desc1750_p_O_DFFX1post_norm_div_,p_desc1751_p_O_DFFX1post_norm_div_,p_desc1752_p_O_DFFX1post_norm_div_,p_desc1753_p_O_DFFX1post_norm_div_,p_desc1754_p_O_DFFX1post_norm_div_,p_desc1755_p_O_DFFX1post_norm_div_,p_desc1756_p_O_DFFX1post_norm_div_,p_desc1757_p_O_DFFX1post_norm_div_,p_desc1758_p_O_DFFX1post_norm_div_,p_desc1849_p_O_DFFX1post_norm_div_,p_desc1850_p_O_DFFX1post_norm_div_,p_desc1851_p_O_DFFX1post_norm_div_,p_desc1852_p_O_DFFX1post_norm_div_,p_desc1853_p_O_DFFX1post_norm_div_,p_desc1854_p_O_DFFX1post_norm_div_,p_desc1855_p_O_DFFX1post_norm_div_,p_desc1856_p_O_DFFX1post_norm_div_,p_desc1857_p_O_DFFX1post_norm_div_,p_desc1858_p_O_DFFX1post_norm_div_,p_desc1859_p_O_DFFX1post_norm_div_,p_desc1860_p_O_DFFX1post_norm_div_,p_desc1861_p_O_DFFX1post_norm_div_,p_desc1862_p_O_DFFX1post_norm_div_,p_desc1863_p_O_DFFX1post_norm_div_,p_desc1864_p_O_DFFX1post_norm_div_,p_desc1865_p_O_DFFX1post_norm_div_,p_desc1866_p_O_DFFX1post_norm_div_,p_desc1867_p_O_DFFX1post_norm_div_,p_desc1868_p_O_DFFX1post_norm_div_,p_desc1869_p_O_DFFX1post_norm_div_);
input [31:0] opa_i ;
input [31:0] opb_i ;
input [2:0] fpu_op_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input clk_i ;
input start_i ;
output ready_o ;
output ine_o ;
output overflow_o ;
output underflow_o ;
output div_zero_o ;
output inf_o ;
output zero_o ;
output qnan_o ;
output snan_o ;
wire addsub_sign_o ;
wire postnorm_addsub_ine_o ;
wire mul_24_sign ;
wire s_start_i ;
wire post_norm_mul_ine ;
wire serial_div_sign ;
wire serial_div_div_zero ;
wire post_norm_div_ine ;
wire sqrt_ine_o ;
wire post_norm_sqrt_ine_o ;
wire s_ine_o ;
wire s_state ;
wire N35 ;
wire N36 ;
wire N37 ;
wire N38 ;
wire N39 ;
wire N40 ;
wire N41 ;
wire N42 ;
wire N43 ;
wire N44 ;
wire N45 ;
wire N46 ;
wire N47 ;
wire N48 ;
wire N49 ;
wire N50 ;
wire N51 ;
wire N52 ;
wire N53 ;
wire N54 ;
wire N55 ;
wire N56 ;
wire N57 ;
wire N58 ;
wire N59 ;
wire N60 ;
wire N61 ;
wire N62 ;
wire N63 ;
wire N64 ;
wire N65 ;
wire N66 ;
wire N342 ;
wire N343 ;
wire N344 ;
wire N345 ;
wire N346 ;
wire N347 ;
wire N348 ;
wire N349 ;
wire N350 ;
wire N351 ;
wire N352 ;
wire N353 ;
wire N354 ;
wire N355 ;
wire N356 ;
wire N357 ;
wire N358 ;
wire N359 ;
wire N360 ;
wire N361 ;
wire N362 ;
wire N363 ;
wire N364 ;
wire N365 ;
wire N366 ;
wire N367 ;
wire N368 ;
wire N369 ;
wire N370 ;
wire N371 ;
wire N372 ;
wire N373 ;
wire N374 ;
wire N546 ;
wire N547 ;
wire N549 ;
wire N581 ;
wire n1 ;
wire n3 ;
wire n9 ;
wire n10 ;
wire n11 ;
wire n13 ;
wire n24 ;
wire n25 ;
wire n26 ;
wire n27 ;
wire n28 ;
wire n29 ;
wire n30 ;
wire n33 ;
wire n37 ;
wire n38 ;
wire n40 ;
wire n41 ;
wire n42 ;
wire n43 ;
wire n44 ;
wire n45 ;
wire n47 ;
wire n48 ;
wire n50 ;
wire n51 ;
wire n52 ;
wire n53 ;
wire n54 ;
wire n55 ;
wire n56 ;
wire n57 ;
wire n58 ;
wire n59 ;
wire n60 ;
wire n61 ;
wire n62 ;
wire n63 ;
wire n64 ;
wire n65 ;
wire n66 ;
wire n67 ;
wire n68 ;
wire n69 ;
wire n70 ;
wire n71 ;
wire n72 ;
wire n73 ;
wire n74 ;
wire n75 ;
wire n76 ;
wire n77 ;
wire n78 ;
wire n79 ;
wire n80 ;
wire n81 ;
wire n82 ;
wire n83 ;
wire n84 ;
wire n85 ;
wire n86 ;
wire n87 ;
wire n88 ;
wire n89 ;
wire n94 ;
wire n95 ;
wire n96 ;
wire n97 ;
wire n98 ;
wire n99 ;
wire n100 ;
wire n101 ;
wire n102 ;
wire n103 ;
wire n104 ;
wire n105 ;
wire n106 ;
wire n107 ;
wire n108 ;
wire n109 ;
wire n110 ;
wire n111 ;
wire n112 ;
wire n113 ;
wire n114 ;
wire n115 ;
wire n116 ;
wire n117 ;
wire n118 ;
wire n119 ;
wire n120 ;
wire n121 ;
wire n122 ;
wire n123 ;
wire n124 ;
wire n125 ;
wire n126 ;
wire n127 ;
wire n128 ;
wire n131 ;
wire n132 ;
wire n133 ;
wire n134 ;
wire n135 ;
wire n136 ;
wire n137 ;
wire n138 ;
wire n139 ;
wire n140 ;
wire n141 ;
wire n142 ;
wire n143 ;
wire n144 ;
wire n145 ;
wire n146 ;
wire n147 ;
wire n148 ;
wire n149 ;
wire n150 ;
wire n151 ;
wire n152 ;
wire n153 ;
wire n154 ;
wire n155 ;
wire n156 ;
wire n157 ;
wire n158 ;
wire n159 ;
wire n160 ;
wire n161 ;
wire n162 ;
wire n163 ;
wire n164 ;
wire n165 ;
wire n166 ;
wire n167 ;
wire n168 ;
wire n169 ;
wire n170 ;
wire n171 ;
wire n172 ;
wire n173 ;
wire n174 ;
wire n175 ;
wire n176 ;
wire n177 ;
wire n178 ;
wire n179 ;
wire n180 ;
wire n181 ;
wire n182 ;
wire n183 ;
wire n184 ;
wire n185 ;
wire n186 ;
wire n187 ;
wire n188 ;
wire n189 ;
wire n190 ;
wire n191 ;
wire n192 ;
wire n193 ;
wire n194 ;
wire n195 ;
wire n196 ;
wire n197 ;
wire n198 ;
wire n199 ;
wire n200 ;
wire n201 ;
wire n202 ;
wire n203 ;
wire n204 ;
wire n205 ;
wire n206 ;
wire n207 ;
wire n208 ;
wire n209 ;
wire n210 ;
wire n211 ;
wire n212 ;
wire n213 ;
wire n214 ;
wire n215 ;
wire n216 ;
wire n217 ;
wire n218 ;
wire n219 ;
wire n220 ;
wire n221 ;
wire n222 ;
wire n223 ;
wire n224 ;
wire n225 ;
wire n226 ;
wire n227 ;
wire n228 ;
wire n229 ;
wire n230 ;
wire n231 ;
wire n232 ;
wire n233 ;
wire n234 ;
wire n235 ;
wire n236 ;
wire n237 ;
wire n238 ;
wire n239 ;
wire n240 ;
wire n241 ;
wire n242 ;
wire n243 ;
wire n244 ;
wire n245 ;
wire n246 ;
wire n247 ;
wire n248 ;
wire n249 ;
wire n250 ;
wire n251 ;
wire n252 ;
wire n253 ;
wire n254 ;
wire n255 ;
wire n256 ;
wire n257 ;
wire n258 ;
wire n259 ;
wire n260 ;
wire n261 ;
wire n262 ;
wire n263 ;
wire n264 ;
wire n265 ;
wire n266 ;
wire n267 ;
wire n268 ;
wire n269 ;
wire n270 ;
wire n271 ;
wire n272 ;
wire n273 ;
wire n274 ;
wire n275 ;
wire n276 ;
wire [31:0] s_opa_i ;
wire [31:0] s_opb_i ;
wire [27:0] prenorm_addsub_fracta_28_o ;
wire [27:0] prenorm_addsub_fractb_28_o ;
wire [7:0] prenorm_addsub_exp_o ;
wire [2:0] s_fpu_op_i ;
wire [27:0] addsub_fract_o ;
wire [1:0] s_rmode_i ;
wire [31:0] postnorm_addsub_output_o ;
wire [9:0] pre_norm_mul_exp_10 ;
wire [23:0] pre_norm_mul_fracta_24 ;
wire [23:0] pre_norm_mul_fractb_24 ;
wire [47:0] mul_24_fract_48 ;
wire [31:0] post_norm_mul_output ;
wire [9:0] pre_norm_div_exp ;
wire [49:0] pre_norm_div_dvdnd ;
wire [26:0] pre_norm_div_dvsor ;
wire [26:0] serial_div_qutnt ;
wire [26:0] serial_div_rmndr ;
wire [31:0] post_norm_div_output ;
wire [51:0] pre_norm_sqrt_fracta_o ;
wire [7:0] pre_norm_sqrt_exp_o ;
wire [25:0] sqrt_sqr_o ;
wire [31:0] post_norm_sqrt_output ;
wire [31:0] s_output_o ;
wire [31:0] s_count ;
wire [31:0] s_output1 ;
wire SYNOPSYS_UNCONNECTED__0 ;
wire SYNOPSYS_UNCONNECTED__1 ;
wire SYNOPSYS_UNCONNECTED__2 ;
wire SYNOPSYS_UNCONNECTED__3 ;
wire SYNOPSYS_UNCONNECTED__4 ;
wire SYNOPSYS_UNCONNECTED__5 ;
wire SYNOPSYS_UNCONNECTED__6 ;
wire SYNOPSYS_UNCONNECTED__7 ;
wire SYNOPSYS_UNCONNECTED__8 ;
wire SYNOPSYS_UNCONNECTED__9 ;
wire SYNOPSYS_UNCONNECTED__10 ;
wire SYNOPSYS_UNCONNECTED__11 ;
wire SYNOPSYS_UNCONNECTED__12 ;
wire SYNOPSYS_UNCONNECTED__13 ;
wire SYNOPSYS_UNCONNECTED__14 ;
wire SYNOPSYS_UNCONNECTED__15 ;
wire SYNOPSYS_UNCONNECTED__16 ;
wire SYNOPSYS_UNCONNECTED__17 ;
wire SYNOPSYS_UNCONNECTED__18 ;
wire SYNOPSYS_UNCONNECTED__19 ;
wire SYNOPSYS_UNCONNECTED__20 ;
wire SYNOPSYS_UNCONNECTED__21 ;
wire SYNOPSYS_UNCONNECTED__22 ;
wire SYNOPSYS_UNCONNECTED__23 ;
wire SYNOPSYS_UNCONNECTED__24 ;
wire SYNOPSYS_UNCONNECTED__25 ;
wire SYNOPSYS_UNCONNECTED__26 ;
wire SYNOPSYS_UNCONNECTED__27 ;
wire SYNOPSYS_UNCONNECTED__28 ;
wire SYNOPSYS_UNCONNECTED__29 ;
wire SYNOPSYS_UNCONNECTED__30 ;
wire SYNOPSYS_UNCONNECTED__31 ;
wire SYNOPSYS_UNCONNECTED__32 ;
wire SYNOPSYS_UNCONNECTED__33 ;
wire SYNOPSYS_UNCONNECTED__34 ;
wire SYNOPSYS_UNCONNECTED__35 ;
wire SYNOPSYS_UNCONNECTED__36 ;
wire SYNOPSYS_UNCONNECTED__37 ;
wire SYNOPSYS_UNCONNECTED__38 ;
wire SYNOPSYS_UNCONNECTED__39 ;
wire SYNOPSYS_UNCONNECTED__40 ;
wire SYNOPSYS_UNCONNECTED__41 ;
wire SYNOPSYS_UNCONNECTED__42 ;
wire SYNOPSYS_UNCONNECTED__43 ;
wire SYNOPSYS_UNCONNECTED__44 ;
wire SYNOPSYS_UNCONNECTED__45 ;
wire SYNOPSYS_UNCONNECTED__46 ;
wire SYNOPSYS_UNCONNECTED__47 ;
wire SYNOPSYS_UNCONNECTED__48 ;
wire SYNOPSYS_UNCONNECTED__49 ;
wire SYNOPSYS_UNCONNECTED__50 ;
wire SYNOPSYS_UNCONNECTED__51 ;
wire SYNOPSYS_UNCONNECTED__52 ;
wire SYNOPSYS_UNCONNECTED__53 ;
wire SYNOPSYS_UNCONNECTED__54 ;
wire SYNOPSYS_UNCONNECTED__55 ;
wire SYNOPSYS_UNCONNECTED__56 ;
wire SYNOPSYS_UNCONNECTED__57 ;
input p_desc1176_p_O_DFFX1pre_norm_div_ ;
input p_desc1177_p_O_DFFX1pre_norm_div_ ;
input p_desc1178_p_O_DFFX1pre_norm_div_ ;
input p_desc1179_p_O_DFFX1pre_norm_div_ ;
input p_desc1180_p_O_DFFX1pre_norm_div_ ;
input p_desc1181_p_O_DFFX1pre_norm_div_ ;
input p_desc1182_p_O_DFFX1pre_norm_div_ ;
input p_desc1183_p_O_DFFX1pre_norm_div_ ;
input p_desc1184_p_O_DFFX1pre_norm_div_ ;
input p_desc1185_p_O_DFFX1pre_norm_div_ ;
input p_desc1186_p_O_DFFX1pre_norm_div_ ;
input p_desc1187_p_O_DFFX1pre_norm_div_ ;
input p_desc1188_p_O_DFFX1pre_norm_div_ ;
input p_desc1189_p_O_DFFX1pre_norm_div_ ;
input p_desc1190_p_O_DFFX1pre_norm_div_ ;
input p_desc1191_p_O_DFFX1pre_norm_div_ ;
input p_desc1192_p_O_DFFX1pre_norm_div_ ;
input p_desc1193_p_O_DFFX1pre_norm_div_ ;
input p_desc1194_p_O_DFFX1pre_norm_div_ ;
input p_desc1195_p_O_DFFX1pre_norm_div_ ;
input p_desc1196_p_O_DFFX1pre_norm_div_ ;
input p_desc1197_p_O_DFFX1pre_norm_div_ ;
input p_desc1198_p_O_DFFX1pre_norm_div_ ;
input p_desc1199_p_O_DFFX1pre_norm_div_ ;
input p_desc1200_p_O_DFFX1pre_norm_div_ ;
input p_desc1201_p_O_DFFX1pre_norm_div_ ;
input p_desc1202_p_O_DFFX1pre_norm_div_ ;
input p_desc1203_p_O_DFFX1pre_norm_div_ ;
input p_desc1204_p_O_DFFX1pre_norm_div_ ;
input p_desc1205_p_O_DFFX1pre_norm_div_ ;
input p_desc1206_p_O_DFFX1pre_norm_div_ ;
input p_desc1207_p_O_DFFX1pre_norm_div_ ;
input p_desc1208_p_O_DFFX1pre_norm_div_ ;
input p_desc1209_p_O_DFFX1pre_norm_div_ ;
input p_desc1210_p_O_DFFX1pre_norm_div_ ;
input p_desc1211_p_O_DFFX1pre_norm_div_ ;
input p_desc1212_p_O_DFFX1pre_norm_div_ ;
input p_desc1213_p_O_DFFX1pre_norm_div_ ;
input p_desc1368_p_O_DFFX1serial_div_ ;
input p_desc1369_p_O_DFFX1serial_div_ ;
input p_desc1370_p_O_DFFX1serial_div_ ;
input p_desc1371_p_O_DFFX1serial_div_ ;
input p_desc1372_p_O_DFFX1serial_div_ ;
input p_desc1373_p_O_DFFX1serial_div_ ;
input p_desc1374_p_O_DFFX1serial_div_ ;
input p_desc1375_p_O_DFFX1serial_div_ ;
input p_desc1376_p_O_DFFX1serial_div_ ;
input p_desc1377_p_O_DFFX1serial_div_ ;
input p_desc1378_p_O_DFFX1serial_div_ ;
input p_desc1379_p_O_DFFX1serial_div_ ;
input p_desc1380_p_O_DFFX1serial_div_ ;
input p_desc1381_p_O_DFFX1serial_div_ ;
input p_desc1382_p_O_DFFX1serial_div_ ;
input p_desc1383_p_O_DFFX1serial_div_ ;
input p_desc1384_p_O_DFFX1serial_div_ ;
input p_desc1385_p_O_DFFX1serial_div_ ;
input p_desc1386_p_O_DFFX1serial_div_ ;
input p_desc1387_p_O_DFFX1serial_div_ ;
input p_desc1388_p_O_DFFX1serial_div_ ;
input p_desc1389_p_O_DFFX1serial_div_ ;
input p_desc1390_p_O_DFFX1serial_div_ ;
input p_desc1391_p_O_DFFX1serial_div_ ;
input p_desc1392_p_O_DFFX1serial_div_ ;
input p_desc1393_p_O_DFFX1serial_div_ ;
input p_desc1394_p_O_DFFX1serial_div_ ;
input p_desc1395_p_O_DFFX1serial_div_ ;
input p_desc1396_p_O_DFFX1serial_div_ ;
input p_desc1397_p_O_DFFX1serial_div_ ;
input p_desc1398_p_O_DFFX1serial_div_ ;
input p_desc1399_p_O_DFFX1serial_div_ ;
input p_desc1400_p_O_DFFX1serial_div_ ;
input p_desc1401_p_O_DFFX1serial_div_ ;
input p_desc1402_p_O_DFFX1serial_div_ ;
input p_desc1403_p_O_DFFX1serial_div_ ;
input p_desc1404_p_O_DFFX1serial_div_ ;
input p_desc1405_p_O_DFFX1serial_div_ ;
input p_desc1406_p_O_DFFX1serial_div_ ;
input p_desc1407_p_O_DFFX1serial_div_ ;
input p_desc1408_p_O_DFFX1serial_div_ ;
input p_desc1409_p_O_DFFX1serial_div_ ;
input p_desc1410_p_O_DFFX1serial_div_ ;
input p_desc1411_p_O_DFFX1serial_div_ ;
input p_desc1412_p_O_DFFX1serial_div_ ;
input p_desc1413_p_O_DFFX1serial_div_ ;
input p_desc1414_p_O_DFFX1serial_div_ ;
input p_desc1415_p_O_DFFX1serial_div_ ;
input p_desc1416_p_O_DFFX1serial_div_ ;
input p_desc1417_p_O_DFFX1serial_div_ ;
input p_desc1418_p_O_DFFX1serial_div_ ;
input p_desc1419_p_O_DFFX1serial_div_ ;
input p_desc1420_p_O_DFFX1serial_div_ ;
input p_desc1421_p_O_DFFX1serial_div_ ;
input p_desc1422_p_O_DFFX1serial_div_ ;
input p_desc1423_p_O_DFFX1serial_div_ ;
input p_desc1424_p_O_DFFX1serial_div_ ;
input p_desc1425_p_O_DFFX1serial_div_ ;
input p_desc1426_p_O_DFFX1serial_div_ ;
input p_desc1427_p_O_DFFX1serial_div_ ;
input p_desc1428_p_O_DFFX1serial_div_ ;
input p_desc1429_p_O_DFFX1serial_div_ ;
input p_desc1430_p_O_DFFX1serial_div_ ;
input p_desc1431_p_O_DFFX1serial_div_ ;
input p_desc1432_p_O_DFFX1serial_div_ ;
input p_desc1433_p_O_DFFX1serial_div_ ;
input p_desc1434_p_O_DFFX1serial_div_ ;
input p_desc1435_p_O_DFFX1serial_div_ ;
input p_desc1436_p_O_DFFX1serial_div_ ;
input p_desc1437_p_O_DFFX1serial_div_ ;
input p_desc1438_p_O_DFFX1serial_div_ ;
input p_desc1439_p_O_DFFX1serial_div_ ;
input p_desc1440_p_O_DFFX1serial_div_ ;
input p_desc1441_p_O_DFFX1serial_div_ ;
input p_desc1442_p_O_DFFX1serial_div_ ;
input p_desc1443_p_O_DFFX1serial_div_ ;
input p_desc1444_p_O_DFFX1serial_div_ ;
input p_s_start_i_reg_p_O_DFFX1serial_div_ ;
input p_s_ready_o_reg_p_O_DFFX1serial_div_ ;
input p_desc1445_p_O_DFFX1serial_div_ ;
input p_desc1446_p_O_DFFX1serial_div_ ;
input p_desc1447_p_O_DFFX1serial_div_ ;
input p_desc1448_p_O_DFFX1serial_div_ ;
input p_desc1449_p_O_DFFX1serial_div_ ;
input p_desc1450_p_O_DFFX1serial_div_ ;
input p_desc1451_p_O_DFFX1serial_div_ ;
input p_desc1452_p_O_DFFX1serial_div_ ;
input p_desc1453_p_O_DFFX1serial_div_ ;
input p_desc1454_p_O_DFFX1serial_div_ ;
input p_desc1455_p_O_DFFX1serial_div_ ;
input p_desc1456_p_O_DFFX1serial_div_ ;
input p_desc1457_p_O_DFFX1serial_div_ ;
input p_desc1458_p_O_DFFX1serial_div_ ;
input p_desc1459_p_O_DFFX1serial_div_ ;
input p_desc1460_p_O_DFFX1serial_div_ ;
input p_desc1461_p_O_DFFX1serial_div_ ;
input p_desc1462_p_O_DFFX1serial_div_ ;
input p_desc1463_p_O_DFFX1serial_div_ ;
input p_desc1464_p_O_DFFX1serial_div_ ;
input p_desc1465_p_O_DFFX1serial_div_ ;
input p_desc1466_p_O_DFFX1serial_div_ ;
input p_desc1467_p_O_DFFX1serial_div_ ;
input p_desc1468_p_O_DFFX1serial_div_ ;
input p_desc1469_p_O_DFFX1serial_div_ ;
input p_desc1470_p_O_DFFX1serial_div_ ;
input p_desc1471_p_O_DFFX1serial_div_ ;
input p_desc1472_p_O_DFFX1serial_div_ ;
input p_desc1473_p_O_DFFX1serial_div_ ;
input p_desc1474_p_O_DFFX1serial_div_ ;
input p_desc1475_p_O_DFFX1serial_div_ ;
input p_desc1476_p_O_DFFX1serial_div_ ;
input p_desc1477_p_O_DFFX1serial_div_ ;
input p_desc1478_p_O_DFFX1serial_div_ ;
input p_desc1479_p_O_DFFX1serial_div_ ;
input p_desc1480_p_O_DFFX1serial_div_ ;
input p_desc1481_p_O_DFFX1serial_div_ ;
input p_desc1482_p_O_DFFX1serial_div_ ;
input p_desc1483_p_O_DFFX1serial_div_ ;
input p_desc1484_p_O_DFFX1serial_div_ ;
input p_desc1485_p_O_DFFX1serial_div_ ;
input p_desc1486_p_O_DFFX1serial_div_ ;
input p_desc1487_p_O_DFFX1serial_div_ ;
input p_desc1488_p_O_DFFX1serial_div_ ;
input p_desc1489_p_O_DFFX1serial_div_ ;
input p_desc1490_p_O_DFFX1serial_div_ ;
input p_desc1491_p_O_DFFX1serial_div_ ;
input p_desc1492_p_O_DFFX1serial_div_ ;
input p_desc1493_p_O_DFFX1serial_div_ ;
input p_desc1494_p_O_DFFX1serial_div_ ;
input p_desc1495_p_O_DFFX1serial_div_ ;
input p_desc1496_p_O_DFFX1serial_div_ ;
input p_desc1497_p_O_DFFX1serial_div_ ;
input p_desc1498_p_O_DFFX1serial_div_ ;
input p_desc1499_p_O_DFFX1serial_div_ ;
input p_desc1500_p_O_DFFX1serial_div_ ;
input p_desc1501_p_O_DFFX1serial_div_ ;
input p_desc1502_p_O_DFFX1serial_div_ ;
input p_desc1503_p_O_DFFX1serial_div_ ;
input p_desc1504_p_O_DFFX1serial_div_ ;
input p_desc1505_p_O_DFFX1serial_div_ ;
input p_desc1506_p_O_DFFX1serial_div_ ;
input p_desc1507_p_O_DFFX1serial_div_ ;
input p_desc1508_p_O_DFFX1serial_div_ ;
input p_desc1509_p_O_DFFX1serial_div_ ;
input p_desc1510_p_O_DFFX1serial_div_ ;
input p_desc1511_p_O_DFFX1serial_div_ ;
input p_desc1512_p_O_DFFX1serial_div_ ;
input p_desc1513_p_O_DFFX1serial_div_ ;
input p_desc1514_p_O_DFFX1serial_div_ ;
input p_desc1515_p_O_DFFX1serial_div_ ;
input p_desc1516_p_O_DFFX1serial_div_ ;
input p_desc1517_p_O_DFFX1serial_div_ ;
input p_desc1518_p_O_DFFX1serial_div_ ;
input p_desc1519_p_O_DFFX1serial_div_ ;
input p_desc1520_p_O_DFFX1serial_div_ ;
input p_desc1521_p_O_DFFX1serial_div_ ;
input p_desc1522_p_O_DFFX1serial_div_ ;
input p_desc1523_p_O_DFFX1serial_div_ ;
input p_desc1524_p_O_DFFX1serial_div_ ;
input p_desc1525_p_O_DFFX1serial_div_ ;
input p_desc1526_p_O_DFFX1serial_div_ ;
input p_desc1527_p_O_DFFX1serial_div_ ;
input p_desc1528_p_O_DFFX1serial_div_ ;
input p_s_state_reg_p_O_DFFX1serial_div_ ;
input p_desc1529_p_O_DFFX1serial_div_ ;
input p_desc1530_p_O_DFFX1post_norm_div_ ;
input p_desc1531_p_O_DFFX1post_norm_div_ ;
input p_desc1532_p_O_DFFX1post_norm_div_ ;
input p_desc1533_p_O_DFFX1post_norm_div_ ;
input p_desc1534_p_O_DFFX1post_norm_div_ ;
input p_desc1535_p_O_DFFX1post_norm_div_ ;
input p_desc1536_p_O_DFFX1post_norm_div_ ;
input p_desc1537_p_O_DFFX1post_norm_div_ ;
input p_desc1538_p_O_DFFX1post_norm_div_ ;
input p_desc1539_p_O_DFFX1post_norm_div_ ;
input p_desc1540_p_O_DFFX1post_norm_div_ ;
input p_desc1541_p_O_DFFX1post_norm_div_ ;
input p_desc1542_p_O_DFFX1post_norm_div_ ;
input p_desc1543_p_O_DFFX1post_norm_div_ ;
input p_desc1544_p_O_DFFX1post_norm_div_ ;
input p_desc1545_p_O_DFFX1post_norm_div_ ;
input p_desc1546_p_O_DFFX1post_norm_div_ ;
input p_desc1547_p_O_DFFX1post_norm_div_ ;
input p_desc1548_p_O_DFFX1post_norm_div_ ;
input p_desc1549_p_O_DFFX1post_norm_div_ ;
input p_desc1550_p_O_DFFX1post_norm_div_ ;
input p_desc1551_p_O_DFFX1post_norm_div_ ;
input p_desc1552_p_O_DFFX1post_norm_div_ ;
input p_desc1553_p_O_DFFX1post_norm_div_ ;
input p_desc1554_p_O_DFFX1post_norm_div_ ;
input p_desc1555_p_O_DFFX1post_norm_div_ ;
input p_desc1556_p_O_DFFX1post_norm_div_ ;
input p_desc1557_p_O_DFFX1post_norm_div_ ;
input p_desc1558_p_O_DFFX1post_norm_div_ ;
input p_desc1559_p_O_DFFX1post_norm_div_ ;
input p_desc1560_p_O_DFFX1post_norm_div_ ;
input p_desc1561_p_O_DFFX1post_norm_div_ ;
input p_desc1562_p_O_DFFX1post_norm_div_ ;
input p_desc1563_p_O_DFFX1post_norm_div_ ;
input p_desc1564_p_O_DFFX1post_norm_div_ ;
input p_desc1565_p_O_DFFX1post_norm_div_ ;
input p_desc1566_p_O_DFFX1post_norm_div_ ;
input p_desc1567_p_O_DFFX1post_norm_div_ ;
input p_desc1568_p_O_DFFX1post_norm_div_ ;
input p_desc1569_p_O_DFFX1post_norm_div_ ;
input p_desc1570_p_O_DFFX1post_norm_div_ ;
input p_desc1571_p_O_DFFX1post_norm_div_ ;
input p_desc1572_p_O_DFFX1post_norm_div_ ;
input p_desc1573_p_O_DFFX1post_norm_div_ ;
input p_desc1574_p_O_DFFX1post_norm_div_ ;
input p_desc1575_p_O_DFFX1post_norm_div_ ;
input p_desc1576_p_O_DFFX1post_norm_div_ ;
input p_desc1577_p_O_DFFX1post_norm_div_ ;
input p_desc1578_p_O_DFFX1post_norm_div_ ;
input p_desc1579_p_O_DFFX1post_norm_div_ ;
input p_desc1580_p_O_DFFX1post_norm_div_ ;
input p_desc1581_p_O_DFFX1post_norm_div_ ;
input p_desc1582_p_O_DFFX1post_norm_div_ ;
input p_desc1583_p_O_DFFX1post_norm_div_ ;
input p_desc1584_p_O_DFFX1post_norm_div_ ;
input p_desc1585_p_O_DFFX1post_norm_div_ ;
input p_desc1586_p_O_DFFX1post_norm_div_ ;
input p_desc1587_p_O_DFFX1post_norm_div_ ;
input p_desc1588_p_O_DFFX1post_norm_div_ ;
input p_desc1589_p_O_DFFX1post_norm_div_ ;
input p_desc1590_p_O_DFFX1post_norm_div_ ;
input p_desc1591_p_O_DFFX1post_norm_div_ ;
input p_desc1592_p_O_DFFX1post_norm_div_ ;
input p_desc1593_p_O_DFFX1post_norm_div_ ;
input p_desc1594_p_O_DFFX1post_norm_div_ ;
input p_desc1595_p_O_DFFX1post_norm_div_ ;
input p_desc1596_p_O_DFFX1post_norm_div_ ;
input p_desc1597_p_O_DFFX1post_norm_div_ ;
input p_desc1598_p_O_DFFX1post_norm_div_ ;
input p_desc1599_p_O_DFFX1post_norm_div_ ;
input p_desc1600_p_O_DFFX1post_norm_div_ ;
input p_desc1601_p_O_DFFX1post_norm_div_ ;
input p_desc1602_p_O_DFFX1post_norm_div_ ;
input p_desc1603_p_O_DFFX1post_norm_div_ ;
input p_desc1604_p_O_DFFX1post_norm_div_ ;
input p_desc1605_p_O_DFFX1post_norm_div_ ;
input p_desc1606_p_O_DFFX1post_norm_div_ ;
input p_desc1607_p_O_DFFX1post_norm_div_ ;
input p_desc1608_p_O_DFFX1post_norm_div_ ;
input p_desc1609_p_O_DFFX1post_norm_div_ ;
input p_desc1610_p_O_DFFX1post_norm_div_ ;
input p_desc1611_p_O_DFFX1post_norm_div_ ;
input p_desc1612_p_O_DFFX1post_norm_div_ ;
input p_desc1613_p_O_DFFX1post_norm_div_ ;
input p_desc1614_p_O_DFFX1post_norm_div_ ;
input p_desc1615_p_O_DFFX1post_norm_div_ ;
input p_desc1616_p_O_DFFX1post_norm_div_ ;
input p_desc1617_p_O_DFFX1post_norm_div_ ;
input p_desc1618_p_O_DFFX1post_norm_div_ ;
input p_desc1619_p_O_DFFX1post_norm_div_ ;
input p_desc1620_p_O_DFFX1post_norm_div_ ;
input p_desc1621_p_O_DFFX1post_norm_div_ ;
input p_desc1622_p_O_DFFX1post_norm_div_ ;
input p_desc1623_p_O_DFFX1post_norm_div_ ;
input p_desc1624_p_O_DFFX1post_norm_div_ ;
input p_desc1625_p_O_DFFX1post_norm_div_ ;
input p_desc1626_p_O_DFFX1post_norm_div_ ;
input p_desc1627_p_O_DFFX1post_norm_div_ ;
input p_desc1628_p_O_DFFX1post_norm_div_ ;
input p_desc1629_p_O_DFFX1post_norm_div_ ;
input p_desc1630_p_O_DFFX1post_norm_div_ ;
input p_desc1631_p_O_DFFX1post_norm_div_ ;
input p_desc1632_p_O_DFFX1post_norm_div_ ;
input p_desc1633_p_O_DFFX1post_norm_div_ ;
input p_desc1634_p_O_DFFX1post_norm_div_ ;
input p_desc1635_p_O_DFFX1post_norm_div_ ;
input p_desc1636_p_O_DFFX1post_norm_div_ ;
input p_desc1637_p_O_DFFX1post_norm_div_ ;
input p_desc1638_p_O_DFFX1post_norm_div_ ;
input p_desc1639_p_O_DFFX1post_norm_div_ ;
input p_desc1640_p_O_DFFX1post_norm_div_ ;
input p_desc1641_p_O_DFFX1post_norm_div_ ;
input p_desc1642_p_O_DFFX1post_norm_div_ ;
input p_desc1643_p_O_DFFX1post_norm_div_ ;
input p_desc1644_p_O_DFFX1post_norm_div_ ;
input p_desc1645_p_O_DFFX1post_norm_div_ ;
input p_desc1646_p_O_DFFX1post_norm_div_ ;
input p_desc1647_p_O_DFFX1post_norm_div_ ;
input p_desc1648_p_O_DFFX1post_norm_div_ ;
input p_desc1649_p_O_DFFX1post_norm_div_ ;
input p_desc1650_p_O_DFFX1post_norm_div_ ;
input p_desc1651_p_O_DFFX1post_norm_div_ ;
input p_s_sign_i_reg_p_O_DFFX1post_norm_div_ ;
input p_desc1652_p_O_DFFX1post_norm_div_ ;
input p_desc1653_p_O_DFFX1post_norm_div_ ;
input p_desc1654_p_O_DFFX1post_norm_div_ ;
input p_desc1658_p_O_DFFX1post_norm_div_ ;
input p_desc1659_p_O_DFFX1post_norm_div_ ;
input p_desc1663_p_O_DFFX1post_norm_div_ ;
input p_desc1664_p_O_DFFX1post_norm_div_ ;
input p_desc1665_p_O_DFFX1post_norm_div_ ;
input p_desc1666_p_O_DFFX1post_norm_div_ ;
input p_desc1667_p_O_DFFX1post_norm_div_ ;
input p_desc1668_p_O_DFFX1post_norm_div_ ;
input p_desc1669_p_O_DFFX1post_norm_div_ ;
input p_desc1670_p_O_DFFX1post_norm_div_ ;
input p_desc1671_p_O_DFFX1post_norm_div_ ;
input p_desc1672_p_O_DFFX1post_norm_div_ ;
input p_desc1673_p_O_DFFX1post_norm_div_ ;
input p_desc1674_p_O_DFFX1post_norm_div_ ;
input p_desc1675_p_O_DFFX1post_norm_div_ ;
input p_desc1676_p_O_DFFX1post_norm_div_ ;
input p_desc1677_p_O_DFFX1post_norm_div_ ;
input p_desc1678_p_O_DFFX1post_norm_div_ ;
input p_desc1679_p_O_DFFX1post_norm_div_ ;
input p_desc1680_p_O_DFFX1post_norm_div_ ;
input p_desc1681_p_O_DFFX1post_norm_div_ ;
input p_desc1682_p_O_DFFX1post_norm_div_ ;
input p_desc1683_p_O_DFFX1post_norm_div_ ;
input p_desc1684_p_O_DFFX1post_norm_div_ ;
input p_desc1685_p_O_DFFX1post_norm_div_ ;
input p_desc1686_p_O_DFFX1post_norm_div_ ;
input p_desc1687_p_O_DFFX1post_norm_div_ ;
input p_desc1688_p_O_DFFX1post_norm_div_ ;
input p_desc1689_p_O_DFFX1post_norm_div_ ;
input p_desc1690_p_O_DFFX1post_norm_div_ ;
input p_desc1691_p_O_DFFX1post_norm_div_ ;
input p_desc1692_p_O_DFFX1post_norm_div_ ;
input p_desc1693_p_O_DFFX1post_norm_div_ ;
input p_desc1694_p_O_DFFX1post_norm_div_ ;
input p_desc1695_p_O_DFFX1post_norm_div_ ;
input p_desc1696_p_O_DFFX1post_norm_div_ ;
input p_desc1697_p_O_DFFX1post_norm_div_ ;
input p_desc1698_p_O_DFFX1post_norm_div_ ;
input p_desc1699_p_O_DFFX1post_norm_div_ ;
input p_desc1700_p_O_DFFX1post_norm_div_ ;
input p_desc1701_p_O_DFFX1post_norm_div_ ;
input p_desc1702_p_O_DFFX1post_norm_div_ ;
input p_desc1703_p_O_DFFX1post_norm_div_ ;
input p_desc1704_p_O_DFFX1post_norm_div_ ;
input p_desc1705_p_O_DFFX1post_norm_div_ ;
input p_desc1706_p_O_DFFX1post_norm_div_ ;
input p_desc1707_p_O_DFFX1post_norm_div_ ;
input p_desc1708_p_O_DFFX1post_norm_div_ ;
input p_desc1709_p_O_DFFX1post_norm_div_ ;
input p_desc1710_p_O_DFFX1post_norm_div_ ;
input p_desc1711_p_O_DFFX1post_norm_div_ ;
input p_desc1712_p_O_DFFX1post_norm_div_ ;
input p_desc1713_p_O_DFFX1post_norm_div_ ;
input p_desc1714_p_O_DFFX1post_norm_div_ ;
input p_desc1715_p_O_DFFX1post_norm_div_ ;
input p_desc1716_p_O_DFFX1post_norm_div_ ;
input p_desc1717_p_O_DFFX1post_norm_div_ ;
input p_desc1718_p_O_DFFX1post_norm_div_ ;
input p_desc1719_p_O_DFFX1post_norm_div_ ;
input p_desc1720_p_O_DFFX1post_norm_div_ ;
input p_desc1721_p_O_DFFX1post_norm_div_ ;
input p_desc1722_p_O_DFFX1post_norm_div_ ;
input p_desc1723_p_O_DFFX1post_norm_div_ ;
input p_desc1724_p_O_DFFX1post_norm_div_ ;
input p_desc1725_p_O_DFFX1post_norm_div_ ;
input p_desc1726_p_O_DFFX1post_norm_div_ ;
input p_desc1727_p_O_DFFX1post_norm_div_ ;
input p_desc1728_p_O_DFFX1post_norm_div_ ;
input p_ine_o_reg_p_O_DFFX1post_norm_div_ ;
input p_desc1729_p_O_DFFX1post_norm_div_ ;
input p_desc1737_p_O_DFFX1post_norm_div_ ;
input p_desc1738_p_O_DFFX1post_norm_div_ ;
input p_desc1739_p_O_DFFX1post_norm_div_ ;
input p_desc1740_p_O_DFFX1post_norm_div_ ;
input p_desc1741_p_O_DFFX1post_norm_div_ ;
input p_desc1742_p_O_DFFX1post_norm_div_ ;
input p_desc1743_p_O_DFFX1post_norm_div_ ;
input p_desc1744_p_O_DFFX1post_norm_div_ ;
input p_desc1745_p_O_DFFX1post_norm_div_ ;
input p_desc1746_p_O_DFFX1post_norm_div_ ;
input p_desc1747_p_O_DFFX1post_norm_div_ ;
input p_desc1748_p_O_DFFX1post_norm_div_ ;
input p_desc1749_p_O_DFFX1post_norm_div_ ;
input p_desc1750_p_O_DFFX1post_norm_div_ ;
input p_desc1751_p_O_DFFX1post_norm_div_ ;
input p_desc1752_p_O_DFFX1post_norm_div_ ;
input p_desc1753_p_O_DFFX1post_norm_div_ ;
input p_desc1754_p_O_DFFX1post_norm_div_ ;
input p_desc1755_p_O_DFFX1post_norm_div_ ;
input p_desc1756_p_O_DFFX1post_norm_div_ ;
input p_desc1757_p_O_DFFX1post_norm_div_ ;
input p_desc1758_p_O_DFFX1post_norm_div_ ;
input p_desc1849_p_O_DFFX1post_norm_div_ ;
input p_desc1850_p_O_DFFX1post_norm_div_ ;
input p_desc1851_p_O_DFFX1post_norm_div_ ;
input p_desc1852_p_O_DFFX1post_norm_div_ ;
input p_desc1853_p_O_DFFX1post_norm_div_ ;
input p_desc1854_p_O_DFFX1post_norm_div_ ;
input p_desc1855_p_O_DFFX1post_norm_div_ ;
input p_desc1856_p_O_DFFX1post_norm_div_ ;
input p_desc1857_p_O_DFFX1post_norm_div_ ;
input p_desc1858_p_O_DFFX1post_norm_div_ ;
input p_desc1859_p_O_DFFX1post_norm_div_ ;
input p_desc1860_p_O_DFFX1post_norm_div_ ;
input p_desc1861_p_O_DFFX1post_norm_div_ ;
input p_desc1862_p_O_DFFX1post_norm_div_ ;
input p_desc1863_p_O_DFFX1post_norm_div_ ;
input p_desc1864_p_O_DFFX1post_norm_div_ ;
input p_desc1865_p_O_DFFX1post_norm_div_ ;
input p_desc1866_p_O_DFFX1post_norm_div_ ;
input p_desc1867_p_O_DFFX1post_norm_div_ ;
input p_desc1868_p_O_DFFX1post_norm_div_ ;
input p_desc1869_p_O_DFFX1post_norm_div_ ;
// instances
  DFFX1 desc2406(.D(opa_i[31:31]),.CLK(clk_i),.Q(s_opa_i[31:31]));
  DFFX1 desc2407(.D(opa_i[30:30]),.CLK(clk_i),.Q(s_opa_i[30:30]));
  DFFX1 desc2408(.D(opa_i[29:29]),.CLK(clk_i),.Q(s_opa_i[29:29]));
  DFFX1 desc2409(.D(opa_i[28:28]),.CLK(clk_i),.Q(s_opa_i[28:28]),.QN(n154));
  DFFX1 desc2410(.D(opa_i[27:27]),.CLK(clk_i),.Q(s_opa_i[27:27]),.QN(n153));
  DFFX1 desc2411(.D(opa_i[26:26]),.CLK(clk_i),.Q(s_opa_i[26:26]),.QN(n152));
  DFFX1 desc2412(.D(opa_i[25:25]),.CLK(clk_i),.Q(s_opa_i[25:25]),.QN(n151));
  DFFX1 desc2413(.D(opa_i[24:24]),.CLK(clk_i),.Q(s_opa_i[24:24]),.QN(n162));
  DFFX1 desc2414(.D(opa_i[23:23]),.CLK(clk_i),.Q(s_opa_i[23:23]),.QN(n161));
  DFFX1 desc2415(.D(opa_i[22:22]),.CLK(clk_i),.Q(s_opa_i[22:22]),.QN(n144));
  DFFX1 desc2416(.D(opa_i[21:21]),.CLK(clk_i),.Q(s_opa_i[21:21]));
  DFFX1 desc2417(.D(opa_i[20:20]),.CLK(clk_i),.Q(s_opa_i[20:20]));
  DFFX1 desc2418(.D(opa_i[19:19]),.CLK(clk_i),.Q(s_opa_i[19:19]),.QN(n143));
  DFFX1 desc2419(.D(opa_i[18:18]),.CLK(clk_i),.Q(s_opa_i[18:18]),.QN(n142));
  DFFX1 desc2420(.D(opa_i[17:17]),.CLK(clk_i),.Q(s_opa_i[17:17]),.QN(n141));
  DFFX1 desc2421(.D(opa_i[16:16]),.CLK(clk_i),.Q(s_opa_i[16:16]));
  DFFX1 desc2422(.D(opa_i[15:15]),.CLK(clk_i),.Q(s_opa_i[15:15]));
  DFFX1 desc2423(.D(opa_i[14:14]),.CLK(clk_i),.Q(s_opa_i[14:14]));
  DFFX1 desc2424(.D(opa_i[13:13]),.CLK(clk_i),.Q(s_opa_i[13:13]));
  DFFX1 desc2425(.D(opa_i[12:12]),.CLK(clk_i),.Q(s_opa_i[12:12]));
  DFFX1 desc2426(.D(opa_i[11:11]),.CLK(clk_i),.Q(s_opa_i[11:11]));
  DFFX1 desc2427(.D(opa_i[10:10]),.CLK(clk_i),.Q(s_opa_i[10:10]),.QN(n150));
  DFFX1 desc2428(.D(opa_i[9:9]),.CLK(clk_i),.Q(s_opa_i[9:9]),.QN(n149));
  DFFX1 desc2429(.D(opa_i[8:8]),.CLK(clk_i),.Q(s_opa_i[8:8]),.QN(n148));
  DFFX1 desc2430(.D(opa_i[7:7]),.CLK(clk_i),.Q(s_opa_i[7:7]),.QN(n147));
  DFFX1 desc2431(.D(opa_i[6:6]),.CLK(clk_i),.Q(s_opa_i[6:6]));
  DFFX1 desc2432(.D(opa_i[5:5]),.CLK(clk_i),.Q(s_opa_i[5:5]));
  DFFX1 desc2433(.D(opa_i[4:4]),.CLK(clk_i),.Q(s_opa_i[4:4]));
  DFFX1 desc2434(.D(opa_i[3:3]),.CLK(clk_i),.Q(s_opa_i[3:3]),.QN(n146));
  DFFX1 desc2435(.D(opa_i[2:2]),.CLK(clk_i),.Q(s_opa_i[2:2]),.QN(n145));
  DFFX1 desc2436(.D(opa_i[1:1]),.CLK(clk_i),.Q(s_opa_i[1:1]));
  DFFX1 desc2437(.D(opa_i[0:0]),.CLK(clk_i),.Q(s_opa_i[0:0]));
  DFFX1 desc2438(.D(opb_i[31:31]),.CLK(clk_i),.Q(s_opb_i[31:31]));
  DFFX1 desc2439(.D(opb_i[30:30]),.CLK(clk_i),.Q(s_opb_i[30:30]));
  DFFX1 desc2440(.D(opb_i[29:29]),.CLK(clk_i),.Q(s_opb_i[29:29]));
  DFFX1 desc2441(.D(opb_i[28:28]),.CLK(clk_i),.Q(s_opb_i[28:28]),.QN(n158));
  DFFX1 desc2442(.D(opb_i[27:27]),.CLK(clk_i),.Q(s_opb_i[27:27]),.QN(n157));
  DFFX1 desc2443(.D(opb_i[26:26]),.CLK(clk_i),.Q(s_opb_i[26:26]),.QN(n156));
  DFFX1 desc2444(.D(opb_i[25:25]),.CLK(clk_i),.Q(s_opb_i[25:25]),.QN(n155));
  DFFX1 desc2445(.D(opb_i[24:24]),.CLK(clk_i),.Q(s_opb_i[24:24]),.QN(n160));
  DFFX1 desc2446(.D(opb_i[23:23]),.CLK(clk_i),.Q(s_opb_i[23:23]),.QN(n159));
  DFFX1 desc2447(.D(opb_i[22:22]),.CLK(clk_i),.Q(s_opb_i[22:22]),.QN(n134));
  DFFX1 desc2448(.D(opb_i[21:21]),.CLK(clk_i),.Q(s_opb_i[21:21]));
  DFFX1 desc2449(.D(opb_i[20:20]),.CLK(clk_i),.Q(s_opb_i[20:20]));
  DFFX1 desc2450(.D(opb_i[19:19]),.CLK(clk_i),.Q(s_opb_i[19:19]),.QN(n133));
  DFFX1 desc2451(.D(opb_i[18:18]),.CLK(clk_i),.Q(s_opb_i[18:18]),.QN(n132));
  DFFX1 desc2452(.D(opb_i[17:17]),.CLK(clk_i),.Q(s_opb_i[17:17]),.QN(n131));
  DFFX1 desc2453(.D(opb_i[16:16]),.CLK(clk_i),.Q(s_opb_i[16:16]));
  DFFX1 desc2454(.D(opb_i[15:15]),.CLK(clk_i),.Q(s_opb_i[15:15]));
  DFFX1 desc2455(.D(opb_i[14:14]),.CLK(clk_i),.Q(s_opb_i[14:14]));
  DFFX1 desc2456(.D(opb_i[13:13]),.CLK(clk_i),.Q(s_opb_i[13:13]));
  DFFX1 desc2457(.D(opb_i[12:12]),.CLK(clk_i),.Q(s_opb_i[12:12]));
  DFFX1 desc2458(.D(opb_i[11:11]),.CLK(clk_i),.Q(s_opb_i[11:11]));
  DFFX1 desc2459(.D(opb_i[10:10]),.CLK(clk_i),.Q(s_opb_i[10:10]),.QN(n140));
  DFFX1 desc2460(.D(opb_i[9:9]),.CLK(clk_i),.Q(s_opb_i[9:9]),.QN(n139));
  DFFX1 desc2461(.D(opb_i[8:8]),.CLK(clk_i),.Q(s_opb_i[8:8]),.QN(n138));
  DFFX1 desc2462(.D(opb_i[7:7]),.CLK(clk_i),.Q(s_opb_i[7:7]),.QN(n137));
  DFFX1 desc2463(.D(opb_i[6:6]),.CLK(clk_i),.Q(s_opb_i[6:6]));
  DFFX1 desc2464(.D(opb_i[5:5]),.CLK(clk_i),.Q(s_opb_i[5:5]));
  DFFX1 desc2465(.D(opb_i[4:4]),.CLK(clk_i),.Q(s_opb_i[4:4]));
  DFFX1 desc2466(.D(opb_i[3:3]),.CLK(clk_i),.Q(s_opb_i[3:3]),.QN(n136));
  DFFX1 desc2467(.D(opb_i[2:2]),.CLK(clk_i),.Q(s_opb_i[2:2]),.QN(n135));
  DFFX1 desc2468(.D(opb_i[1:1]),.CLK(clk_i),.Q(s_opb_i[1:1]));
  DFFX1 desc2469(.D(opb_i[0:0]),.CLK(clk_i),.Q(s_opb_i[0:0]));
  DFFX1 desc2470(.D(fpu_op_i[2:2]),.CLK(clk_i),.Q(s_fpu_op_i[2:2]));
  DFFX1 desc2471(.D(fpu_op_i[1:1]),.CLK(clk_i),.Q(s_fpu_op_i[1:1]));
  DFFX1 desc2472(.D(fpu_op_i[0:0]),.CLK(clk_i),.Q(s_fpu_op_i[0:0]));
  DFFX1 desc2473(.D(rmode_i[1:1]),.CLK(clk_i),.Q(s_rmode_i[1:1]),.QN(n215));
  DFFX1 desc2474(.D(rmode_i[0:0]),.CLK(clk_i),.Q(s_rmode_i[0:0]));
  DFFX1 s_start_i_reg(.D(start_i),.CLK(clk_i),.Q(s_start_i),.QN(n218));
  DFFX1 div_zero_o_reg(.D(n197),.CLK(clk_i),.Q(div_zero_o));
  DFFX1 snan_o_reg(.D(N581),.CLK(clk_i),.Q(snan_o));
  DFFX1 s_ine_o_reg(.D(N374),.CLK(clk_i),.Q(s_ine_o),.QN(n217));
  DFFX1 ine_o_reg(.D(s_ine_o),.CLK(clk_i),.Q(ine_o));
  DFFX1 desc2475(.D(N373),.CLK(clk_i),.Q(s_output1[31:31]),.QN(n219));
  DFFX1 desc2476(.D(N372),.CLK(clk_i),.Q(s_output_o[30:30]),.QN(n224));
  DFFX1 desc2477(.D(s_output_o[30:30]),.CLK(clk_i),.Q(output_o[30:30]));
  DFFX1 desc2478(.D(N371),.CLK(clk_i),.Q(s_output_o[29:29]),.QN(n225));
  DFFX1 desc2479(.D(s_output_o[29:29]),.CLK(clk_i),.Q(output_o[29:29]));
  DFFX1 desc2480(.D(N370),.CLK(clk_i),.Q(s_output_o[28:28]));
  DFFX1 desc2481(.D(s_output_o[28:28]),.CLK(clk_i),.Q(output_o[28:28]));
  DFFX1 desc2482(.D(N369),.CLK(clk_i),.Q(s_output_o[27:27]));
  DFFX1 desc2483(.D(s_output_o[27:27]),.CLK(clk_i),.Q(output_o[27:27]));
  DFFX1 desc2484(.D(N368),.CLK(clk_i),.Q(s_output_o[26:26]));
  DFFX1 desc2485(.D(s_output_o[26:26]),.CLK(clk_i),.Q(output_o[26:26]));
  DFFX1 desc2486(.D(N367),.CLK(clk_i),.Q(s_output_o[25:25]));
  DFFX1 desc2487(.D(s_output_o[25:25]),.CLK(clk_i),.Q(output_o[25:25]));
  DFFX1 desc2488(.D(N366),.CLK(clk_i),.Q(s_output_o[24:24]),.QN(n216));
  DFFX1 desc2489(.D(s_output_o[24:24]),.CLK(clk_i),.Q(output_o[24:24]));
  DFFX1 desc2490(.D(N365),.CLK(clk_i),.Q(s_output1[23:23]),.QN(n207));
  DFFX1 underflow_o_reg(.D(N546),.CLK(clk_i),.Q(underflow_o));
  DFFX1 overflow_o_reg(.D(N547),.CLK(clk_i),.Q(overflow_o));
  DFFX1 desc2491(.D(N364),.CLK(clk_i),.Q(s_output1[22:22]),.QN(n214));
  DFFX1 desc2492(.D(N363),.CLK(clk_i),.Q(s_output1[21:21]));
  DFFX1 desc2493(.D(N362),.CLK(clk_i),.QN(n203));
  DFFX1 desc2494(.D(N361),.CLK(clk_i),.QN(n204));
  DFFX1 desc2495(.D(N360),.CLK(clk_i),.QN(n211));
  DFFX1 desc2496(.D(N359),.CLK(clk_i),.QN(n200));
  DFFX1 desc2497(.D(N358),.CLK(clk_i),.Q(s_output1[16:16]));
  DFFX1 desc2498(.D(N357),.CLK(clk_i),.Q(s_output1[15:15]));
  DFFX1 desc2499(.D(N356),.CLK(clk_i),.Q(s_output1[14:14]));
  DFFX1 desc2500(.D(N355),.CLK(clk_i),.Q(s_output1[13:13]));
  DFFX1 desc2501(.D(N354),.CLK(clk_i),.Q(s_output1[12:12]));
  DFFX1 desc2502(.D(N353),.CLK(clk_i),.Q(s_output1[11:11]));
  DFFX1 desc2503(.D(N352),.CLK(clk_i),.QN(n202));
  DFFX1 desc2504(.D(N351),.CLK(clk_i),.QN(n205));
  DFFX1 desc2505(.D(N350),.CLK(clk_i),.QN(n212));
  DFFX1 desc2506(.D(N349),.CLK(clk_i),.QN(n201));
  DFFX1 desc2507(.D(N348),.CLK(clk_i),.Q(s_output1[6:6]));
  DFFX1 desc2508(.D(N347),.CLK(clk_i),.Q(s_output1[5:5]));
  DFFX1 desc2509(.D(N346),.CLK(clk_i),.Q(s_output1[4:4]));
  DFFX1 desc2510(.D(N345),.CLK(clk_i),.Q(s_output1[3:3]));
  DFFX1 desc2511(.D(N344),.CLK(clk_i),.Q(s_output1[2:2]));
  DFFX1 desc2512(.D(N343),.CLK(clk_i),.QN(n210));
  DFFX1 desc2513(.D(N342),.CLK(clk_i),.QN(n209));
  DFFX1 zero_o_reg(.D(n199),.CLK(clk_i),.Q(zero_o));
  DFFX1 desc2514(.D(s_output_o[31:31]),.CLK(clk_i),.Q(output_o[31:31]));
  DFFX1 desc2515(.D(s_output_o[23:23]),.CLK(clk_i),.Q(output_o[23:23]));
  DFFX1 desc2516(.D(s_output_o[11:11]),.CLK(clk_i),.Q(output_o[11:11]));
  DFFX1 desc2517(.D(s_output_o[12:12]),.CLK(clk_i),.Q(output_o[12:12]));
  DFFX1 desc2518(.D(s_output_o[13:13]),.CLK(clk_i),.Q(output_o[13:13]));
  DFFX1 desc2519(.D(s_output_o[14:14]),.CLK(clk_i),.Q(output_o[14:14]));
  DFFX1 desc2520(.D(s_output_o[15:15]),.CLK(clk_i),.Q(output_o[15:15]));
  DFFX1 desc2521(.D(s_output_o[16:16]),.CLK(clk_i),.Q(output_o[16:16]));
  DFFX1 desc2522(.D(s_output_o[21:21]),.CLK(clk_i),.Q(output_o[21:21]));
  DFFX1 desc2523(.D(s_output_o[2:2]),.CLK(clk_i),.Q(output_o[2:2]));
  DFFX1 desc2524(.D(s_output_o[3:3]),.CLK(clk_i),.Q(output_o[3:3]));
  DFFX1 desc2525(.D(s_output_o[4:4]),.CLK(clk_i),.Q(output_o[4:4]));
  DFFX1 desc2526(.D(s_output_o[5:5]),.CLK(clk_i),.Q(output_o[5:5]));
  DFFX1 desc2527(.D(s_output_o[6:6]),.CLK(clk_i),.Q(output_o[6:6]));
  DFFX1 desc2528(.D(s_output_o[9:9]),.CLK(clk_i),.Q(output_o[9:9]));
  DFFX1 desc2529(.D(s_output_o[8:8]),.CLK(clk_i),.Q(output_o[8:8]));
  DFFX1 desc2530(.D(s_output_o[7:7]),.CLK(clk_i),.Q(output_o[7:7]));
  DFFX1 desc2531(.D(s_output_o[22:22]),.CLK(clk_i),.Q(output_o[22:22]));
  DFFX1 desc2532(.D(s_output_o[20:20]),.CLK(clk_i),.Q(output_o[20:20]));
  DFFX1 desc2533(.D(s_output_o[1:1]),.CLK(clk_i),.Q(output_o[1:1]));
  DFFX1 desc2534(.D(s_output_o[19:19]),.CLK(clk_i),.Q(output_o[19:19]));
  DFFX1 desc2535(.D(s_output_o[18:18]),.CLK(clk_i),.Q(output_o[18:18]));
  DFFX1 desc2536(.D(s_output_o[17:17]),.CLK(clk_i),.Q(output_o[17:17]));
  DFFX1 desc2537(.D(s_output_o[10:10]),.CLK(clk_i),.Q(output_o[10:10]));
  DFFX1 desc2538(.D(s_output_o[0:0]),.CLK(clk_i),.Q(output_o[0:0]));
  DFFX1 inf_o_reg(.D(N549),.CLK(clk_i),.Q(inf_o));
  DFFX1 qnan_o_reg(.D(n198),.CLK(clk_i),.Q(qnan_o));
  DFFX1 desc2539(.D(n196),.CLK(clk_i),.Q(s_count[0:0]));
  DFFX1 ready_o_reg(.D(n195),.CLK(clk_i),.Q(ready_o));
  DFFX1 s_state_reg(.D(n194),.CLK(clk_i),.Q(s_state));
  DFFX1 desc2540(.D(n193),.CLK(clk_i),.Q(s_count[31:31]));
  DFFX1 desc2541(.D(n192),.CLK(clk_i),.Q(s_count[1:1]),.QN(n206));
  DFFX1 desc2542(.D(n191),.CLK(clk_i),.Q(s_count[2:2]),.QN(n208));
  DFFX1 desc2543(.D(n190),.CLK(clk_i),.Q(s_count[3:3]),.QN(n213));
  DFFX1 desc2544(.D(n189),.CLK(clk_i),.Q(s_count[4:4]));
  DFFX1 desc2545(.D(n188),.CLK(clk_i),.Q(s_count[5:5]),.QN(n221));
  DFFX1 desc2546(.D(n187),.CLK(clk_i),.Q(s_count[6:6]));
  DFFX1 desc2547(.D(n186),.CLK(clk_i),.Q(s_count[7:7]));
  DFFX1 desc2548(.D(n185),.CLK(clk_i),.Q(s_count[8:8]));
  DFFX1 desc2549(.D(n184),.CLK(clk_i),.Q(s_count[9:9]));
  DFFX1 desc2550(.D(n183),.CLK(clk_i),.Q(s_count[10:10]));
  DFFX1 desc2551(.D(n182),.CLK(clk_i),.Q(s_count[11:11]));
  DFFX1 desc2552(.D(n181),.CLK(clk_i),.Q(s_count[12:12]));
  DFFX1 desc2553(.D(n180),.CLK(clk_i),.Q(s_count[13:13]));
  DFFX1 desc2554(.D(n179),.CLK(clk_i),.Q(s_count[14:14]));
  DFFX1 desc2555(.D(n178),.CLK(clk_i),.Q(s_count[15:15]));
  DFFX1 desc2556(.D(n177),.CLK(clk_i),.Q(s_count[16:16]));
  DFFX1 desc2557(.D(n176),.CLK(clk_i),.Q(s_count[17:17]));
  DFFX1 desc2558(.D(n175),.CLK(clk_i),.Q(s_count[18:18]));
  DFFX1 desc2559(.D(n174),.CLK(clk_i),.Q(s_count[19:19]));
  DFFX1 desc2560(.D(n173),.CLK(clk_i),.Q(s_count[20:20]));
  DFFX1 desc2561(.D(n172),.CLK(clk_i),.Q(s_count[21:21]));
  DFFX1 desc2562(.D(n171),.CLK(clk_i),.Q(s_count[22:22]));
  DFFX1 desc2563(.D(n170),.CLK(clk_i),.Q(s_count[23:23]));
  DFFX1 desc2564(.D(n169),.CLK(clk_i),.Q(s_count[24:24]));
  DFFX1 desc2565(.D(n168),.CLK(clk_i),.Q(s_count[25:25]));
  DFFX1 desc2566(.D(n167),.CLK(clk_i),.Q(s_count[26:26]));
  DFFX1 desc2567(.D(n166),.CLK(clk_i),.Q(s_count[27:27]));
  DFFX1 desc2568(.D(n165),.CLK(clk_i),.Q(s_count[28:28]));
  DFFX1 desc2569(.D(n164),.CLK(clk_i),.Q(s_count[29:29]));
  DFFX1 desc2570(.D(n163),.CLK(clk_i),.Q(s_count[30:30]));
  AO21X1 U3(.IN1(s_state),.IN2(n1),.IN3(s_start_i),.Q(n194));
  OR2X1 U7(.IN1(s_output1[6:6]),.IN2(n272),.Q(s_output_o[6:6]));
  OR2X1 U8(.IN1(s_output1[5:5]),.IN2(n272),.Q(s_output_o[5:5]));
  OR2X1 U9(.IN1(s_output1[4:4]),.IN2(n272),.Q(s_output_o[4:4]));
  OR2X1 U10(.IN1(s_output1[3:3]),.IN2(n272),.Q(s_output_o[3:3]));
  NOR4X0 U13(.IN1(s_fpu_op_i[2:2]),.IN2(s_fpu_op_i[1:1]),.IN3(n11),.IN4(n215),.QN(n10));
  XOR2X1 U16(.IN1(s_opb_i[31:31]),.IN2(s_fpu_op_i[0:0]),.Q(n13));
  OR2X1 U18(.IN1(s_output1[2:2]),.IN2(n272),.Q(s_output_o[2:2]));
  OR2X1 U21(.IN1(s_output1[21:21]),.IN2(n272),.Q(s_output_o[21:21]));
  OR2X1 U27(.IN1(s_output1[16:16]),.IN2(n272),.Q(s_output_o[16:16]));
  OR2X1 U28(.IN1(s_output1[15:15]),.IN2(n272),.Q(s_output_o[15:15]));
  OR2X1 U29(.IN1(s_output1[14:14]),.IN2(n272),.Q(s_output_o[14:14]));
  OR2X1 U30(.IN1(s_output1[13:13]),.IN2(n272),.Q(s_output_o[13:13]));
  OR2X1 U31(.IN1(s_output1[12:12]),.IN2(n272),.Q(s_output_o[12:12]));
  OR2X1 U32(.IN1(s_output1[11:11]),.IN2(n272),.Q(s_output_o[11:11]));
  NOR4X0 U37(.IN1(n198),.IN2(n25),.IN3(n26),.IN4(n197),.QN(n9));
  XNOR2X1 U38(.IN1(s_rmode_i[0:0]),.IN2(n27),.Q(n24));
  AO22X1 U41(.IN1(s_count[9:9]),.IN2(n250),.IN3(N44),.IN4(n247),.Q(n184));
  AO22X1 U42(.IN1(s_count[8:8]),.IN2(n251),.IN3(N43),.IN4(n247),.Q(n185));
  AO22X1 U43(.IN1(s_count[7:7]),.IN2(n251),.IN3(N42),.IN4(n247),.Q(n186));
  AO22X1 U44(.IN1(s_count[6:6]),.IN2(n251),.IN3(N41),.IN4(n247),.Q(n187));
  AO22X1 U45(.IN1(n250),.IN2(s_count[5:5]),.IN3(N40),.IN4(n247),.Q(n188));
  AO22X1 U46(.IN1(s_count[4:4]),.IN2(n251),.IN3(N39),.IN4(n247),.Q(n189));
  AO22X1 U47(.IN1(n250),.IN2(s_count[3:3]),.IN3(N38),.IN4(n247),.Q(n190));
  AO22X1 U48(.IN1(s_count[31:31]),.IN2(n251),.IN3(N66),.IN4(n247),.Q(n193));
  AO22X1 U49(.IN1(s_count[30:30]),.IN2(n251),.IN3(N65),.IN4(n247),.Q(n163));
  AO22X1 U50(.IN1(n250),.IN2(s_count[2:2]),.IN3(N37),.IN4(n247),.Q(n191));
  AO22X1 U51(.IN1(s_count[29:29]),.IN2(n251),.IN3(N64),.IN4(n247),.Q(n164));
  AO22X1 U52(.IN1(s_count[28:28]),.IN2(n251),.IN3(N63),.IN4(n247),.Q(n165));
  AO22X1 U53(.IN1(s_count[27:27]),.IN2(n251),.IN3(N62),.IN4(n248),.Q(n166));
  AO22X1 U54(.IN1(s_count[26:26]),.IN2(n251),.IN3(N61),.IN4(n248),.Q(n167));
  AO22X1 U55(.IN1(s_count[25:25]),.IN2(n251),.IN3(N60),.IN4(n248),.Q(n168));
  AO22X1 U56(.IN1(s_count[24:24]),.IN2(n251),.IN3(N59),.IN4(n248),.Q(n169));
  AO22X1 U57(.IN1(s_count[23:23]),.IN2(n251),.IN3(N58),.IN4(n248),.Q(n170));
  AO22X1 U58(.IN1(s_count[22:22]),.IN2(n250),.IN3(N57),.IN4(n248),.Q(n171));
  AO22X1 U59(.IN1(s_count[21:21]),.IN2(n250),.IN3(N56),.IN4(n248),.Q(n172));
  AO22X1 U60(.IN1(s_count[20:20]),.IN2(n250),.IN3(N55),.IN4(n248),.Q(n173));
  AO22X1 U61(.IN1(n250),.IN2(s_count[1:1]),.IN3(N36),.IN4(n248),.Q(n192));
  AO22X1 U62(.IN1(s_count[19:19]),.IN2(n250),.IN3(N54),.IN4(n248),.Q(n174));
  AO22X1 U63(.IN1(s_count[18:18]),.IN2(n250),.IN3(N53),.IN4(n248),.Q(n175));
  AO22X1 U64(.IN1(s_count[17:17]),.IN2(n250),.IN3(N52),.IN4(n248),.Q(n176));
  AO22X1 U65(.IN1(s_count[16:16]),.IN2(n250),.IN3(N51),.IN4(n249),.Q(n177));
  AO22X1 U66(.IN1(s_count[15:15]),.IN2(n250),.IN3(N50),.IN4(n249),.Q(n178));
  AO22X1 U67(.IN1(s_count[14:14]),.IN2(n250),.IN3(N49),.IN4(n249),.Q(n179));
  AO22X1 U68(.IN1(s_count[13:13]),.IN2(n250),.IN3(N48),.IN4(n249),.Q(n180));
  AO22X1 U69(.IN1(s_count[12:12]),.IN2(n250),.IN3(N47),.IN4(n249),.Q(n181));
  AO22X1 U70(.IN1(s_count[11:11]),.IN2(n250),.IN3(N46),.IN4(n249),.Q(n182));
  AO22X1 U71(.IN1(s_count[10:10]),.IN2(n250),.IN3(N45),.IN4(n249),.Q(n183));
  AO22X1 U72(.IN1(n250),.IN2(s_count[0:0]),.IN3(N35),.IN4(n249),.Q(n196));
  NOR3X0 U73(.IN1(n250),.IN2(s_start_i),.IN3(n273),.QN(n30));
  NOR3X0 U74(.IN1(s_start_i),.IN2(s_state),.IN3(n273),.QN(n29));
  AO22X1 U75(.IN1(n273),.IN2(n218),.IN3(ready_o),.IN4(n33),.Q(n195));
  OR2X1 U76(.IN1(s_state),.IN2(s_start_i),.Q(n33));
  NAND3X0 U82(.IN1(n244),.IN2(n41),.IN3(s_count[3:3]),.QN(n38));
  NAND4X0 U83(.IN1(s_count[2:2]),.IN2(n241),.IN3(n43),.IN4(n44),.QN(n37));
  OR2X1 U88(.IN1(n239),.IN2(n236),.Q(n45));
  AND3X1 U89(.IN1(n44),.IN2(n208),.IN3(s_count[0:0]),.Q(n41));
  AND4X1 U91(.IN1(n50),.IN2(n51),.IN3(n52),.IN4(n53),.Q(n44));
  NOR4X0 U92(.IN1(n54),.IN2(s_count[30:30]),.IN3(s_count[4:4]),.IN4(s_count[31:31]),.QN(n53));
  OR4X1 U93(.IN1(s_count[6:6]),.IN2(s_count[7:7]),.IN3(s_count[8:8]),.IN4(s_count[9:9]),.Q(n54));
  NOR4X0 U94(.IN1(n55),.IN2(s_count[23:23]),.IN3(s_count[25:25]),.IN4(s_count[24:24]),.QN(n52));
  OR4X1 U95(.IN1(s_count[26:26]),.IN2(s_count[27:27]),.IN3(s_count[28:28]),.IN4(s_count[29:29]),.Q(n55));
  NOR4X0 U96(.IN1(n56),.IN2(s_count[16:16]),.IN3(s_count[18:18]),.IN4(s_count[17:17]),.QN(n51));
  OR4X1 U97(.IN1(s_count[19:19]),.IN2(s_count[20:20]),.IN3(s_count[21:21]),.IN4(s_count[22:22]),.Q(n56));
  NOR4X0 U98(.IN1(n57),.IN2(s_count[10:10]),.IN3(s_count[12:12]),.IN4(s_count[11:11]),.QN(n50));
  OR3X1 U99(.IN1(s_count[14:14]),.IN2(s_count[15:15]),.IN3(s_count[13:13]),.Q(n57));
  AND2X1 U100(.IN1(serial_div_div_zero),.IN2(n239),.Q(n197));
  NOR3X0 U101(.IN1(n58),.IN2(s_output1[22:22]),.IN3(n59),.QN(n199));
  NOR3X0 U102(.IN1(n28),.IN2(N581),.IN3(n198),.QN(N549));
  NOR3X0 U103(.IN1(n58),.IN2(n28),.IN3(n214),.QN(n198));
  NAND4X0 U105(.IN1(n60),.IN2(n61),.IN3(n62),.IN4(n63),.QN(n58));
  NOR4X0 U106(.IN1(n64),.IN2(s_output1[4:4]),.IN3(s_output1[6:6]),.IN4(s_output1[5:5]),.QN(n63));
  NAND3X0 U107(.IN1(n212),.IN2(n205),.IN3(n201),.QN(n64));
  NOR4X0 U111(.IN1(n65),.IN2(s_output1[21:21]),.IN3(s_output1[3:3]),.IN4(s_output1[2:2]),.QN(n62));
  NOR4X0 U115(.IN1(n66),.IN2(s_output1[14:14]),.IN3(s_output1[16:16]),.IN4(s_output1[15:15]),.QN(n61));
  NAND3X0 U116(.IN1(n211),.IN2(n204),.IN3(n200),.QN(n66));
  NOR4X0 U120(.IN1(n67),.IN2(s_output1[11:11]),.IN3(s_output1[13:13]),.IN4(s_output1[12:12]),.QN(n60));
  NAND4X0 U125(.IN1(n70),.IN2(n71),.IN3(n72),.IN4(n73),.QN(n69));
  NOR4X0 U126(.IN1(n74),.IN2(n255),.IN3(n257),.IN4(n256),.QN(n73));
  NAND3X0 U127(.IN1(n148),.IN2(n149),.IN3(n147),.QN(n74));
  NOR4X0 U128(.IN1(n75),.IN2(n252),.IN3(s_opa_i[21:21]),.IN4(n235),.QN(n72));
  NAND3X0 U129(.IN1(n145),.IN2(n146),.IN3(n144),.QN(n75));
  NOR4X0 U130(.IN1(n76),.IN2(n264),.IN3(n266),.IN4(n265),.QN(n71));
  NAND3X0 U131(.IN1(n142),.IN2(n143),.IN3(n141),.QN(n76));
  NOR4X0 U132(.IN1(n77),.IN2(n262),.IN3(n263),.IN4(n232),.QN(n70));
  NAND3X0 U133(.IN1(n25),.IN2(n150),.IN3(s_opa_i[0:0]),.QN(n77));
  AND4X1 U134(.IN1(n229),.IN2(n270),.IN3(n78),.IN4(n79),.Q(n25));
  NOR4X0 U135(.IN1(n161),.IN2(n162),.IN3(n151),.IN4(n152),.QN(n79));
  NAND4X0 U137(.IN1(n80),.IN2(n81),.IN3(n82),.IN4(n83),.QN(n68));
  NOR4X0 U138(.IN1(n84),.IN2(s_opb_i[4:4]),.IN3(s_opb_i[6:6]),.IN4(s_opb_i[5:5]),.QN(n83));
  NAND3X0 U139(.IN1(n138),.IN2(n139),.IN3(n137),.QN(n84));
  NOR4X0 U140(.IN1(n85),.IN2(s_opb_i[1:1]),.IN3(s_opb_i[21:21]),.IN4(s_opb_i[20:20]),.QN(n82));
  NAND3X0 U141(.IN1(n135),.IN2(n136),.IN3(n134),.QN(n85));
  NOR4X0 U142(.IN1(n86),.IN2(s_opb_i[14:14]),.IN3(s_opb_i[16:16]),.IN4(s_opb_i[15:15]),.QN(n81));
  NAND3X0 U143(.IN1(n132),.IN2(n133),.IN3(n131),.QN(n86));
  NOR4X0 U144(.IN1(n87),.IN2(s_opb_i[11:11]),.IN3(s_opb_i[13:13]),.IN4(s_opb_i[12:12]),.QN(n80));
  NAND3X0 U145(.IN1(n26),.IN2(n140),.IN3(s_opb_i[0:0]),.QN(n87));
  AND4X1 U146(.IN1(s_opb_i[30:30]),.IN2(s_opb_i[29:29]),.IN3(n88),.IN4(n89),.Q(n26));
  NOR4X0 U147(.IN1(n159),.IN2(n160),.IN3(n155),.IN4(n156),.QN(n89));
  NAND4X0 U155(.IN1(n207),.IN2(n216),.IN3(n94),.IN4(n95),.QN(n59));
  NOR4X0 U156(.IN1(s_output_o[30:30]),.IN2(s_output_o[29:29]),.IN3(s_output_o[28:28]),.IN4(s_output_o[27:27]),.QN(n95));
  AO221X1 U160(.IN1(postnorm_addsub_ine_o),.IN2(n241),.IN3(post_norm_sqrt_ine_o),.IN4(n236),.IN5(n96),.Q(N374));
  AO22X1 U161(.IN1(post_norm_div_ine),.IN2(n239),.IN3(post_norm_mul_ine),.IN4(n244),.Q(n96));
  AO221X1 U162(.IN1(postnorm_addsub_output_o[31:31]),.IN2(n241),.IN3(post_norm_sqrt_output[31:31]),.IN4(n236),.IN5(n97),.Q(N373));
  AO22X1 U163(.IN1(post_norm_div_output[31:31]),.IN2(n239),.IN3(post_norm_mul_output[31:31]),.IN4(n244),.Q(n97));
  AO221X1 U164(.IN1(postnorm_addsub_output_o[30:30]),.IN2(n241),.IN3(post_norm_sqrt_output[30:30]),.IN4(n236),.IN5(n98),.Q(N372));
  AO22X1 U165(.IN1(post_norm_div_output[30:30]),.IN2(n239),.IN3(post_norm_mul_output[30:30]),.IN4(n244),.Q(n98));
  AO221X1 U166(.IN1(postnorm_addsub_output_o[29:29]),.IN2(n241),.IN3(post_norm_sqrt_output[29:29]),.IN4(n236),.IN5(n99),.Q(N371));
  AO22X1 U167(.IN1(post_norm_div_output[29:29]),.IN2(n239),.IN3(post_norm_mul_output[29:29]),.IN4(n244),.Q(n99));
  AO221X1 U168(.IN1(postnorm_addsub_output_o[28:28]),.IN2(n241),.IN3(post_norm_sqrt_output[28:28]),.IN4(n236),.IN5(n100),.Q(N370));
  AO22X1 U169(.IN1(post_norm_div_output[28:28]),.IN2(n239),.IN3(post_norm_mul_output[28:28]),.IN4(n244),.Q(n100));
  AO221X1 U170(.IN1(postnorm_addsub_output_o[27:27]),.IN2(n241),.IN3(post_norm_sqrt_output[27:27]),.IN4(n236),.IN5(n101),.Q(N369));
  AO22X1 U171(.IN1(post_norm_div_output[27:27]),.IN2(n239),.IN3(post_norm_mul_output[27:27]),.IN4(n244),.Q(n101));
  AO221X1 U172(.IN1(postnorm_addsub_output_o[26:26]),.IN2(n241),.IN3(post_norm_sqrt_output[26:26]),.IN4(n236),.IN5(n102),.Q(N368));
  AO22X1 U173(.IN1(post_norm_div_output[26:26]),.IN2(n239),.IN3(post_norm_mul_output[26:26]),.IN4(n244),.Q(n102));
  AO221X1 U174(.IN1(postnorm_addsub_output_o[25:25]),.IN2(n241),.IN3(post_norm_sqrt_output[25:25]),.IN4(n236),.IN5(n103),.Q(N367));
  AO22X1 U175(.IN1(post_norm_div_output[25:25]),.IN2(n239),.IN3(post_norm_mul_output[25:25]),.IN4(n244),.Q(n103));
  AO221X1 U176(.IN1(postnorm_addsub_output_o[24:24]),.IN2(n241),.IN3(post_norm_sqrt_output[24:24]),.IN4(n236),.IN5(n104),.Q(N366));
  AO22X1 U177(.IN1(post_norm_div_output[24:24]),.IN2(n239),.IN3(post_norm_mul_output[24:24]),.IN4(n244),.Q(n104));
  AO221X1 U178(.IN1(postnorm_addsub_output_o[23:23]),.IN2(n241),.IN3(post_norm_sqrt_output[23:23]),.IN4(n236),.IN5(n105),.Q(N365));
  AO22X1 U179(.IN1(post_norm_div_output[23:23]),.IN2(n239),.IN3(post_norm_mul_output[23:23]),.IN4(n244),.Q(n105));
  AO221X1 U180(.IN1(postnorm_addsub_output_o[22:22]),.IN2(n241),.IN3(post_norm_sqrt_output[22:22]),.IN4(n236),.IN5(n106),.Q(N364));
  AO22X1 U181(.IN1(post_norm_div_output[22:22]),.IN2(n239),.IN3(post_norm_mul_output[22:22]),.IN4(n244),.Q(n106));
  AO221X1 U182(.IN1(postnorm_addsub_output_o[21:21]),.IN2(n241),.IN3(post_norm_sqrt_output[21:21]),.IN4(n236),.IN5(n107),.Q(N363));
  AO22X1 U183(.IN1(post_norm_div_output[21:21]),.IN2(n239),.IN3(post_norm_mul_output[21:21]),.IN4(n244),.Q(n107));
  AO221X1 U184(.IN1(postnorm_addsub_output_o[20:20]),.IN2(n241),.IN3(post_norm_sqrt_output[20:20]),.IN4(n236),.IN5(n108),.Q(N362));
  AO22X1 U185(.IN1(post_norm_div_output[20:20]),.IN2(n239),.IN3(post_norm_mul_output[20:20]),.IN4(n244),.Q(n108));
  AO221X1 U186(.IN1(postnorm_addsub_output_o[19:19]),.IN2(n241),.IN3(post_norm_sqrt_output[19:19]),.IN4(n236),.IN5(n109),.Q(N361));
  AO22X1 U187(.IN1(post_norm_div_output[19:19]),.IN2(n239),.IN3(post_norm_mul_output[19:19]),.IN4(n244),.Q(n109));
  AO221X1 U188(.IN1(postnorm_addsub_output_o[18:18]),.IN2(n241),.IN3(post_norm_sqrt_output[18:18]),.IN4(n237),.IN5(n110),.Q(N360));
  AO22X1 U189(.IN1(post_norm_div_output[18:18]),.IN2(n239),.IN3(post_norm_mul_output[18:18]),.IN4(n244),.Q(n110));
  AO221X1 U190(.IN1(postnorm_addsub_output_o[17:17]),.IN2(n242),.IN3(post_norm_sqrt_output[17:17]),.IN4(n237),.IN5(n111),.Q(N359));
  AO22X1 U191(.IN1(post_norm_div_output[17:17]),.IN2(n239),.IN3(post_norm_mul_output[17:17]),.IN4(n245),.Q(n111));
  AO221X1 U192(.IN1(postnorm_addsub_output_o[16:16]),.IN2(n242),.IN3(post_norm_sqrt_output[16:16]),.IN4(n237),.IN5(n112),.Q(N358));
  AO22X1 U193(.IN1(post_norm_div_output[16:16]),.IN2(n239),.IN3(post_norm_mul_output[16:16]),.IN4(n245),.Q(n112));
  AO221X1 U194(.IN1(postnorm_addsub_output_o[15:15]),.IN2(n242),.IN3(post_norm_sqrt_output[15:15]),.IN4(n237),.IN5(n113),.Q(N357));
  AO22X1 U195(.IN1(post_norm_div_output[15:15]),.IN2(n240),.IN3(post_norm_mul_output[15:15]),.IN4(n245),.Q(n113));
  AO221X1 U196(.IN1(postnorm_addsub_output_o[14:14]),.IN2(n242),.IN3(post_norm_sqrt_output[14:14]),.IN4(n237),.IN5(n114),.Q(N356));
  AO22X1 U197(.IN1(post_norm_div_output[14:14]),.IN2(n240),.IN3(post_norm_mul_output[14:14]),.IN4(n245),.Q(n114));
  AO221X1 U198(.IN1(postnorm_addsub_output_o[13:13]),.IN2(n242),.IN3(post_norm_sqrt_output[13:13]),.IN4(n237),.IN5(n115),.Q(N355));
  AO22X1 U199(.IN1(post_norm_div_output[13:13]),.IN2(n240),.IN3(post_norm_mul_output[13:13]),.IN4(n245),.Q(n115));
  AO221X1 U200(.IN1(postnorm_addsub_output_o[12:12]),.IN2(n242),.IN3(post_norm_sqrt_output[12:12]),.IN4(n237),.IN5(n116),.Q(N354));
  AO22X1 U201(.IN1(post_norm_div_output[12:12]),.IN2(n240),.IN3(post_norm_mul_output[12:12]),.IN4(n245),.Q(n116));
  AO221X1 U202(.IN1(postnorm_addsub_output_o[11:11]),.IN2(n242),.IN3(post_norm_sqrt_output[11:11]),.IN4(n237),.IN5(n117),.Q(N353));
  AO22X1 U203(.IN1(post_norm_div_output[11:11]),.IN2(n240),.IN3(post_norm_mul_output[11:11]),.IN4(n245),.Q(n117));
  AO221X1 U204(.IN1(postnorm_addsub_output_o[10:10]),.IN2(n242),.IN3(post_norm_sqrt_output[10:10]),.IN4(n237),.IN5(n118),.Q(N352));
  AO22X1 U205(.IN1(post_norm_div_output[10:10]),.IN2(n240),.IN3(post_norm_mul_output[10:10]),.IN4(n245),.Q(n118));
  AO221X1 U206(.IN1(postnorm_addsub_output_o[9:9]),.IN2(n242),.IN3(post_norm_sqrt_output[9:9]),.IN4(n237),.IN5(n119),.Q(N351));
  AO22X1 U207(.IN1(post_norm_div_output[9:9]),.IN2(n240),.IN3(post_norm_mul_output[9:9]),.IN4(n245),.Q(n119));
  AO221X1 U208(.IN1(postnorm_addsub_output_o[8:8]),.IN2(n242),.IN3(post_norm_sqrt_output[8:8]),.IN4(n237),.IN5(n120),.Q(N350));
  AO22X1 U209(.IN1(post_norm_div_output[8:8]),.IN2(n240),.IN3(post_norm_mul_output[8:8]),.IN4(n245),.Q(n120));
  AO221X1 U210(.IN1(postnorm_addsub_output_o[7:7]),.IN2(n242),.IN3(post_norm_sqrt_output[7:7]),.IN4(n237),.IN5(n121),.Q(N349));
  AO22X1 U211(.IN1(post_norm_div_output[7:7]),.IN2(n240),.IN3(post_norm_mul_output[7:7]),.IN4(n245),.Q(n121));
  AO221X1 U212(.IN1(postnorm_addsub_output_o[6:6]),.IN2(n242),.IN3(post_norm_sqrt_output[6:6]),.IN4(n237),.IN5(n122),.Q(N348));
  AO22X1 U213(.IN1(post_norm_div_output[6:6]),.IN2(n240),.IN3(post_norm_mul_output[6:6]),.IN4(n245),.Q(n122));
  AO221X1 U214(.IN1(postnorm_addsub_output_o[5:5]),.IN2(n242),.IN3(post_norm_sqrt_output[5:5]),.IN4(n237),.IN5(n123),.Q(N347));
  AO22X1 U215(.IN1(post_norm_div_output[5:5]),.IN2(n240),.IN3(post_norm_mul_output[5:5]),.IN4(n245),.Q(n123));
  AO221X1 U216(.IN1(postnorm_addsub_output_o[4:4]),.IN2(n242),.IN3(post_norm_sqrt_output[4:4]),.IN4(n237),.IN5(n124),.Q(N346));
  AO22X1 U217(.IN1(post_norm_div_output[4:4]),.IN2(n240),.IN3(post_norm_mul_output[4:4]),.IN4(n245),.Q(n124));
  AO221X1 U218(.IN1(postnorm_addsub_output_o[3:3]),.IN2(n242),.IN3(post_norm_sqrt_output[3:3]),.IN4(n237),.IN5(n125),.Q(N345));
  AO22X1 U219(.IN1(post_norm_div_output[3:3]),.IN2(n240),.IN3(post_norm_mul_output[3:3]),.IN4(n245),.Q(n125));
  AO221X1 U220(.IN1(postnorm_addsub_output_o[2:2]),.IN2(n242),.IN3(post_norm_sqrt_output[2:2]),.IN4(n238),.IN5(n126),.Q(N344));
  AO22X1 U221(.IN1(post_norm_div_output[2:2]),.IN2(n240),.IN3(post_norm_mul_output[2:2]),.IN4(n245),.Q(n126));
  AO221X1 U222(.IN1(postnorm_addsub_output_o[1:1]),.IN2(n243),.IN3(post_norm_sqrt_output[1:1]),.IN4(n238),.IN5(n127),.Q(N343));
  AO22X1 U223(.IN1(post_norm_div_output[1:1]),.IN2(n240),.IN3(post_norm_mul_output[1:1]),.IN4(n246),.Q(n127));
  AO221X1 U224(.IN1(postnorm_addsub_output_o[0:0]),.IN2(n243),.IN3(post_norm_sqrt_output[0:0]),.IN4(n238),.IN5(n128),.Q(N342));
  AO22X1 U225(.IN1(post_norm_div_output[0:0]),.IN2(n240),.IN3(post_norm_mul_output[0:0]),.IN4(n246),.Q(n128));
  NOR3X0 U226(.IN1(fpu_op_i[0:0]),.IN2(fpu_op_i[2:2]),.IN3(n275),.QN(n40));
  AND3X1 U228(.IN1(fpu_op_i[1:1]),.IN2(n274),.IN3(fpu_op_i[0:0]),.Q(n47));
  NOR3X0 U229(.IN1(fpu_op_i[0:0]),.IN2(fpu_op_i[1:1]),.IN3(n274),.QN(n48));
  pre_norm_addsub_inj i_prenorm_addsub(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n228,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n235,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n232,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.fracta_28_o({SYNOPSYS_UNCONNECTED__0,prenorm_addsub_fracta_28_o[26:0]}),.fractb_28_o({SYNOPSYS_UNCONNECTED__1,prenorm_addsub_fractb_28_o[26:0]}),.exp_o(prenorm_addsub_exp_o));
  addsub_28_inj i_addsub(.clk_i(clk_i),.fpu_op_i(s_fpu_op_i[0:0]),.fracta_i({1'b0,prenorm_addsub_fracta_28_o[26:0]}),.fractb_i({1'b0,prenorm_addsub_fractb_28_o[26:0]}),.signa_i(s_opa_i[31:31]),.signb_i(s_opb_i[31:31]),.fract_o(addsub_fract_o),.sign_o(addsub_sign_o));
  post_norm_addsub_inj i_postnorm_addsub(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n234,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n231,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.fract_28_i(addsub_fract_o),.exp_i(prenorm_addsub_exp_o),.sign_i(addsub_sign_o),.fpu_op_i(s_fpu_op_i[0:0]),.rmode_i(s_rmode_i),.output_o(postnorm_addsub_output_o),.ine_o(postnorm_addsub_ine_o));
  pre_norm_mul_inj i_pre_norm_mul(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n233,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n230,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.exp_10_o(pre_norm_mul_exp_10),.fracta_24_o(pre_norm_mul_fracta_24),.fractb_24_o(pre_norm_mul_fractb_24));
  mul_24_inj i_mul_24(.clk_i(clk_i),.fracta_i(pre_norm_mul_fracta_24),.fractb_i(pre_norm_mul_fractb_24),.signa_i(s_opa_i[31:31]),.signb_i(s_opb_i[31:31]),.start_i(start_i),.fract_o(mul_24_fract_48),.sign_o(mul_24_sign));
  serial_mul_inj i_serial_mul(.clk_i(clk_i),.fracta_i(pre_norm_mul_fracta_24),.fractb_i(pre_norm_mul_fractb_24),.signa_i(s_opa_i[31:31]),.signb_i(s_opb_i[31:31]),.start_i(s_start_i));
  post_norm_mul_inj i_post_norm_mul(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n235,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n232,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.exp_10_i(pre_norm_mul_exp_10),.fract_48_i(mul_24_fract_48),.sign_i(mul_24_sign),.rmode_i(s_rmode_i),.output_o(post_norm_mul_output),.ine_o(post_norm_mul_ine));
  pre_norm_div_inj i_pre_norm_div(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n234,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n231,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.exp_10_o(pre_norm_div_exp),.dvdnd_50_o({pre_norm_div_dvdnd[49:26],SYNOPSYS_UNCONNECTED__2,SYNOPSYS_UNCONNECTED__3,SYNOPSYS_UNCONNECTED__4,SYNOPSYS_UNCONNECTED__5,SYNOPSYS_UNCONNECTED__6,SYNOPSYS_UNCONNECTED__7,SYNOPSYS_UNCONNECTED__8,SYNOPSYS_UNCONNECTED__9,SYNOPSYS_UNCONNECTED__10,SYNOPSYS_UNCONNECTED__11,SYNOPSYS_UNCONNECTED__12,SYNOPSYS_UNCONNECTED__13,SYNOPSYS_UNCONNECTED__14,SYNOPSYS_UNCONNECTED__15,SYNOPSYS_UNCONNECTED__16,SYNOPSYS_UNCONNECTED__17,SYNOPSYS_UNCONNECTED__18,SYNOPSYS_UNCONNECTED__19,SYNOPSYS_UNCONNECTED__20,SYNOPSYS_UNCONNECTED__21,SYNOPSYS_UNCONNECTED__22,SYNOPSYS_UNCONNECTED__23,SYNOPSYS_UNCONNECTED__24,SYNOPSYS_UNCONNECTED__25,SYNOPSYS_UNCONNECTED__26,SYNOPSYS_UNCONNECTED__27}),.dvsor_27_o({SYNOPSYS_UNCONNECTED__28,SYNOPSYS_UNCONNECTED__29,SYNOPSYS_UNCONNECTED__30,pre_norm_div_dvsor[23:0]}),.p_desc1176_p_O_DFFX1(p_desc1176_p_O_DFFX1pre_norm_div_),.p_desc1177_p_O_DFFX1(p_desc1177_p_O_DFFX1pre_norm_div_),.p_desc1178_p_O_DFFX1(p_desc1178_p_O_DFFX1pre_norm_div_),.p_desc1179_p_O_DFFX1(p_desc1179_p_O_DFFX1pre_norm_div_),.p_desc1180_p_O_DFFX1(p_desc1180_p_O_DFFX1pre_norm_div_),.p_desc1181_p_O_DFFX1(p_desc1181_p_O_DFFX1pre_norm_div_),.p_desc1182_p_O_DFFX1(p_desc1182_p_O_DFFX1pre_norm_div_),.p_desc1183_p_O_DFFX1(p_desc1183_p_O_DFFX1pre_norm_div_),.p_desc1184_p_O_DFFX1(p_desc1184_p_O_DFFX1pre_norm_div_),.p_desc1185_p_O_DFFX1(p_desc1185_p_O_DFFX1pre_norm_div_),.p_desc1186_p_O_DFFX1(p_desc1186_p_O_DFFX1pre_norm_div_),.p_desc1187_p_O_DFFX1(p_desc1187_p_O_DFFX1pre_norm_div_),.p_desc1188_p_O_DFFX1(p_desc1188_p_O_DFFX1pre_norm_div_),.p_desc1189_p_O_DFFX1(p_desc1189_p_O_DFFX1pre_norm_div_),.p_desc1190_p_O_DFFX1(p_desc1190_p_O_DFFX1pre_norm_div_),.p_desc1191_p_O_DFFX1(p_desc1191_p_O_DFFX1pre_norm_div_),.p_desc1192_p_O_DFFX1(p_desc1192_p_O_DFFX1pre_norm_div_),.p_desc1193_p_O_DFFX1(p_desc1193_p_O_DFFX1pre_norm_div_),.p_desc1194_p_O_DFFX1(p_desc1194_p_O_DFFX1pre_norm_div_),.p_desc1195_p_O_DFFX1(p_desc1195_p_O_DFFX1pre_norm_div_),.p_desc1196_p_O_DFFX1(p_desc1196_p_O_DFFX1pre_norm_div_),.p_desc1197_p_O_DFFX1(p_desc1197_p_O_DFFX1pre_norm_div_),.p_desc1198_p_O_DFFX1(p_desc1198_p_O_DFFX1pre_norm_div_),.p_desc1199_p_O_DFFX1(p_desc1199_p_O_DFFX1pre_norm_div_),.p_desc1200_p_O_DFFX1(p_desc1200_p_O_DFFX1pre_norm_div_),.p_desc1201_p_O_DFFX1(p_desc1201_p_O_DFFX1pre_norm_div_),.p_desc1202_p_O_DFFX1(p_desc1202_p_O_DFFX1pre_norm_div_),.p_desc1203_p_O_DFFX1(p_desc1203_p_O_DFFX1pre_norm_div_),.p_desc1204_p_O_DFFX1(p_desc1204_p_O_DFFX1pre_norm_div_),.p_desc1205_p_O_DFFX1(p_desc1205_p_O_DFFX1pre_norm_div_),.p_desc1206_p_O_DFFX1(p_desc1206_p_O_DFFX1pre_norm_div_),.p_desc1207_p_O_DFFX1(p_desc1207_p_O_DFFX1pre_norm_div_),.p_desc1208_p_O_DFFX1(p_desc1208_p_O_DFFX1pre_norm_div_),.p_desc1209_p_O_DFFX1(p_desc1209_p_O_DFFX1pre_norm_div_),.p_desc1210_p_O_DFFX1(p_desc1210_p_O_DFFX1pre_norm_div_),.p_desc1211_p_O_DFFX1(p_desc1211_p_O_DFFX1pre_norm_div_),.p_desc1212_p_O_DFFX1(p_desc1212_p_O_DFFX1pre_norm_div_),.p_desc1213_p_O_DFFX1(p_desc1213_p_O_DFFX1pre_norm_div_));
  serial_div_inj i_serial_div(.clk_i(clk_i),.dvdnd_i({pre_norm_div_dvdnd[49:26],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.dvsor_i({1'b0,1'b0,1'b0,pre_norm_div_dvsor[23:0]}),.sign_dvd_i(s_opa_i[31:31]),.sign_div_i(s_opb_i[31:31]),.start_i(s_start_i),.qutnt_o(serial_div_qutnt),.rmndr_o(serial_div_rmndr),.sign_o(serial_div_sign),.div_zero_o(serial_div_div_zero),.p_desc1368_p_O_DFFX1(p_desc1368_p_O_DFFX1serial_div_),.p_desc1369_p_O_DFFX1(p_desc1369_p_O_DFFX1serial_div_),.p_desc1370_p_O_DFFX1(p_desc1370_p_O_DFFX1serial_div_),.p_desc1371_p_O_DFFX1(p_desc1371_p_O_DFFX1serial_div_),.p_desc1372_p_O_DFFX1(p_desc1372_p_O_DFFX1serial_div_),.p_desc1373_p_O_DFFX1(p_desc1373_p_O_DFFX1serial_div_),.p_desc1374_p_O_DFFX1(p_desc1374_p_O_DFFX1serial_div_),.p_desc1375_p_O_DFFX1(p_desc1375_p_O_DFFX1serial_div_),.p_desc1376_p_O_DFFX1(p_desc1376_p_O_DFFX1serial_div_),.p_desc1377_p_O_DFFX1(p_desc1377_p_O_DFFX1serial_div_),.p_desc1378_p_O_DFFX1(p_desc1378_p_O_DFFX1serial_div_),.p_desc1379_p_O_DFFX1(p_desc1379_p_O_DFFX1serial_div_),.p_desc1380_p_O_DFFX1(p_desc1380_p_O_DFFX1serial_div_),.p_desc1381_p_O_DFFX1(p_desc1381_p_O_DFFX1serial_div_),.p_desc1382_p_O_DFFX1(p_desc1382_p_O_DFFX1serial_div_),.p_desc1383_p_O_DFFX1(p_desc1383_p_O_DFFX1serial_div_),.p_desc1384_p_O_DFFX1(p_desc1384_p_O_DFFX1serial_div_),.p_desc1385_p_O_DFFX1(p_desc1385_p_O_DFFX1serial_div_),.p_desc1386_p_O_DFFX1(p_desc1386_p_O_DFFX1serial_div_),.p_desc1387_p_O_DFFX1(p_desc1387_p_O_DFFX1serial_div_),.p_desc1388_p_O_DFFX1(p_desc1388_p_O_DFFX1serial_div_),.p_desc1389_p_O_DFFX1(p_desc1389_p_O_DFFX1serial_div_),.p_desc1390_p_O_DFFX1(p_desc1390_p_O_DFFX1serial_div_),.p_desc1391_p_O_DFFX1(p_desc1391_p_O_DFFX1serial_div_),.p_desc1392_p_O_DFFX1(p_desc1392_p_O_DFFX1serial_div_),.p_desc1393_p_O_DFFX1(p_desc1393_p_O_DFFX1serial_div_),.p_desc1394_p_O_DFFX1(p_desc1394_p_O_DFFX1serial_div_),.p_desc1395_p_O_DFFX1(p_desc1395_p_O_DFFX1serial_div_),.p_desc1396_p_O_DFFX1(p_desc1396_p_O_DFFX1serial_div_),.p_desc1397_p_O_DFFX1(p_desc1397_p_O_DFFX1serial_div_),.p_desc1398_p_O_DFFX1(p_desc1398_p_O_DFFX1serial_div_),.p_desc1399_p_O_DFFX1(p_desc1399_p_O_DFFX1serial_div_),.p_desc1400_p_O_DFFX1(p_desc1400_p_O_DFFX1serial_div_),.p_desc1401_p_O_DFFX1(p_desc1401_p_O_DFFX1serial_div_),.p_desc1402_p_O_DFFX1(p_desc1402_p_O_DFFX1serial_div_),.p_desc1403_p_O_DFFX1(p_desc1403_p_O_DFFX1serial_div_),.p_desc1404_p_O_DFFX1(p_desc1404_p_O_DFFX1serial_div_),.p_desc1405_p_O_DFFX1(p_desc1405_p_O_DFFX1serial_div_),.p_desc1406_p_O_DFFX1(p_desc1406_p_O_DFFX1serial_div_),.p_desc1407_p_O_DFFX1(p_desc1407_p_O_DFFX1serial_div_),.p_desc1408_p_O_DFFX1(p_desc1408_p_O_DFFX1serial_div_),.p_desc1409_p_O_DFFX1(p_desc1409_p_O_DFFX1serial_div_),.p_desc1410_p_O_DFFX1(p_desc1410_p_O_DFFX1serial_div_),.p_desc1411_p_O_DFFX1(p_desc1411_p_O_DFFX1serial_div_),.p_desc1412_p_O_DFFX1(p_desc1412_p_O_DFFX1serial_div_),.p_desc1413_p_O_DFFX1(p_desc1413_p_O_DFFX1serial_div_),.p_desc1414_p_O_DFFX1(p_desc1414_p_O_DFFX1serial_div_),.p_desc1415_p_O_DFFX1(p_desc1415_p_O_DFFX1serial_div_),.p_desc1416_p_O_DFFX1(p_desc1416_p_O_DFFX1serial_div_),.p_desc1417_p_O_DFFX1(p_desc1417_p_O_DFFX1serial_div_),.p_desc1418_p_O_DFFX1(p_desc1418_p_O_DFFX1serial_div_),.p_desc1419_p_O_DFFX1(p_desc1419_p_O_DFFX1serial_div_),.p_desc1420_p_O_DFFX1(p_desc1420_p_O_DFFX1serial_div_),.p_desc1421_p_O_DFFX1(p_desc1421_p_O_DFFX1serial_div_),.p_desc1422_p_O_DFFX1(p_desc1422_p_O_DFFX1serial_div_),.p_desc1423_p_O_DFFX1(p_desc1423_p_O_DFFX1serial_div_),.p_desc1424_p_O_DFFX1(p_desc1424_p_O_DFFX1serial_div_),.p_desc1425_p_O_DFFX1(p_desc1425_p_O_DFFX1serial_div_),.p_desc1426_p_O_DFFX1(p_desc1426_p_O_DFFX1serial_div_),.p_desc1427_p_O_DFFX1(p_desc1427_p_O_DFFX1serial_div_),.p_desc1428_p_O_DFFX1(p_desc1428_p_O_DFFX1serial_div_),.p_desc1429_p_O_DFFX1(p_desc1429_p_O_DFFX1serial_div_),.p_desc1430_p_O_DFFX1(p_desc1430_p_O_DFFX1serial_div_),.p_desc1431_p_O_DFFX1(p_desc1431_p_O_DFFX1serial_div_),.p_desc1432_p_O_DFFX1(p_desc1432_p_O_DFFX1serial_div_),.p_desc1433_p_O_DFFX1(p_desc1433_p_O_DFFX1serial_div_),.p_desc1434_p_O_DFFX1(p_desc1434_p_O_DFFX1serial_div_),.p_desc1435_p_O_DFFX1(p_desc1435_p_O_DFFX1serial_div_),.p_desc1436_p_O_DFFX1(p_desc1436_p_O_DFFX1serial_div_),.p_desc1437_p_O_DFFX1(p_desc1437_p_O_DFFX1serial_div_),.p_desc1438_p_O_DFFX1(p_desc1438_p_O_DFFX1serial_div_),.p_desc1439_p_O_DFFX1(p_desc1439_p_O_DFFX1serial_div_),.p_desc1440_p_O_DFFX1(p_desc1440_p_O_DFFX1serial_div_),.p_desc1441_p_O_DFFX1(p_desc1441_p_O_DFFX1serial_div_),.p_desc1442_p_O_DFFX1(p_desc1442_p_O_DFFX1serial_div_),.p_desc1443_p_O_DFFX1(p_desc1443_p_O_DFFX1serial_div_),.p_desc1444_p_O_DFFX1(p_desc1444_p_O_DFFX1serial_div_),.p_s_start_i_reg_p_O_DFFX1(p_s_start_i_reg_p_O_DFFX1serial_div_),.p_s_ready_o_reg_p_O_DFFX1(p_s_ready_o_reg_p_O_DFFX1serial_div_),.p_desc1445_p_O_DFFX1(p_desc1445_p_O_DFFX1serial_div_),.p_desc1446_p_O_DFFX1(p_desc1446_p_O_DFFX1serial_div_),.p_desc1447_p_O_DFFX1(p_desc1447_p_O_DFFX1serial_div_),.p_desc1448_p_O_DFFX1(p_desc1448_p_O_DFFX1serial_div_),.p_desc1449_p_O_DFFX1(p_desc1449_p_O_DFFX1serial_div_),.p_desc1450_p_O_DFFX1(p_desc1450_p_O_DFFX1serial_div_),.p_desc1451_p_O_DFFX1(p_desc1451_p_O_DFFX1serial_div_),.p_desc1452_p_O_DFFX1(p_desc1452_p_O_DFFX1serial_div_),.p_desc1453_p_O_DFFX1(p_desc1453_p_O_DFFX1serial_div_),.p_desc1454_p_O_DFFX1(p_desc1454_p_O_DFFX1serial_div_),.p_desc1455_p_O_DFFX1(p_desc1455_p_O_DFFX1serial_div_),.p_desc1456_p_O_DFFX1(p_desc1456_p_O_DFFX1serial_div_),.p_desc1457_p_O_DFFX1(p_desc1457_p_O_DFFX1serial_div_),.p_desc1458_p_O_DFFX1(p_desc1458_p_O_DFFX1serial_div_),.p_desc1459_p_O_DFFX1(p_desc1459_p_O_DFFX1serial_div_),.p_desc1460_p_O_DFFX1(p_desc1460_p_O_DFFX1serial_div_),.p_desc1461_p_O_DFFX1(p_desc1461_p_O_DFFX1serial_div_),.p_desc1462_p_O_DFFX1(p_desc1462_p_O_DFFX1serial_div_),.p_desc1463_p_O_DFFX1(p_desc1463_p_O_DFFX1serial_div_),.p_desc1464_p_O_DFFX1(p_desc1464_p_O_DFFX1serial_div_),.p_desc1465_p_O_DFFX1(p_desc1465_p_O_DFFX1serial_div_),.p_desc1466_p_O_DFFX1(p_desc1466_p_O_DFFX1serial_div_),.p_desc1467_p_O_DFFX1(p_desc1467_p_O_DFFX1serial_div_),.p_desc1468_p_O_DFFX1(p_desc1468_p_O_DFFX1serial_div_),.p_desc1469_p_O_DFFX1(p_desc1469_p_O_DFFX1serial_div_),.p_desc1470_p_O_DFFX1(p_desc1470_p_O_DFFX1serial_div_),.p_desc1471_p_O_DFFX1(p_desc1471_p_O_DFFX1serial_div_),.p_desc1472_p_O_DFFX1(p_desc1472_p_O_DFFX1serial_div_),.p_desc1473_p_O_DFFX1(p_desc1473_p_O_DFFX1serial_div_),.p_desc1474_p_O_DFFX1(p_desc1474_p_O_DFFX1serial_div_),.p_desc1475_p_O_DFFX1(p_desc1475_p_O_DFFX1serial_div_),.p_desc1476_p_O_DFFX1(p_desc1476_p_O_DFFX1serial_div_),.p_desc1477_p_O_DFFX1(p_desc1477_p_O_DFFX1serial_div_),.p_desc1478_p_O_DFFX1(p_desc1478_p_O_DFFX1serial_div_),.p_desc1479_p_O_DFFX1(p_desc1479_p_O_DFFX1serial_div_),.p_desc1480_p_O_DFFX1(p_desc1480_p_O_DFFX1serial_div_),.p_desc1481_p_O_DFFX1(p_desc1481_p_O_DFFX1serial_div_),.p_desc1482_p_O_DFFX1(p_desc1482_p_O_DFFX1serial_div_),.p_desc1483_p_O_DFFX1(p_desc1483_p_O_DFFX1serial_div_),.p_desc1484_p_O_DFFX1(p_desc1484_p_O_DFFX1serial_div_),.p_desc1485_p_O_DFFX1(p_desc1485_p_O_DFFX1serial_div_),.p_desc1486_p_O_DFFX1(p_desc1486_p_O_DFFX1serial_div_),.p_desc1487_p_O_DFFX1(p_desc1487_p_O_DFFX1serial_div_),.p_desc1488_p_O_DFFX1(p_desc1488_p_O_DFFX1serial_div_),.p_desc1489_p_O_DFFX1(p_desc1489_p_O_DFFX1serial_div_),.p_desc1490_p_O_DFFX1(p_desc1490_p_O_DFFX1serial_div_),.p_desc1491_p_O_DFFX1(p_desc1491_p_O_DFFX1serial_div_),.p_desc1492_p_O_DFFX1(p_desc1492_p_O_DFFX1serial_div_),.p_desc1493_p_O_DFFX1(p_desc1493_p_O_DFFX1serial_div_),.p_desc1494_p_O_DFFX1(p_desc1494_p_O_DFFX1serial_div_),.p_desc1495_p_O_DFFX1(p_desc1495_p_O_DFFX1serial_div_),.p_desc1496_p_O_DFFX1(p_desc1496_p_O_DFFX1serial_div_),.p_desc1497_p_O_DFFX1(p_desc1497_p_O_DFFX1serial_div_),.p_desc1498_p_O_DFFX1(p_desc1498_p_O_DFFX1serial_div_),.p_desc1499_p_O_DFFX1(p_desc1499_p_O_DFFX1serial_div_),.p_desc1500_p_O_DFFX1(p_desc1500_p_O_DFFX1serial_div_),.p_desc1501_p_O_DFFX1(p_desc1501_p_O_DFFX1serial_div_),.p_desc1502_p_O_DFFX1(p_desc1502_p_O_DFFX1serial_div_),.p_desc1503_p_O_DFFX1(p_desc1503_p_O_DFFX1serial_div_),.p_desc1504_p_O_DFFX1(p_desc1504_p_O_DFFX1serial_div_),.p_desc1505_p_O_DFFX1(p_desc1505_p_O_DFFX1serial_div_),.p_desc1506_p_O_DFFX1(p_desc1506_p_O_DFFX1serial_div_),.p_desc1507_p_O_DFFX1(p_desc1507_p_O_DFFX1serial_div_),.p_desc1508_p_O_DFFX1(p_desc1508_p_O_DFFX1serial_div_),.p_desc1509_p_O_DFFX1(p_desc1509_p_O_DFFX1serial_div_),.p_desc1510_p_O_DFFX1(p_desc1510_p_O_DFFX1serial_div_),.p_desc1511_p_O_DFFX1(p_desc1511_p_O_DFFX1serial_div_),.p_desc1512_p_O_DFFX1(p_desc1512_p_O_DFFX1serial_div_),.p_desc1513_p_O_DFFX1(p_desc1513_p_O_DFFX1serial_div_),.p_desc1514_p_O_DFFX1(p_desc1514_p_O_DFFX1serial_div_),.p_desc1515_p_O_DFFX1(p_desc1515_p_O_DFFX1serial_div_),.p_desc1516_p_O_DFFX1(p_desc1516_p_O_DFFX1serial_div_),.p_desc1517_p_O_DFFX1(p_desc1517_p_O_DFFX1serial_div_),.p_desc1518_p_O_DFFX1(p_desc1518_p_O_DFFX1serial_div_),.p_desc1519_p_O_DFFX1(p_desc1519_p_O_DFFX1serial_div_),.p_desc1520_p_O_DFFX1(p_desc1520_p_O_DFFX1serial_div_),.p_desc1521_p_O_DFFX1(p_desc1521_p_O_DFFX1serial_div_),.p_desc1522_p_O_DFFX1(p_desc1522_p_O_DFFX1serial_div_),.p_desc1523_p_O_DFFX1(p_desc1523_p_O_DFFX1serial_div_),.p_desc1524_p_O_DFFX1(p_desc1524_p_O_DFFX1serial_div_),.p_desc1525_p_O_DFFX1(p_desc1525_p_O_DFFX1serial_div_),.p_desc1526_p_O_DFFX1(p_desc1526_p_O_DFFX1serial_div_),.p_desc1527_p_O_DFFX1(p_desc1527_p_O_DFFX1serial_div_),.p_desc1528_p_O_DFFX1(p_desc1528_p_O_DFFX1serial_div_),.p_s_state_reg_p_O_DFFX1(p_s_state_reg_p_O_DFFX1serial_div_),.p_desc1529_p_O_DFFX1(p_desc1529_p_O_DFFX1serial_div_));
  post_norm_div_inj i_post_norm_div(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n234,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n231,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.opb_i(s_opb_i),.qutnt_i(serial_div_qutnt),.rmndr_i(serial_div_rmndr),.exp_10_i(pre_norm_div_exp),.sign_i(serial_div_sign),.rmode_i(s_rmode_i),.output_o(post_norm_div_output),.ine_o(post_norm_div_ine),.p_desc1530_p_O_DFFX1(p_desc1530_p_O_DFFX1post_norm_div_),.p_desc1531_p_O_DFFX1(p_desc1531_p_O_DFFX1post_norm_div_),.p_desc1532_p_O_DFFX1(p_desc1532_p_O_DFFX1post_norm_div_),.p_desc1533_p_O_DFFX1(p_desc1533_p_O_DFFX1post_norm_div_),.p_desc1534_p_O_DFFX1(p_desc1534_p_O_DFFX1post_norm_div_),.p_desc1535_p_O_DFFX1(p_desc1535_p_O_DFFX1post_norm_div_),.p_desc1536_p_O_DFFX1(p_desc1536_p_O_DFFX1post_norm_div_),.p_desc1537_p_O_DFFX1(p_desc1537_p_O_DFFX1post_norm_div_),.p_desc1538_p_O_DFFX1(p_desc1538_p_O_DFFX1post_norm_div_),.p_desc1539_p_O_DFFX1(p_desc1539_p_O_DFFX1post_norm_div_),.p_desc1540_p_O_DFFX1(p_desc1540_p_O_DFFX1post_norm_div_),.p_desc1541_p_O_DFFX1(p_desc1541_p_O_DFFX1post_norm_div_),.p_desc1542_p_O_DFFX1(p_desc1542_p_O_DFFX1post_norm_div_),.p_desc1543_p_O_DFFX1(p_desc1543_p_O_DFFX1post_norm_div_),.p_desc1544_p_O_DFFX1(p_desc1544_p_O_DFFX1post_norm_div_),.p_desc1545_p_O_DFFX1(p_desc1545_p_O_DFFX1post_norm_div_),.p_desc1546_p_O_DFFX1(p_desc1546_p_O_DFFX1post_norm_div_),.p_desc1547_p_O_DFFX1(p_desc1547_p_O_DFFX1post_norm_div_),.p_desc1548_p_O_DFFX1(p_desc1548_p_O_DFFX1post_norm_div_),.p_desc1549_p_O_DFFX1(p_desc1549_p_O_DFFX1post_norm_div_),.p_desc1550_p_O_DFFX1(p_desc1550_p_O_DFFX1post_norm_div_),.p_desc1551_p_O_DFFX1(p_desc1551_p_O_DFFX1post_norm_div_),.p_desc1552_p_O_DFFX1(p_desc1552_p_O_DFFX1post_norm_div_),.p_desc1553_p_O_DFFX1(p_desc1553_p_O_DFFX1post_norm_div_),.p_desc1554_p_O_DFFX1(p_desc1554_p_O_DFFX1post_norm_div_),.p_desc1555_p_O_DFFX1(p_desc1555_p_O_DFFX1post_norm_div_),.p_desc1556_p_O_DFFX1(p_desc1556_p_O_DFFX1post_norm_div_),.p_desc1557_p_O_DFFX1(p_desc1557_p_O_DFFX1post_norm_div_),.p_desc1558_p_O_DFFX1(p_desc1558_p_O_DFFX1post_norm_div_),.p_desc1559_p_O_DFFX1(p_desc1559_p_O_DFFX1post_norm_div_),.p_desc1560_p_O_DFFX1(p_desc1560_p_O_DFFX1post_norm_div_),.p_desc1561_p_O_DFFX1(p_desc1561_p_O_DFFX1post_norm_div_),.p_desc1562_p_O_DFFX1(p_desc1562_p_O_DFFX1post_norm_div_),.p_desc1563_p_O_DFFX1(p_desc1563_p_O_DFFX1post_norm_div_),.p_desc1564_p_O_DFFX1(p_desc1564_p_O_DFFX1post_norm_div_),.p_desc1565_p_O_DFFX1(p_desc1565_p_O_DFFX1post_norm_div_),.p_desc1566_p_O_DFFX1(p_desc1566_p_O_DFFX1post_norm_div_),.p_desc1567_p_O_DFFX1(p_desc1567_p_O_DFFX1post_norm_div_),.p_desc1568_p_O_DFFX1(p_desc1568_p_O_DFFX1post_norm_div_),.p_desc1569_p_O_DFFX1(p_desc1569_p_O_DFFX1post_norm_div_),.p_desc1570_p_O_DFFX1(p_desc1570_p_O_DFFX1post_norm_div_),.p_desc1571_p_O_DFFX1(p_desc1571_p_O_DFFX1post_norm_div_),.p_desc1572_p_O_DFFX1(p_desc1572_p_O_DFFX1post_norm_div_),.p_desc1573_p_O_DFFX1(p_desc1573_p_O_DFFX1post_norm_div_),.p_desc1574_p_O_DFFX1(p_desc1574_p_O_DFFX1post_norm_div_),.p_desc1575_p_O_DFFX1(p_desc1575_p_O_DFFX1post_norm_div_),.p_desc1576_p_O_DFFX1(p_desc1576_p_O_DFFX1post_norm_div_),.p_desc1577_p_O_DFFX1(p_desc1577_p_O_DFFX1post_norm_div_),.p_desc1578_p_O_DFFX1(p_desc1578_p_O_DFFX1post_norm_div_),.p_desc1579_p_O_DFFX1(p_desc1579_p_O_DFFX1post_norm_div_),.p_desc1580_p_O_DFFX1(p_desc1580_p_O_DFFX1post_norm_div_),.p_desc1581_p_O_DFFX1(p_desc1581_p_O_DFFX1post_norm_div_),.p_desc1582_p_O_DFFX1(p_desc1582_p_O_DFFX1post_norm_div_),.p_desc1583_p_O_DFFX1(p_desc1583_p_O_DFFX1post_norm_div_),.p_desc1584_p_O_DFFX1(p_desc1584_p_O_DFFX1post_norm_div_),.p_desc1585_p_O_DFFX1(p_desc1585_p_O_DFFX1post_norm_div_),.p_desc1586_p_O_DFFX1(p_desc1586_p_O_DFFX1post_norm_div_),.p_desc1587_p_O_DFFX1(p_desc1587_p_O_DFFX1post_norm_div_),.p_desc1588_p_O_DFFX1(p_desc1588_p_O_DFFX1post_norm_div_),.p_desc1589_p_O_DFFX1(p_desc1589_p_O_DFFX1post_norm_div_),.p_desc1590_p_O_DFFX1(p_desc1590_p_O_DFFX1post_norm_div_),.p_desc1591_p_O_DFFX1(p_desc1591_p_O_DFFX1post_norm_div_),.p_desc1592_p_O_DFFX1(p_desc1592_p_O_DFFX1post_norm_div_),.p_desc1593_p_O_DFFX1(p_desc1593_p_O_DFFX1post_norm_div_),.p_desc1594_p_O_DFFX1(p_desc1594_p_O_DFFX1post_norm_div_),.p_desc1595_p_O_DFFX1(p_desc1595_p_O_DFFX1post_norm_div_),.p_desc1596_p_O_DFFX1(p_desc1596_p_O_DFFX1post_norm_div_),.p_desc1597_p_O_DFFX1(p_desc1597_p_O_DFFX1post_norm_div_),.p_desc1598_p_O_DFFX1(p_desc1598_p_O_DFFX1post_norm_div_),.p_desc1599_p_O_DFFX1(p_desc1599_p_O_DFFX1post_norm_div_),.p_desc1600_p_O_DFFX1(p_desc1600_p_O_DFFX1post_norm_div_),.p_desc1601_p_O_DFFX1(p_desc1601_p_O_DFFX1post_norm_div_),.p_desc1602_p_O_DFFX1(p_desc1602_p_O_DFFX1post_norm_div_),.p_desc1603_p_O_DFFX1(p_desc1603_p_O_DFFX1post_norm_div_),.p_desc1604_p_O_DFFX1(p_desc1604_p_O_DFFX1post_norm_div_),.p_desc1605_p_O_DFFX1(p_desc1605_p_O_DFFX1post_norm_div_),.p_desc1606_p_O_DFFX1(p_desc1606_p_O_DFFX1post_norm_div_),.p_desc1607_p_O_DFFX1(p_desc1607_p_O_DFFX1post_norm_div_),.p_desc1608_p_O_DFFX1(p_desc1608_p_O_DFFX1post_norm_div_),.p_desc1609_p_O_DFFX1(p_desc1609_p_O_DFFX1post_norm_div_),.p_desc1610_p_O_DFFX1(p_desc1610_p_O_DFFX1post_norm_div_),.p_desc1611_p_O_DFFX1(p_desc1611_p_O_DFFX1post_norm_div_),.p_desc1612_p_O_DFFX1(p_desc1612_p_O_DFFX1post_norm_div_),.p_desc1613_p_O_DFFX1(p_desc1613_p_O_DFFX1post_norm_div_),.p_desc1614_p_O_DFFX1(p_desc1614_p_O_DFFX1post_norm_div_),.p_desc1615_p_O_DFFX1(p_desc1615_p_O_DFFX1post_norm_div_),.p_desc1616_p_O_DFFX1(p_desc1616_p_O_DFFX1post_norm_div_),.p_desc1617_p_O_DFFX1(p_desc1617_p_O_DFFX1post_norm_div_),.p_desc1618_p_O_DFFX1(p_desc1618_p_O_DFFX1post_norm_div_),.p_desc1619_p_O_DFFX1(p_desc1619_p_O_DFFX1post_norm_div_),.p_desc1620_p_O_DFFX1(p_desc1620_p_O_DFFX1post_norm_div_),.p_desc1621_p_O_DFFX1(p_desc1621_p_O_DFFX1post_norm_div_),.p_desc1622_p_O_DFFX1(p_desc1622_p_O_DFFX1post_norm_div_),.p_desc1623_p_O_DFFX1(p_desc1623_p_O_DFFX1post_norm_div_),.p_desc1624_p_O_DFFX1(p_desc1624_p_O_DFFX1post_norm_div_),.p_desc1625_p_O_DFFX1(p_desc1625_p_O_DFFX1post_norm_div_),.p_desc1626_p_O_DFFX1(p_desc1626_p_O_DFFX1post_norm_div_),.p_desc1627_p_O_DFFX1(p_desc1627_p_O_DFFX1post_norm_div_),.p_desc1628_p_O_DFFX1(p_desc1628_p_O_DFFX1post_norm_div_),.p_desc1629_p_O_DFFX1(p_desc1629_p_O_DFFX1post_norm_div_),.p_desc1630_p_O_DFFX1(p_desc1630_p_O_DFFX1post_norm_div_),.p_desc1631_p_O_DFFX1(p_desc1631_p_O_DFFX1post_norm_div_),.p_desc1632_p_O_DFFX1(p_desc1632_p_O_DFFX1post_norm_div_),.p_desc1633_p_O_DFFX1(p_desc1633_p_O_DFFX1post_norm_div_),.p_desc1634_p_O_DFFX1(p_desc1634_p_O_DFFX1post_norm_div_),.p_desc1635_p_O_DFFX1(p_desc1635_p_O_DFFX1post_norm_div_),.p_desc1636_p_O_DFFX1(p_desc1636_p_O_DFFX1post_norm_div_),.p_desc1637_p_O_DFFX1(p_desc1637_p_O_DFFX1post_norm_div_),.p_desc1638_p_O_DFFX1(p_desc1638_p_O_DFFX1post_norm_div_),.p_desc1639_p_O_DFFX1(p_desc1639_p_O_DFFX1post_norm_div_),.p_desc1640_p_O_DFFX1(p_desc1640_p_O_DFFX1post_norm_div_),.p_desc1641_p_O_DFFX1(p_desc1641_p_O_DFFX1post_norm_div_),.p_desc1642_p_O_DFFX1(p_desc1642_p_O_DFFX1post_norm_div_),.p_desc1643_p_O_DFFX1(p_desc1643_p_O_DFFX1post_norm_div_),.p_desc1644_p_O_DFFX1(p_desc1644_p_O_DFFX1post_norm_div_),.p_desc1645_p_O_DFFX1(p_desc1645_p_O_DFFX1post_norm_div_),.p_desc1646_p_O_DFFX1(p_desc1646_p_O_DFFX1post_norm_div_),.p_desc1647_p_O_DFFX1(p_desc1647_p_O_DFFX1post_norm_div_),.p_desc1648_p_O_DFFX1(p_desc1648_p_O_DFFX1post_norm_div_),.p_desc1649_p_O_DFFX1(p_desc1649_p_O_DFFX1post_norm_div_),.p_desc1650_p_O_DFFX1(p_desc1650_p_O_DFFX1post_norm_div_),.p_desc1651_p_O_DFFX1(p_desc1651_p_O_DFFX1post_norm_div_),.p_s_sign_i_reg_p_O_DFFX1(p_s_sign_i_reg_p_O_DFFX1post_norm_div_),.p_desc1652_p_O_DFFX1(p_desc1652_p_O_DFFX1post_norm_div_),.p_desc1653_p_O_DFFX1(p_desc1653_p_O_DFFX1post_norm_div_),.p_desc1654_p_O_DFFX1(p_desc1654_p_O_DFFX1post_norm_div_),.p_desc1658_p_O_DFFX1(p_desc1658_p_O_DFFX1post_norm_div_),.p_desc1659_p_O_DFFX1(p_desc1659_p_O_DFFX1post_norm_div_),.p_desc1663_p_O_DFFX1(p_desc1663_p_O_DFFX1post_norm_div_),.p_desc1664_p_O_DFFX1(p_desc1664_p_O_DFFX1post_norm_div_),.p_desc1665_p_O_DFFX1(p_desc1665_p_O_DFFX1post_norm_div_),.p_desc1666_p_O_DFFX1(p_desc1666_p_O_DFFX1post_norm_div_),.p_desc1667_p_O_DFFX1(p_desc1667_p_O_DFFX1post_norm_div_),.p_desc1668_p_O_DFFX1(p_desc1668_p_O_DFFX1post_norm_div_),.p_desc1669_p_O_DFFX1(p_desc1669_p_O_DFFX1post_norm_div_),.p_desc1670_p_O_DFFX1(p_desc1670_p_O_DFFX1post_norm_div_),.p_desc1671_p_O_DFFX1(p_desc1671_p_O_DFFX1post_norm_div_),.p_desc1672_p_O_DFFX1(p_desc1672_p_O_DFFX1post_norm_div_),.p_desc1673_p_O_DFFX1(p_desc1673_p_O_DFFX1post_norm_div_),.p_desc1674_p_O_DFFX1(p_desc1674_p_O_DFFX1post_norm_div_),.p_desc1675_p_O_DFFX1(p_desc1675_p_O_DFFX1post_norm_div_),.p_desc1676_p_O_DFFX1(p_desc1676_p_O_DFFX1post_norm_div_),.p_desc1677_p_O_DFFX1(p_desc1677_p_O_DFFX1post_norm_div_),.p_desc1678_p_O_DFFX1(p_desc1678_p_O_DFFX1post_norm_div_),.p_desc1679_p_O_DFFX1(p_desc1679_p_O_DFFX1post_norm_div_),.p_desc1680_p_O_DFFX1(p_desc1680_p_O_DFFX1post_norm_div_),.p_desc1681_p_O_DFFX1(p_desc1681_p_O_DFFX1post_norm_div_),.p_desc1682_p_O_DFFX1(p_desc1682_p_O_DFFX1post_norm_div_),.p_desc1683_p_O_DFFX1(p_desc1683_p_O_DFFX1post_norm_div_),.p_desc1684_p_O_DFFX1(p_desc1684_p_O_DFFX1post_norm_div_),.p_desc1685_p_O_DFFX1(p_desc1685_p_O_DFFX1post_norm_div_),.p_desc1686_p_O_DFFX1(p_desc1686_p_O_DFFX1post_norm_div_),.p_desc1687_p_O_DFFX1(p_desc1687_p_O_DFFX1post_norm_div_),.p_desc1688_p_O_DFFX1(p_desc1688_p_O_DFFX1post_norm_div_),.p_desc1689_p_O_DFFX1(p_desc1689_p_O_DFFX1post_norm_div_),.p_desc1690_p_O_DFFX1(p_desc1690_p_O_DFFX1post_norm_div_),.p_desc1691_p_O_DFFX1(p_desc1691_p_O_DFFX1post_norm_div_),.p_desc1692_p_O_DFFX1(p_desc1692_p_O_DFFX1post_norm_div_),.p_desc1693_p_O_DFFX1(p_desc1693_p_O_DFFX1post_norm_div_),.p_desc1694_p_O_DFFX1(p_desc1694_p_O_DFFX1post_norm_div_),.p_desc1695_p_O_DFFX1(p_desc1695_p_O_DFFX1post_norm_div_),.p_desc1696_p_O_DFFX1(p_desc1696_p_O_DFFX1post_norm_div_),.p_desc1697_p_O_DFFX1(p_desc1697_p_O_DFFX1post_norm_div_),.p_desc1698_p_O_DFFX1(p_desc1698_p_O_DFFX1post_norm_div_),.p_desc1699_p_O_DFFX1(p_desc1699_p_O_DFFX1post_norm_div_),.p_desc1700_p_O_DFFX1(p_desc1700_p_O_DFFX1post_norm_div_),.p_desc1701_p_O_DFFX1(p_desc1701_p_O_DFFX1post_norm_div_),.p_desc1702_p_O_DFFX1(p_desc1702_p_O_DFFX1post_norm_div_),.p_desc1703_p_O_DFFX1(p_desc1703_p_O_DFFX1post_norm_div_),.p_desc1704_p_O_DFFX1(p_desc1704_p_O_DFFX1post_norm_div_),.p_desc1705_p_O_DFFX1(p_desc1705_p_O_DFFX1post_norm_div_),.p_desc1706_p_O_DFFX1(p_desc1706_p_O_DFFX1post_norm_div_),.p_desc1707_p_O_DFFX1(p_desc1707_p_O_DFFX1post_norm_div_),.p_desc1708_p_O_DFFX1(p_desc1708_p_O_DFFX1post_norm_div_),.p_desc1709_p_O_DFFX1(p_desc1709_p_O_DFFX1post_norm_div_),.p_desc1710_p_O_DFFX1(p_desc1710_p_O_DFFX1post_norm_div_),.p_desc1711_p_O_DFFX1(p_desc1711_p_O_DFFX1post_norm_div_),.p_desc1712_p_O_DFFX1(p_desc1712_p_O_DFFX1post_norm_div_),.p_desc1713_p_O_DFFX1(p_desc1713_p_O_DFFX1post_norm_div_),.p_desc1714_p_O_DFFX1(p_desc1714_p_O_DFFX1post_norm_div_),.p_desc1715_p_O_DFFX1(p_desc1715_p_O_DFFX1post_norm_div_),.p_desc1716_p_O_DFFX1(p_desc1716_p_O_DFFX1post_norm_div_),.p_desc1717_p_O_DFFX1(p_desc1717_p_O_DFFX1post_norm_div_),.p_desc1718_p_O_DFFX1(p_desc1718_p_O_DFFX1post_norm_div_),.p_desc1719_p_O_DFFX1(p_desc1719_p_O_DFFX1post_norm_div_),.p_desc1720_p_O_DFFX1(p_desc1720_p_O_DFFX1post_norm_div_),.p_desc1721_p_O_DFFX1(p_desc1721_p_O_DFFX1post_norm_div_),.p_desc1722_p_O_DFFX1(p_desc1722_p_O_DFFX1post_norm_div_),.p_desc1723_p_O_DFFX1(p_desc1723_p_O_DFFX1post_norm_div_),.p_desc1724_p_O_DFFX1(p_desc1724_p_O_DFFX1post_norm_div_),.p_desc1725_p_O_DFFX1(p_desc1725_p_O_DFFX1post_norm_div_),.p_desc1726_p_O_DFFX1(p_desc1726_p_O_DFFX1post_norm_div_),.p_desc1727_p_O_DFFX1(p_desc1727_p_O_DFFX1post_norm_div_),.p_desc1728_p_O_DFFX1(p_desc1728_p_O_DFFX1post_norm_div_),.p_ine_o_reg_p_O_DFFX1(p_ine_o_reg_p_O_DFFX1post_norm_div_),.p_desc1729_p_O_DFFX1(p_desc1729_p_O_DFFX1post_norm_div_),.p_desc1737_p_O_DFFX1(p_desc1737_p_O_DFFX1post_norm_div_),.p_desc1738_p_O_DFFX1(p_desc1738_p_O_DFFX1post_norm_div_),.p_desc1739_p_O_DFFX1(p_desc1739_p_O_DFFX1post_norm_div_),.p_desc1740_p_O_DFFX1(p_desc1740_p_O_DFFX1post_norm_div_),.p_desc1741_p_O_DFFX1(p_desc1741_p_O_DFFX1post_norm_div_),.p_desc1742_p_O_DFFX1(p_desc1742_p_O_DFFX1post_norm_div_),.p_desc1743_p_O_DFFX1(p_desc1743_p_O_DFFX1post_norm_div_),.p_desc1744_p_O_DFFX1(p_desc1744_p_O_DFFX1post_norm_div_),.p_desc1745_p_O_DFFX1(p_desc1745_p_O_DFFX1post_norm_div_),.p_desc1746_p_O_DFFX1(p_desc1746_p_O_DFFX1post_norm_div_),.p_desc1747_p_O_DFFX1(p_desc1747_p_O_DFFX1post_norm_div_),.p_desc1748_p_O_DFFX1(p_desc1748_p_O_DFFX1post_norm_div_),.p_desc1749_p_O_DFFX1(p_desc1749_p_O_DFFX1post_norm_div_),.p_desc1750_p_O_DFFX1(p_desc1750_p_O_DFFX1post_norm_div_),.p_desc1751_p_O_DFFX1(p_desc1751_p_O_DFFX1post_norm_div_),.p_desc1752_p_O_DFFX1(p_desc1752_p_O_DFFX1post_norm_div_),.p_desc1753_p_O_DFFX1(p_desc1753_p_O_DFFX1post_norm_div_),.p_desc1754_p_O_DFFX1(p_desc1754_p_O_DFFX1post_norm_div_),.p_desc1755_p_O_DFFX1(p_desc1755_p_O_DFFX1post_norm_div_),.p_desc1756_p_O_DFFX1(p_desc1756_p_O_DFFX1post_norm_div_),.p_desc1757_p_O_DFFX1(p_desc1757_p_O_DFFX1post_norm_div_),.p_desc1758_p_O_DFFX1(p_desc1758_p_O_DFFX1post_norm_div_),.p_desc1849_p_O_DFFX1(p_desc1849_p_O_DFFX1post_norm_div_),.p_desc1850_p_O_DFFX1(p_desc1850_p_O_DFFX1post_norm_div_),.p_desc1851_p_O_DFFX1(p_desc1851_p_O_DFFX1post_norm_div_),.p_desc1852_p_O_DFFX1(p_desc1852_p_O_DFFX1post_norm_div_),.p_desc1853_p_O_DFFX1(p_desc1853_p_O_DFFX1post_norm_div_),.p_desc1854_p_O_DFFX1(p_desc1854_p_O_DFFX1post_norm_div_),.p_desc1855_p_O_DFFX1(p_desc1855_p_O_DFFX1post_norm_div_),.p_desc1856_p_O_DFFX1(p_desc1856_p_O_DFFX1post_norm_div_),.p_desc1857_p_O_DFFX1(p_desc1857_p_O_DFFX1post_norm_div_),.p_desc1858_p_O_DFFX1(p_desc1858_p_O_DFFX1post_norm_div_),.p_desc1859_p_O_DFFX1(p_desc1859_p_O_DFFX1post_norm_div_),.p_desc1860_p_O_DFFX1(p_desc1860_p_O_DFFX1post_norm_div_),.p_desc1861_p_O_DFFX1(p_desc1861_p_O_DFFX1post_norm_div_),.p_desc1862_p_O_DFFX1(p_desc1862_p_O_DFFX1post_norm_div_),.p_desc1863_p_O_DFFX1(p_desc1863_p_O_DFFX1post_norm_div_),.p_desc1864_p_O_DFFX1(p_desc1864_p_O_DFFX1post_norm_div_),.p_desc1865_p_O_DFFX1(p_desc1865_p_O_DFFX1post_norm_div_),.p_desc1866_p_O_DFFX1(p_desc1866_p_O_DFFX1post_norm_div_),.p_desc1867_p_O_DFFX1(p_desc1867_p_O_DFFX1post_norm_div_),.p_desc1868_p_O_DFFX1(p_desc1868_p_O_DFFX1post_norm_div_),.p_desc1869_p_O_DFFX1(p_desc1869_p_O_DFFX1post_norm_div_));
  pre_norm_sqrt_inj i_pre_norm_sqrt(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n233,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n230,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.fracta_52_o({pre_norm_sqrt_fracta_o[51:27],SYNOPSYS_UNCONNECTED__31,SYNOPSYS_UNCONNECTED__32,SYNOPSYS_UNCONNECTED__33,SYNOPSYS_UNCONNECTED__34,SYNOPSYS_UNCONNECTED__35,SYNOPSYS_UNCONNECTED__36,SYNOPSYS_UNCONNECTED__37,SYNOPSYS_UNCONNECTED__38,SYNOPSYS_UNCONNECTED__39,SYNOPSYS_UNCONNECTED__40,SYNOPSYS_UNCONNECTED__41,SYNOPSYS_UNCONNECTED__42,SYNOPSYS_UNCONNECTED__43,SYNOPSYS_UNCONNECTED__44,SYNOPSYS_UNCONNECTED__45,SYNOPSYS_UNCONNECTED__46,SYNOPSYS_UNCONNECTED__47,SYNOPSYS_UNCONNECTED__48,SYNOPSYS_UNCONNECTED__49,SYNOPSYS_UNCONNECTED__50,SYNOPSYS_UNCONNECTED__51,SYNOPSYS_UNCONNECTED__52,SYNOPSYS_UNCONNECTED__53,SYNOPSYS_UNCONNECTED__54,SYNOPSYS_UNCONNECTED__55,SYNOPSYS_UNCONNECTED__56,SYNOPSYS_UNCONNECTED__57}),.exp_o(pre_norm_sqrt_exp_o));
  sqrt_RD_WIDTH52_SQ_WIDTH26_inj i_sqrt(.clk_i(clk_i),.rad_i({pre_norm_sqrt_fracta_o[51:27],1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0}),.start_i(s_start_i),.sqr_o(sqrt_sqr_o),.ine_o(sqrt_ine_o));
  post_norm_sqrt_inj i_post_norm_sqrt(.clk_i(clk_i),.opa_i({s_opa_i[31:31],n229,n270,s_opa_i[28:24],n269,s_opa_i[22:21],n233,s_opa_i[19:19],n268,n267,n266,n265,n264,n263,n230,n262,n261,n260,n259,n258,n257,n256,n255,n254,n253,n252,s_opa_i[0:0]}),.fract_26_i(sqrt_sqr_o),.exp_i(pre_norm_sqrt_exp_o),.ine_i(sqrt_ine_o),.rmode_i(s_rmode_i),.output_o(post_norm_sqrt_output),.ine_o(post_norm_sqrt_ine_o));
  fpu_DW01_inc_0_inj add_392(.A(s_count),.SUM({N66,N65,N64,N63,N62,N61,N60,N59,N58,N57,N56,N55,N54,N53,N52,N51,N50,N49,N48,N47,N46,N45,N44,N43,N42,N41,N40,N39,N38,N37,N36,N35}));
  DELLN1X2 U232(.INP(n29),.Z(n250));
  OAI22X2 U233(.IN1(n221),.IN2(n222),.IN3(n223),.IN4(s_count[5:5]),.QN(n1));
  NAND2X1 U234(.IN1(n219),.IN2(n220),.QN(s_output_o[31:31]));
  NAND4X0 U235(.IN1(n9),.IN2(s_rmode_i[0:0]),.IN3(n199),.IN4(n10),.QN(n220));
  NBUFFX2 U236(.INP(n271),.Z(n229));
  NBUFFX2 U237(.INP(n271),.Z(n228));
  INVX0 U238(.INP(n3),.ZN(n272));
  NOR2X0 U239(.IN1(n272),.IN2(n207),.QN(s_output_o[23:23]));
  NBUFFX2 U240(.INP(n30),.Z(n248));
  NBUFFX2 U241(.INP(n30),.Z(n247));
  INVX0 U242(.INP(n1),.ZN(n273));
  NAND2X1 U243(.IN1(n209),.IN2(n202),.QN(n67));
  NBUFFX2 U244(.INP(n30),.Z(n249));
  NAND2X1 U245(.IN1(n209),.IN2(n3),.QN(s_output_o[0:0]));
  NAND2X1 U246(.IN1(n202),.IN2(n3),.QN(s_output_o[10:10]));
  NAND2X1 U247(.IN1(n200),.IN2(n3),.QN(s_output_o[17:17]));
  NAND2X1 U248(.IN1(n211),.IN2(n3),.QN(s_output_o[18:18]));
  NAND2X1 U249(.IN1(n204),.IN2(n3),.QN(s_output_o[19:19]));
  NAND2X1 U250(.IN1(n210),.IN2(n3),.QN(s_output_o[1:1]));
  NAND2X1 U251(.IN1(n203),.IN2(n3),.QN(s_output_o[20:20]));
  NAND2X1 U252(.IN1(n214),.IN2(n3),.QN(s_output_o[22:22]));
  NAND2X1 U253(.IN1(n201),.IN2(n3),.QN(s_output_o[7:7]));
  NAND2X1 U254(.IN1(n212),.IN2(n3),.QN(s_output_o[8:8]));
  NAND2X1 U255(.IN1(n205),.IN2(n3),.QN(s_output_o[9:9]));
  NBUFFX2 U256(.INP(n29),.Z(n251));
  NOR2X0 U257(.IN1(n59),.IN2(n217),.QN(N546));
  NOR2X0 U258(.IN1(n28),.IN2(n217),.QN(N547));
  NBUFFX2 U259(.INP(n48),.Z(n237));
  NBUFFX2 U260(.INP(n47),.Z(n239));
  NBUFFX2 U261(.INP(n48),.Z(n236));
  NBUFFX2 U262(.INP(n40),.Z(n244));
  NBUFFX2 U263(.INP(n40),.Z(n245));
  NBUFFX2 U264(.INP(n42),.Z(n241));
  NBUFFX2 U265(.INP(n42),.Z(n242));
  NBUFFX2 U266(.INP(n47),.Z(n240));
  NBUFFX2 U267(.INP(n48),.Z(n238));
  NBUFFX2 U268(.INP(n40),.Z(n246));
  NBUFFX2 U269(.INP(n42),.Z(n243));
  NBUFFX2 U270(.INP(s_opa_i[20:20]),.Z(n233));
  NBUFFX2 U271(.INP(s_opa_i[20:20]),.Z(n234));
  NAND3X0 U272(.IN1(n276),.IN2(n24),.IN3(n9),.QN(n3));
  INVX0 U273(.INP(n28),.ZN(n276));
  NAND2X0 U274(.IN1(s_rmode_i[1:1]),.IN2(s_output1[31:31]),.QN(n27));
  NBUFFX2 U275(.INP(s_opa_i[23:23]),.Z(n269));
  NOR2X0 U276(.IN1(n153),.IN2(n154),.QN(n78));
  NBUFFX2 U277(.INP(s_opa_i[29:29]),.Z(n270));
  NAND2X1 U278(.IN1(n210),.IN2(n203),.QN(n65));
  DELLN1X2 U279(.INP(s_opa_i[12:12]),.Z(n230));
  NBUFFX2 U280(.INP(s_opa_i[12:12]),.Z(n231));
  AND4X1 U281(.IN1(n41),.IN2(n45),.IN3(n206),.IN4(n213),.Q(n222));
  AOI21X1 U282(.IN1(n37),.IN2(n38),.IN3(n206),.QN(n223));
  NBUFFX2 U283(.INP(s_opa_i[15:15]),.Z(n265));
  NBUFFX2 U284(.INP(s_opa_i[17:17]),.Z(n267));
  NBUFFX2 U285(.INP(s_opa_i[18:18]),.Z(n268));
  NOR2X0 U286(.IN1(s_count[3:3]),.IN2(s_count[0:0]),.QN(n43));
  NBUFFX4 U287(.INP(s_opa_i[14:14]),.Z(n264));
  NBUFFX4 U288(.INP(s_opa_i[6:6]),.Z(n257));
  NBUFFX4 U289(.INP(s_opa_i[16:16]),.Z(n266));
  NBUFFX2 U290(.INP(s_opa_i[2:2]),.Z(n253));
  NBUFFX2 U291(.INP(s_opa_i[3:3]),.Z(n254));
  NBUFFX2 U292(.INP(s_opa_i[11:11]),.Z(n262));
  NBUFFX2 U293(.INP(s_opa_i[12:12]),.Z(n232));
  OR4X1 U294(.IN1(n224),.IN2(n225),.IN3(n226),.IN4(n227),.Q(n28));
  NAND2X0 U295(.IN1(s_output_o[27:27]),.IN2(s_output_o[28:28]),.QN(n226));
  NAND4X0 U296(.IN1(s_output1[23:23]),.IN2(s_output_o[24:24]),.IN3(s_output_o[25:25]),.IN4(s_output_o[26:26]),.QN(n227));
  NAND2X0 U297(.IN1(n68),.IN2(n69),.QN(N581));
  NBUFFX2 U298(.INP(s_opa_i[4:4]),.Z(n255));
  NBUFFX2 U299(.INP(s_opa_i[8:8]),.Z(n259));
  NBUFFX2 U300(.INP(s_opa_i[9:9]),.Z(n260));
  NBUFFX2 U301(.INP(s_opa_i[7:7]),.Z(n258));
  NBUFFX2 U302(.INP(s_opa_i[1:1]),.Z(n252));
  NBUFFX2 U303(.INP(s_opa_i[5:5]),.Z(n256));
  NOR2X0 U304(.IN1(n157),.IN2(n158),.QN(n88));
  NBUFFX2 U305(.INP(s_opa_i[20:20]),.Z(n235));
  NOR2X0 U306(.IN1(s_opa_i[31:31]),.IN2(n13),.QN(n11));
  NOR2X0 U307(.IN1(s_output_o[26:26]),.IN2(s_output_o[25:25]),.QN(n94));
  INVX0 U308(.INP(fpu_op_i[1:1]),.ZN(n275));
  NOR2X0 U309(.IN1(fpu_op_i[1:1]),.IN2(fpu_op_i[2:2]),.QN(n42));
  INVX0 U310(.INP(fpu_op_i[2:2]),.ZN(n274));
  DELLN1X2 U311(.INP(s_opa_i[10:10]),.Z(n261));
  DELLN1X2 U312(.INP(s_opa_i[13:13]),.Z(n263));
  DELLN1X2 U313(.INP(s_opa_i[30:30]),.Z(n271));
endmodule
