`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[441:0] injectionVector;
fpu_inj toplevel_instance (
.opa_i(testVector [31:0]),
.opb_i(testVector [63:32]),
.fpu_op_i(testVector [66:64]),
.rmode_i(testVector [68:67]),
.output_o(resultVector [31:0]),
.clk_i(clk),
.start_i(testVector[69]),
.ready_o(resultVector[32]),
.ine_o(resultVector[33]),
.overflow_o(resultVector[34]),
.underflow_o(resultVector[35]),
.div_zero_o(resultVector[36]),
.inf_o(resultVector[37]),
.zero_o(resultVector[38]),
.qnan_o(resultVector[39]),
.snan_o(resultVector[40]),
.p_desc1176_p_O_DFFX1pre_norm_div_(injectionVector[0]),
.p_desc1177_p_O_DFFX1pre_norm_div_(injectionVector[1]),
.p_desc1178_p_O_DFFX1pre_norm_div_(injectionVector[2]),
.p_desc1179_p_O_DFFX1pre_norm_div_(injectionVector[3]),
.p_desc1180_p_O_DFFX1pre_norm_div_(injectionVector[4]),
.p_desc1181_p_O_DFFX1pre_norm_div_(injectionVector[5]),
.p_desc1182_p_O_DFFX1pre_norm_div_(injectionVector[6]),
.p_desc1183_p_O_DFFX1pre_norm_div_(injectionVector[7]),
.p_desc1184_p_O_DFFX1pre_norm_div_(injectionVector[8]),
.p_desc1185_p_O_DFFX1pre_norm_div_(injectionVector[9]),
.p_desc1186_p_O_DFFX1pre_norm_div_(injectionVector[10]),
.p_desc1187_p_O_DFFX1pre_norm_div_(injectionVector[11]),
.p_desc1188_p_O_DFFX1pre_norm_div_(injectionVector[12]),
.p_desc1189_p_O_DFFX1pre_norm_div_(injectionVector[13]),
.p_desc1190_p_O_DFFX1pre_norm_div_(injectionVector[14]),
.p_desc1191_p_O_DFFX1pre_norm_div_(injectionVector[15]),
.p_desc1192_p_O_DFFX1pre_norm_div_(injectionVector[16]),
.p_desc1193_p_O_DFFX1pre_norm_div_(injectionVector[17]),
.p_desc1194_p_O_DFFX1pre_norm_div_(injectionVector[18]),
.p_desc1195_p_O_DFFX1pre_norm_div_(injectionVector[19]),
.p_desc1196_p_O_DFFX1pre_norm_div_(injectionVector[20]),
.p_desc1197_p_O_DFFX1pre_norm_div_(injectionVector[21]),
.p_desc1198_p_O_DFFX1pre_norm_div_(injectionVector[22]),
.p_desc1199_p_O_DFFX1pre_norm_div_(injectionVector[23]),
.p_desc1200_p_O_DFFX1pre_norm_div_(injectionVector[24]),
.p_desc1201_p_O_DFFX1pre_norm_div_(injectionVector[25]),
.p_desc1202_p_O_DFFX1pre_norm_div_(injectionVector[26]),
.p_desc1203_p_O_DFFX1pre_norm_div_(injectionVector[27]),
.p_desc1204_p_O_DFFX1pre_norm_div_(injectionVector[28]),
.p_desc1205_p_O_DFFX1pre_norm_div_(injectionVector[29]),
.p_desc1206_p_O_DFFX1pre_norm_div_(injectionVector[30]),
.p_desc1207_p_O_DFFX1pre_norm_div_(injectionVector[31]),
.p_desc1208_p_O_DFFX1pre_norm_div_(injectionVector[32]),
.p_desc1209_p_O_DFFX1pre_norm_div_(injectionVector[33]),
.p_desc1210_p_O_DFFX1pre_norm_div_(injectionVector[34]),
.p_desc1211_p_O_DFFX1pre_norm_div_(injectionVector[35]),
.p_desc1212_p_O_DFFX1pre_norm_div_(injectionVector[36]),
.p_desc1213_p_O_DFFX1pre_norm_div_(injectionVector[37]),
.p_desc1368_p_O_DFFX1serial_div_(injectionVector[38]),
.p_desc1369_p_O_DFFX1serial_div_(injectionVector[39]),
.p_desc1370_p_O_DFFX1serial_div_(injectionVector[40]),
.p_desc1371_p_O_DFFX1serial_div_(injectionVector[41]),
.p_desc1372_p_O_DFFX1serial_div_(injectionVector[42]),
.p_desc1373_p_O_DFFX1serial_div_(injectionVector[43]),
.p_desc1374_p_O_DFFX1serial_div_(injectionVector[44]),
.p_desc1375_p_O_DFFX1serial_div_(injectionVector[45]),
.p_desc1376_p_O_DFFX1serial_div_(injectionVector[46]),
.p_desc1377_p_O_DFFX1serial_div_(injectionVector[47]),
.p_desc1378_p_O_DFFX1serial_div_(injectionVector[48]),
.p_desc1379_p_O_DFFX1serial_div_(injectionVector[49]),
.p_desc1380_p_O_DFFX1serial_div_(injectionVector[50]),
.p_desc1381_p_O_DFFX1serial_div_(injectionVector[51]),
.p_desc1382_p_O_DFFX1serial_div_(injectionVector[52]),
.p_desc1383_p_O_DFFX1serial_div_(injectionVector[53]),
.p_desc1384_p_O_DFFX1serial_div_(injectionVector[54]),
.p_desc1385_p_O_DFFX1serial_div_(injectionVector[55]),
.p_desc1386_p_O_DFFX1serial_div_(injectionVector[56]),
.p_desc1387_p_O_DFFX1serial_div_(injectionVector[57]),
.p_desc1388_p_O_DFFX1serial_div_(injectionVector[58]),
.p_desc1389_p_O_DFFX1serial_div_(injectionVector[59]),
.p_desc1390_p_O_DFFX1serial_div_(injectionVector[60]),
.p_desc1391_p_O_DFFX1serial_div_(injectionVector[61]),
.p_desc1392_p_O_DFFX1serial_div_(injectionVector[62]),
.p_desc1393_p_O_DFFX1serial_div_(injectionVector[63]),
.p_desc1394_p_O_DFFX1serial_div_(injectionVector[64]),
.p_desc1395_p_O_DFFX1serial_div_(injectionVector[65]),
.p_desc1396_p_O_DFFX1serial_div_(injectionVector[66]),
.p_desc1397_p_O_DFFX1serial_div_(injectionVector[67]),
.p_desc1398_p_O_DFFX1serial_div_(injectionVector[68]),
.p_desc1399_p_O_DFFX1serial_div_(injectionVector[69]),
.p_desc1400_p_O_DFFX1serial_div_(injectionVector[70]),
.p_desc1401_p_O_DFFX1serial_div_(injectionVector[71]),
.p_desc1402_p_O_DFFX1serial_div_(injectionVector[72]),
.p_desc1403_p_O_DFFX1serial_div_(injectionVector[73]),
.p_desc1404_p_O_DFFX1serial_div_(injectionVector[74]),
.p_desc1405_p_O_DFFX1serial_div_(injectionVector[75]),
.p_desc1406_p_O_DFFX1serial_div_(injectionVector[76]),
.p_desc1407_p_O_DFFX1serial_div_(injectionVector[77]),
.p_desc1408_p_O_DFFX1serial_div_(injectionVector[78]),
.p_desc1409_p_O_DFFX1serial_div_(injectionVector[79]),
.p_desc1410_p_O_DFFX1serial_div_(injectionVector[80]),
.p_desc1411_p_O_DFFX1serial_div_(injectionVector[81]),
.p_desc1412_p_O_DFFX1serial_div_(injectionVector[82]),
.p_desc1413_p_O_DFFX1serial_div_(injectionVector[83]),
.p_desc1414_p_O_DFFX1serial_div_(injectionVector[84]),
.p_desc1415_p_O_DFFX1serial_div_(injectionVector[85]),
.p_desc1416_p_O_DFFX1serial_div_(injectionVector[86]),
.p_desc1417_p_O_DFFX1serial_div_(injectionVector[87]),
.p_desc1418_p_O_DFFX1serial_div_(injectionVector[88]),
.p_desc1419_p_O_DFFX1serial_div_(injectionVector[89]),
.p_desc1420_p_O_DFFX1serial_div_(injectionVector[90]),
.p_desc1421_p_O_DFFX1serial_div_(injectionVector[91]),
.p_desc1422_p_O_DFFX1serial_div_(injectionVector[92]),
.p_desc1423_p_O_DFFX1serial_div_(injectionVector[93]),
.p_desc1424_p_O_DFFX1serial_div_(injectionVector[94]),
.p_desc1425_p_O_DFFX1serial_div_(injectionVector[95]),
.p_desc1426_p_O_DFFX1serial_div_(injectionVector[96]),
.p_desc1427_p_O_DFFX1serial_div_(injectionVector[97]),
.p_desc1428_p_O_DFFX1serial_div_(injectionVector[98]),
.p_desc1429_p_O_DFFX1serial_div_(injectionVector[99]),
.p_desc1430_p_O_DFFX1serial_div_(injectionVector[100]),
.p_desc1431_p_O_DFFX1serial_div_(injectionVector[101]),
.p_desc1432_p_O_DFFX1serial_div_(injectionVector[102]),
.p_desc1433_p_O_DFFX1serial_div_(injectionVector[103]),
.p_desc1434_p_O_DFFX1serial_div_(injectionVector[104]),
.p_desc1435_p_O_DFFX1serial_div_(injectionVector[105]),
.p_desc1436_p_O_DFFX1serial_div_(injectionVector[106]),
.p_desc1437_p_O_DFFX1serial_div_(injectionVector[107]),
.p_desc1438_p_O_DFFX1serial_div_(injectionVector[108]),
.p_desc1439_p_O_DFFX1serial_div_(injectionVector[109]),
.p_desc1440_p_O_DFFX1serial_div_(injectionVector[110]),
.p_desc1441_p_O_DFFX1serial_div_(injectionVector[111]),
.p_desc1442_p_O_DFFX1serial_div_(injectionVector[112]),
.p_desc1443_p_O_DFFX1serial_div_(injectionVector[113]),
.p_desc1444_p_O_DFFX1serial_div_(injectionVector[114]),
.p_s_start_i_reg_p_O_DFFX1serial_div_(injectionVector[115]),
.p_s_ready_o_reg_p_O_DFFX1serial_div_(injectionVector[116]),
.p_desc1445_p_O_DFFX1serial_div_(injectionVector[117]),
.p_desc1446_p_O_DFFX1serial_div_(injectionVector[118]),
.p_desc1447_p_O_DFFX1serial_div_(injectionVector[119]),
.p_desc1448_p_O_DFFX1serial_div_(injectionVector[120]),
.p_desc1449_p_O_DFFX1serial_div_(injectionVector[121]),
.p_desc1450_p_O_DFFX1serial_div_(injectionVector[122]),
.p_desc1451_p_O_DFFX1serial_div_(injectionVector[123]),
.p_desc1452_p_O_DFFX1serial_div_(injectionVector[124]),
.p_desc1453_p_O_DFFX1serial_div_(injectionVector[125]),
.p_desc1454_p_O_DFFX1serial_div_(injectionVector[126]),
.p_desc1455_p_O_DFFX1serial_div_(injectionVector[127]),
.p_desc1456_p_O_DFFX1serial_div_(injectionVector[128]),
.p_desc1457_p_O_DFFX1serial_div_(injectionVector[129]),
.p_desc1458_p_O_DFFX1serial_div_(injectionVector[130]),
.p_desc1459_p_O_DFFX1serial_div_(injectionVector[131]),
.p_desc1460_p_O_DFFX1serial_div_(injectionVector[132]),
.p_desc1461_p_O_DFFX1serial_div_(injectionVector[133]),
.p_desc1462_p_O_DFFX1serial_div_(injectionVector[134]),
.p_desc1463_p_O_DFFX1serial_div_(injectionVector[135]),
.p_desc1464_p_O_DFFX1serial_div_(injectionVector[136]),
.p_desc1465_p_O_DFFX1serial_div_(injectionVector[137]),
.p_desc1466_p_O_DFFX1serial_div_(injectionVector[138]),
.p_desc1467_p_O_DFFX1serial_div_(injectionVector[139]),
.p_desc1468_p_O_DFFX1serial_div_(injectionVector[140]),
.p_desc1469_p_O_DFFX1serial_div_(injectionVector[141]),
.p_desc1470_p_O_DFFX1serial_div_(injectionVector[142]),
.p_desc1471_p_O_DFFX1serial_div_(injectionVector[143]),
.p_desc1472_p_O_DFFX1serial_div_(injectionVector[144]),
.p_desc1473_p_O_DFFX1serial_div_(injectionVector[145]),
.p_desc1474_p_O_DFFX1serial_div_(injectionVector[146]),
.p_desc1475_p_O_DFFX1serial_div_(injectionVector[147]),
.p_desc1476_p_O_DFFX1serial_div_(injectionVector[148]),
.p_desc1477_p_O_DFFX1serial_div_(injectionVector[149]),
.p_desc1478_p_O_DFFX1serial_div_(injectionVector[150]),
.p_desc1479_p_O_DFFX1serial_div_(injectionVector[151]),
.p_desc1480_p_O_DFFX1serial_div_(injectionVector[152]),
.p_desc1481_p_O_DFFX1serial_div_(injectionVector[153]),
.p_desc1482_p_O_DFFX1serial_div_(injectionVector[154]),
.p_desc1483_p_O_DFFX1serial_div_(injectionVector[155]),
.p_desc1484_p_O_DFFX1serial_div_(injectionVector[156]),
.p_desc1485_p_O_DFFX1serial_div_(injectionVector[157]),
.p_desc1486_p_O_DFFX1serial_div_(injectionVector[158]),
.p_desc1487_p_O_DFFX1serial_div_(injectionVector[159]),
.p_desc1488_p_O_DFFX1serial_div_(injectionVector[160]),
.p_desc1489_p_O_DFFX1serial_div_(injectionVector[161]),
.p_desc1490_p_O_DFFX1serial_div_(injectionVector[162]),
.p_desc1491_p_O_DFFX1serial_div_(injectionVector[163]),
.p_desc1492_p_O_DFFX1serial_div_(injectionVector[164]),
.p_desc1493_p_O_DFFX1serial_div_(injectionVector[165]),
.p_desc1494_p_O_DFFX1serial_div_(injectionVector[166]),
.p_desc1495_p_O_DFFX1serial_div_(injectionVector[167]),
.p_desc1496_p_O_DFFX1serial_div_(injectionVector[168]),
.p_desc1497_p_O_DFFX1serial_div_(injectionVector[169]),
.p_desc1498_p_O_DFFX1serial_div_(injectionVector[170]),
.p_desc1499_p_O_DFFX1serial_div_(injectionVector[171]),
.p_desc1500_p_O_DFFX1serial_div_(injectionVector[172]),
.p_desc1501_p_O_DFFX1serial_div_(injectionVector[173]),
.p_desc1502_p_O_DFFX1serial_div_(injectionVector[174]),
.p_desc1503_p_O_DFFX1serial_div_(injectionVector[175]),
.p_desc1504_p_O_DFFX1serial_div_(injectionVector[176]),
.p_desc1505_p_O_DFFX1serial_div_(injectionVector[177]),
.p_desc1506_p_O_DFFX1serial_div_(injectionVector[178]),
.p_desc1507_p_O_DFFX1serial_div_(injectionVector[179]),
.p_desc1508_p_O_DFFX1serial_div_(injectionVector[180]),
.p_desc1509_p_O_DFFX1serial_div_(injectionVector[181]),
.p_desc1510_p_O_DFFX1serial_div_(injectionVector[182]),
.p_desc1511_p_O_DFFX1serial_div_(injectionVector[183]),
.p_desc1512_p_O_DFFX1serial_div_(injectionVector[184]),
.p_desc1513_p_O_DFFX1serial_div_(injectionVector[185]),
.p_desc1514_p_O_DFFX1serial_div_(injectionVector[186]),
.p_desc1515_p_O_DFFX1serial_div_(injectionVector[187]),
.p_desc1516_p_O_DFFX1serial_div_(injectionVector[188]),
.p_desc1517_p_O_DFFX1serial_div_(injectionVector[189]),
.p_desc1518_p_O_DFFX1serial_div_(injectionVector[190]),
.p_desc1519_p_O_DFFX1serial_div_(injectionVector[191]),
.p_desc1520_p_O_DFFX1serial_div_(injectionVector[192]),
.p_desc1521_p_O_DFFX1serial_div_(injectionVector[193]),
.p_desc1522_p_O_DFFX1serial_div_(injectionVector[194]),
.p_desc1523_p_O_DFFX1serial_div_(injectionVector[195]),
.p_desc1524_p_O_DFFX1serial_div_(injectionVector[196]),
.p_desc1525_p_O_DFFX1serial_div_(injectionVector[197]),
.p_desc1526_p_O_DFFX1serial_div_(injectionVector[198]),
.p_desc1527_p_O_DFFX1serial_div_(injectionVector[199]),
.p_desc1528_p_O_DFFX1serial_div_(injectionVector[200]),
.p_s_state_reg_p_O_DFFX1serial_div_(injectionVector[201]),
.p_desc1529_p_O_DFFX1serial_div_(injectionVector[202]),
.p_desc1530_p_O_DFFX1post_norm_div_(injectionVector[203]),
.p_desc1531_p_O_DFFX1post_norm_div_(injectionVector[204]),
.p_desc1532_p_O_DFFX1post_norm_div_(injectionVector[205]),
.p_desc1533_p_O_DFFX1post_norm_div_(injectionVector[206]),
.p_desc1534_p_O_DFFX1post_norm_div_(injectionVector[207]),
.p_desc1535_p_O_DFFX1post_norm_div_(injectionVector[208]),
.p_desc1536_p_O_DFFX1post_norm_div_(injectionVector[209]),
.p_desc1537_p_O_DFFX1post_norm_div_(injectionVector[210]),
.p_desc1538_p_O_DFFX1post_norm_div_(injectionVector[211]),
.p_desc1539_p_O_DFFX1post_norm_div_(injectionVector[212]),
.p_desc1540_p_O_DFFX1post_norm_div_(injectionVector[213]),
.p_desc1541_p_O_DFFX1post_norm_div_(injectionVector[214]),
.p_desc1542_p_O_DFFX1post_norm_div_(injectionVector[215]),
.p_desc1543_p_O_DFFX1post_norm_div_(injectionVector[216]),
.p_desc1544_p_O_DFFX1post_norm_div_(injectionVector[217]),
.p_desc1545_p_O_DFFX1post_norm_div_(injectionVector[218]),
.p_desc1546_p_O_DFFX1post_norm_div_(injectionVector[219]),
.p_desc1547_p_O_DFFX1post_norm_div_(injectionVector[220]),
.p_desc1548_p_O_DFFX1post_norm_div_(injectionVector[221]),
.p_desc1549_p_O_DFFX1post_norm_div_(injectionVector[222]),
.p_desc1550_p_O_DFFX1post_norm_div_(injectionVector[223]),
.p_desc1551_p_O_DFFX1post_norm_div_(injectionVector[224]),
.p_desc1552_p_O_DFFX1post_norm_div_(injectionVector[225]),
.p_desc1553_p_O_DFFX1post_norm_div_(injectionVector[226]),
.p_desc1554_p_O_DFFX1post_norm_div_(injectionVector[227]),
.p_desc1555_p_O_DFFX1post_norm_div_(injectionVector[228]),
.p_desc1556_p_O_DFFX1post_norm_div_(injectionVector[229]),
.p_desc1557_p_O_DFFX1post_norm_div_(injectionVector[230]),
.p_desc1558_p_O_DFFX1post_norm_div_(injectionVector[231]),
.p_desc1559_p_O_DFFX1post_norm_div_(injectionVector[232]),
.p_desc1560_p_O_DFFX1post_norm_div_(injectionVector[233]),
.p_desc1561_p_O_DFFX1post_norm_div_(injectionVector[234]),
.p_desc1562_p_O_DFFX1post_norm_div_(injectionVector[235]),
.p_desc1563_p_O_DFFX1post_norm_div_(injectionVector[236]),
.p_desc1564_p_O_DFFX1post_norm_div_(injectionVector[237]),
.p_desc1565_p_O_DFFX1post_norm_div_(injectionVector[238]),
.p_desc1566_p_O_DFFX1post_norm_div_(injectionVector[239]),
.p_desc1567_p_O_DFFX1post_norm_div_(injectionVector[240]),
.p_desc1568_p_O_DFFX1post_norm_div_(injectionVector[241]),
.p_desc1569_p_O_DFFX1post_norm_div_(injectionVector[242]),
.p_desc1570_p_O_DFFX1post_norm_div_(injectionVector[243]),
.p_desc1571_p_O_DFFX1post_norm_div_(injectionVector[244]),
.p_desc1572_p_O_DFFX1post_norm_div_(injectionVector[245]),
.p_desc1573_p_O_DFFX1post_norm_div_(injectionVector[246]),
.p_desc1574_p_O_DFFX1post_norm_div_(injectionVector[247]),
.p_desc1575_p_O_DFFX1post_norm_div_(injectionVector[248]),
.p_desc1576_p_O_DFFX1post_norm_div_(injectionVector[249]),
.p_desc1577_p_O_DFFX1post_norm_div_(injectionVector[250]),
.p_desc1578_p_O_DFFX1post_norm_div_(injectionVector[251]),
.p_desc1579_p_O_DFFX1post_norm_div_(injectionVector[252]),
.p_desc1580_p_O_DFFX1post_norm_div_(injectionVector[253]),
.p_desc1581_p_O_DFFX1post_norm_div_(injectionVector[254]),
.p_desc1582_p_O_DFFX1post_norm_div_(injectionVector[255]),
.p_desc1583_p_O_DFFX1post_norm_div_(injectionVector[256]),
.p_desc1584_p_O_DFFX1post_norm_div_(injectionVector[257]),
.p_desc1585_p_O_DFFX1post_norm_div_(injectionVector[258]),
.p_desc1586_p_O_DFFX1post_norm_div_(injectionVector[259]),
.p_desc1587_p_O_DFFX1post_norm_div_(injectionVector[260]),
.p_desc1588_p_O_DFFX1post_norm_div_(injectionVector[261]),
.p_desc1589_p_O_DFFX1post_norm_div_(injectionVector[262]),
.p_desc1590_p_O_DFFX1post_norm_div_(injectionVector[263]),
.p_desc1591_p_O_DFFX1post_norm_div_(injectionVector[264]),
.p_desc1592_p_O_DFFX1post_norm_div_(injectionVector[265]),
.p_desc1593_p_O_DFFX1post_norm_div_(injectionVector[266]),
.p_desc1594_p_O_DFFX1post_norm_div_(injectionVector[267]),
.p_desc1595_p_O_DFFX1post_norm_div_(injectionVector[268]),
.p_desc1596_p_O_DFFX1post_norm_div_(injectionVector[269]),
.p_desc1597_p_O_DFFX1post_norm_div_(injectionVector[270]),
.p_desc1598_p_O_DFFX1post_norm_div_(injectionVector[271]),
.p_desc1599_p_O_DFFX1post_norm_div_(injectionVector[272]),
.p_desc1600_p_O_DFFX1post_norm_div_(injectionVector[273]),
.p_desc1601_p_O_DFFX1post_norm_div_(injectionVector[274]),
.p_desc1602_p_O_DFFX1post_norm_div_(injectionVector[275]),
.p_desc1603_p_O_DFFX1post_norm_div_(injectionVector[276]),
.p_desc1604_p_O_DFFX1post_norm_div_(injectionVector[277]),
.p_desc1605_p_O_DFFX1post_norm_div_(injectionVector[278]),
.p_desc1606_p_O_DFFX1post_norm_div_(injectionVector[279]),
.p_desc1607_p_O_DFFX1post_norm_div_(injectionVector[280]),
.p_desc1608_p_O_DFFX1post_norm_div_(injectionVector[281]),
.p_desc1609_p_O_DFFX1post_norm_div_(injectionVector[282]),
.p_desc1610_p_O_DFFX1post_norm_div_(injectionVector[283]),
.p_desc1611_p_O_DFFX1post_norm_div_(injectionVector[284]),
.p_desc1612_p_O_DFFX1post_norm_div_(injectionVector[285]),
.p_desc1613_p_O_DFFX1post_norm_div_(injectionVector[286]),
.p_desc1614_p_O_DFFX1post_norm_div_(injectionVector[287]),
.p_desc1615_p_O_DFFX1post_norm_div_(injectionVector[288]),
.p_desc1616_p_O_DFFX1post_norm_div_(injectionVector[289]),
.p_desc1617_p_O_DFFX1post_norm_div_(injectionVector[290]),
.p_desc1618_p_O_DFFX1post_norm_div_(injectionVector[291]),
.p_desc1619_p_O_DFFX1post_norm_div_(injectionVector[292]),
.p_desc1620_p_O_DFFX1post_norm_div_(injectionVector[293]),
.p_desc1621_p_O_DFFX1post_norm_div_(injectionVector[294]),
.p_desc1622_p_O_DFFX1post_norm_div_(injectionVector[295]),
.p_desc1623_p_O_DFFX1post_norm_div_(injectionVector[296]),
.p_desc1624_p_O_DFFX1post_norm_div_(injectionVector[297]),
.p_desc1625_p_O_DFFX1post_norm_div_(injectionVector[298]),
.p_desc1626_p_O_DFFX1post_norm_div_(injectionVector[299]),
.p_desc1627_p_O_DFFX1post_norm_div_(injectionVector[300]),
.p_desc1628_p_O_DFFX1post_norm_div_(injectionVector[301]),
.p_desc1629_p_O_DFFX1post_norm_div_(injectionVector[302]),
.p_desc1630_p_O_DFFX1post_norm_div_(injectionVector[303]),
.p_desc1631_p_O_DFFX1post_norm_div_(injectionVector[304]),
.p_desc1632_p_O_DFFX1post_norm_div_(injectionVector[305]),
.p_desc1633_p_O_DFFX1post_norm_div_(injectionVector[306]),
.p_desc1634_p_O_DFFX1post_norm_div_(injectionVector[307]),
.p_desc1635_p_O_DFFX1post_norm_div_(injectionVector[308]),
.p_desc1636_p_O_DFFX1post_norm_div_(injectionVector[309]),
.p_desc1637_p_O_DFFX1post_norm_div_(injectionVector[310]),
.p_desc1638_p_O_DFFX1post_norm_div_(injectionVector[311]),
.p_desc1639_p_O_DFFX1post_norm_div_(injectionVector[312]),
.p_desc1640_p_O_DFFX1post_norm_div_(injectionVector[313]),
.p_desc1641_p_O_DFFX1post_norm_div_(injectionVector[314]),
.p_desc1642_p_O_DFFX1post_norm_div_(injectionVector[315]),
.p_desc1643_p_O_DFFX1post_norm_div_(injectionVector[316]),
.p_desc1644_p_O_DFFX1post_norm_div_(injectionVector[317]),
.p_desc1645_p_O_DFFX1post_norm_div_(injectionVector[318]),
.p_desc1646_p_O_DFFX1post_norm_div_(injectionVector[319]),
.p_desc1647_p_O_DFFX1post_norm_div_(injectionVector[320]),
.p_desc1648_p_O_DFFX1post_norm_div_(injectionVector[321]),
.p_desc1649_p_O_DFFX1post_norm_div_(injectionVector[322]),
.p_desc1650_p_O_DFFX1post_norm_div_(injectionVector[323]),
.p_desc1651_p_O_DFFX1post_norm_div_(injectionVector[324]),
.p_s_sign_i_reg_p_O_DFFX1post_norm_div_(injectionVector[325]),
.p_desc1652_p_O_DFFX1post_norm_div_(injectionVector[326]),
.p_desc1653_p_O_DFFX1post_norm_div_(injectionVector[327]),
.p_desc1654_p_O_DFFX1post_norm_div_(injectionVector[328]),
.p_desc1658_p_O_DFFX1post_norm_div_(injectionVector[329]),
.p_desc1659_p_O_DFFX1post_norm_div_(injectionVector[330]),
.p_desc1663_p_O_DFFX1post_norm_div_(injectionVector[331]),
.p_desc1664_p_O_DFFX1post_norm_div_(injectionVector[332]),
.p_desc1665_p_O_DFFX1post_norm_div_(injectionVector[333]),
.p_desc1666_p_O_DFFX1post_norm_div_(injectionVector[334]),
.p_desc1667_p_O_DFFX1post_norm_div_(injectionVector[335]),
.p_desc1668_p_O_DFFX1post_norm_div_(injectionVector[336]),
.p_desc1669_p_O_DFFX1post_norm_div_(injectionVector[337]),
.p_desc1670_p_O_DFFX1post_norm_div_(injectionVector[338]),
.p_desc1671_p_O_DFFX1post_norm_div_(injectionVector[339]),
.p_desc1672_p_O_DFFX1post_norm_div_(injectionVector[340]),
.p_desc1673_p_O_DFFX1post_norm_div_(injectionVector[341]),
.p_desc1674_p_O_DFFX1post_norm_div_(injectionVector[342]),
.p_desc1675_p_O_DFFX1post_norm_div_(injectionVector[343]),
.p_desc1676_p_O_DFFX1post_norm_div_(injectionVector[344]),
.p_desc1677_p_O_DFFX1post_norm_div_(injectionVector[345]),
.p_desc1678_p_O_DFFX1post_norm_div_(injectionVector[346]),
.p_desc1679_p_O_DFFX1post_norm_div_(injectionVector[347]),
.p_desc1680_p_O_DFFX1post_norm_div_(injectionVector[348]),
.p_desc1681_p_O_DFFX1post_norm_div_(injectionVector[349]),
.p_desc1682_p_O_DFFX1post_norm_div_(injectionVector[350]),
.p_desc1683_p_O_DFFX1post_norm_div_(injectionVector[351]),
.p_desc1684_p_O_DFFX1post_norm_div_(injectionVector[352]),
.p_desc1685_p_O_DFFX1post_norm_div_(injectionVector[353]),
.p_desc1686_p_O_DFFX1post_norm_div_(injectionVector[354]),
.p_desc1687_p_O_DFFX1post_norm_div_(injectionVector[355]),
.p_desc1688_p_O_DFFX1post_norm_div_(injectionVector[356]),
.p_desc1689_p_O_DFFX1post_norm_div_(injectionVector[357]),
.p_desc1690_p_O_DFFX1post_norm_div_(injectionVector[358]),
.p_desc1691_p_O_DFFX1post_norm_div_(injectionVector[359]),
.p_desc1692_p_O_DFFX1post_norm_div_(injectionVector[360]),
.p_desc1693_p_O_DFFX1post_norm_div_(injectionVector[361]),
.p_desc1694_p_O_DFFX1post_norm_div_(injectionVector[362]),
.p_desc1695_p_O_DFFX1post_norm_div_(injectionVector[363]),
.p_desc1696_p_O_DFFX1post_norm_div_(injectionVector[364]),
.p_desc1697_p_O_DFFX1post_norm_div_(injectionVector[365]),
.p_desc1698_p_O_DFFX1post_norm_div_(injectionVector[366]),
.p_desc1699_p_O_DFFX1post_norm_div_(injectionVector[367]),
.p_desc1700_p_O_DFFX1post_norm_div_(injectionVector[368]),
.p_desc1701_p_O_DFFX1post_norm_div_(injectionVector[369]),
.p_desc1702_p_O_DFFX1post_norm_div_(injectionVector[370]),
.p_desc1703_p_O_DFFX1post_norm_div_(injectionVector[371]),
.p_desc1704_p_O_DFFX1post_norm_div_(injectionVector[372]),
.p_desc1705_p_O_DFFX1post_norm_div_(injectionVector[373]),
.p_desc1706_p_O_DFFX1post_norm_div_(injectionVector[374]),
.p_desc1707_p_O_DFFX1post_norm_div_(injectionVector[375]),
.p_desc1708_p_O_DFFX1post_norm_div_(injectionVector[376]),
.p_desc1709_p_O_DFFX1post_norm_div_(injectionVector[377]),
.p_desc1710_p_O_DFFX1post_norm_div_(injectionVector[378]),
.p_desc1711_p_O_DFFX1post_norm_div_(injectionVector[379]),
.p_desc1712_p_O_DFFX1post_norm_div_(injectionVector[380]),
.p_desc1713_p_O_DFFX1post_norm_div_(injectionVector[381]),
.p_desc1714_p_O_DFFX1post_norm_div_(injectionVector[382]),
.p_desc1715_p_O_DFFX1post_norm_div_(injectionVector[383]),
.p_desc1716_p_O_DFFX1post_norm_div_(injectionVector[384]),
.p_desc1717_p_O_DFFX1post_norm_div_(injectionVector[385]),
.p_desc1718_p_O_DFFX1post_norm_div_(injectionVector[386]),
.p_desc1719_p_O_DFFX1post_norm_div_(injectionVector[387]),
.p_desc1720_p_O_DFFX1post_norm_div_(injectionVector[388]),
.p_desc1721_p_O_DFFX1post_norm_div_(injectionVector[389]),
.p_desc1722_p_O_DFFX1post_norm_div_(injectionVector[390]),
.p_desc1723_p_O_DFFX1post_norm_div_(injectionVector[391]),
.p_desc1724_p_O_DFFX1post_norm_div_(injectionVector[392]),
.p_desc1725_p_O_DFFX1post_norm_div_(injectionVector[393]),
.p_desc1726_p_O_DFFX1post_norm_div_(injectionVector[394]),
.p_desc1727_p_O_DFFX1post_norm_div_(injectionVector[395]),
.p_desc1728_p_O_DFFX1post_norm_div_(injectionVector[396]),
.p_ine_o_reg_p_O_DFFX1post_norm_div_(injectionVector[397]),
.p_desc1729_p_O_DFFX1post_norm_div_(injectionVector[398]),
.p_desc1737_p_O_DFFX1post_norm_div_(injectionVector[399]),
.p_desc1738_p_O_DFFX1post_norm_div_(injectionVector[400]),
.p_desc1739_p_O_DFFX1post_norm_div_(injectionVector[401]),
.p_desc1740_p_O_DFFX1post_norm_div_(injectionVector[402]),
.p_desc1741_p_O_DFFX1post_norm_div_(injectionVector[403]),
.p_desc1742_p_O_DFFX1post_norm_div_(injectionVector[404]),
.p_desc1743_p_O_DFFX1post_norm_div_(injectionVector[405]),
.p_desc1744_p_O_DFFX1post_norm_div_(injectionVector[406]),
.p_desc1745_p_O_DFFX1post_norm_div_(injectionVector[407]),
.p_desc1746_p_O_DFFX1post_norm_div_(injectionVector[408]),
.p_desc1747_p_O_DFFX1post_norm_div_(injectionVector[409]),
.p_desc1748_p_O_DFFX1post_norm_div_(injectionVector[410]),
.p_desc1749_p_O_DFFX1post_norm_div_(injectionVector[411]),
.p_desc1750_p_O_DFFX1post_norm_div_(injectionVector[412]),
.p_desc1751_p_O_DFFX1post_norm_div_(injectionVector[413]),
.p_desc1752_p_O_DFFX1post_norm_div_(injectionVector[414]),
.p_desc1753_p_O_DFFX1post_norm_div_(injectionVector[415]),
.p_desc1754_p_O_DFFX1post_norm_div_(injectionVector[416]),
.p_desc1755_p_O_DFFX1post_norm_div_(injectionVector[417]),
.p_desc1756_p_O_DFFX1post_norm_div_(injectionVector[418]),
.p_desc1757_p_O_DFFX1post_norm_div_(injectionVector[419]),
.p_desc1758_p_O_DFFX1post_norm_div_(injectionVector[420]),
.p_desc1849_p_O_DFFX1post_norm_div_(injectionVector[421]),
.p_desc1850_p_O_DFFX1post_norm_div_(injectionVector[422]),
.p_desc1851_p_O_DFFX1post_norm_div_(injectionVector[423]),
.p_desc1852_p_O_DFFX1post_norm_div_(injectionVector[424]),
.p_desc1853_p_O_DFFX1post_norm_div_(injectionVector[425]),
.p_desc1854_p_O_DFFX1post_norm_div_(injectionVector[426]),
.p_desc1855_p_O_DFFX1post_norm_div_(injectionVector[427]),
.p_desc1856_p_O_DFFX1post_norm_div_(injectionVector[428]),
.p_desc1857_p_O_DFFX1post_norm_div_(injectionVector[429]),
.p_desc1858_p_O_DFFX1post_norm_div_(injectionVector[430]),
.p_desc1859_p_O_DFFX1post_norm_div_(injectionVector[431]),
.p_desc1860_p_O_DFFX1post_norm_div_(injectionVector[432]),
.p_desc1861_p_O_DFFX1post_norm_div_(injectionVector[433]),
.p_desc1862_p_O_DFFX1post_norm_div_(injectionVector[434]),
.p_desc1863_p_O_DFFX1post_norm_div_(injectionVector[435]),
.p_desc1864_p_O_DFFX1post_norm_div_(injectionVector[436]),
.p_desc1865_p_O_DFFX1post_norm_div_(injectionVector[437]),
.p_desc1866_p_O_DFFX1post_norm_div_(injectionVector[438]),
.p_desc1867_p_O_DFFX1post_norm_div_(injectionVector[439]),
.p_desc1868_p_O_DFFX1post_norm_div_(injectionVector[440]),
.p_desc1869_p_O_DFFX1post_norm_div_(injectionVector[441]));
endmodule