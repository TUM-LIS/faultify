`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[68:0] testVector;
output[4:0] resultVector;
input[577:0] injectionVector;
dec_viterbi_inj toplevel_instance (
.aclk(clk),
.aresetn(rst),
.s_axis_input_tvalid(testVector[0]),
.s_axis_input_tdata(testVector [32:1]),
.s_axis_input_tlast(testVector[33]),
.s_axis_input_tready(resultVector[0]),
.m_axis_output_tvalid(resultVector[1]),
.m_axis_output_tdata(resultVector[2]),
.m_axis_output_tlast(resultVector[3]),
.m_axis_output_tready(testVector[34]),
.s_axis_ctrl_tvalid(testVector[35]),
.s_axis_ctrl_tdata(testVector [67:36]),
.s_axis_ctrl_tlast(testVector[68]),
.s_axis_ctrl_tready(resultVector[4]),
.p_output_valid_reg_Z_p_O_FDRaxi4s_buffer_(injectionVector[0]),
.p_m_axis_output_tlast_Z_p_O_FDRbranch_distanceZ0_(injectionVector[1]),
.p_m_axis_output_tvalid_int_Z_p_O_FDRbranch_distanceZ0_(injectionVector[2]),
.p_desc89_p_O_FDRacsZ0_(injectionVector[3]),
.p_desc90_p_O_FDRacsZ0_(injectionVector[4]),
.p_desc91_p_O_FDRacsZ0_(injectionVector[5]),
.p_desc92_p_O_FDRacsZ0_(injectionVector[6]),
.p_desc93_p_O_FDRacsZ0_(injectionVector[7]),
.p_desc94_p_O_FDRacsZ0_(injectionVector[8]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_(injectionVector[9]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_(injectionVector[10]),
.p_desc128_p_O_FDRacsZ0_1_(injectionVector[11]),
.p_desc129_p_O_FDRacsZ0_1_(injectionVector[12]),
.p_desc130_p_O_FDRacsZ0_1_(injectionVector[13]),
.p_desc131_p_O_FDRacsZ0_1_(injectionVector[14]),
.p_desc132_p_O_FDRacsZ0_1_(injectionVector[15]),
.p_desc133_p_O_FDRacsZ0_1_(injectionVector[16]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_1_(injectionVector[17]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_1_(injectionVector[18]),
.p_desc167_p_O_FDRacsZ0_2_(injectionVector[19]),
.p_desc168_p_O_FDRacsZ0_2_(injectionVector[20]),
.p_desc169_p_O_FDRacsZ0_2_(injectionVector[21]),
.p_desc170_p_O_FDRacsZ0_2_(injectionVector[22]),
.p_desc171_p_O_FDRacsZ0_2_(injectionVector[23]),
.p_desc172_p_O_FDRacsZ0_2_(injectionVector[24]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_2_(injectionVector[25]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_2_(injectionVector[26]),
.p_desc206_p_O_FDRacsZ0_3_(injectionVector[27]),
.p_desc207_p_O_FDRacsZ0_3_(injectionVector[28]),
.p_desc208_p_O_FDRacsZ0_3_(injectionVector[29]),
.p_desc209_p_O_FDRacsZ0_3_(injectionVector[30]),
.p_desc210_p_O_FDRacsZ0_3_(injectionVector[31]),
.p_desc211_p_O_FDRacsZ0_3_(injectionVector[32]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_3_(injectionVector[33]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_3_(injectionVector[34]),
.p_desc245_p_O_FDRacsZ0_4_(injectionVector[35]),
.p_desc246_p_O_FDRacsZ0_4_(injectionVector[36]),
.p_desc247_p_O_FDRacsZ0_4_(injectionVector[37]),
.p_desc248_p_O_FDRacsZ0_4_(injectionVector[38]),
.p_desc249_p_O_FDRacsZ0_4_(injectionVector[39]),
.p_desc250_p_O_FDRacsZ0_4_(injectionVector[40]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_4_(injectionVector[41]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_4_(injectionVector[42]),
.p_desc284_p_O_FDRacsZ0_5_(injectionVector[43]),
.p_desc285_p_O_FDRacsZ0_5_(injectionVector[44]),
.p_desc286_p_O_FDRacsZ0_5_(injectionVector[45]),
.p_desc287_p_O_FDRacsZ0_5_(injectionVector[46]),
.p_desc288_p_O_FDRacsZ0_5_(injectionVector[47]),
.p_desc289_p_O_FDRacsZ0_5_(injectionVector[48]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_5_(injectionVector[49]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_5_(injectionVector[50]),
.p_desc323_p_O_FDRacsZ0_6_(injectionVector[51]),
.p_desc324_p_O_FDRacsZ0_6_(injectionVector[52]),
.p_desc325_p_O_FDRacsZ0_6_(injectionVector[53]),
.p_desc326_p_O_FDRacsZ0_6_(injectionVector[54]),
.p_desc327_p_O_FDRacsZ0_6_(injectionVector[55]),
.p_desc328_p_O_FDRacsZ0_6_(injectionVector[56]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_6_(injectionVector[57]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_6_(injectionVector[58]),
.p_desc362_p_O_FDRacsZ0_7_(injectionVector[59]),
.p_desc363_p_O_FDRacsZ0_7_(injectionVector[60]),
.p_desc364_p_O_FDRacsZ0_7_(injectionVector[61]),
.p_desc365_p_O_FDRacsZ0_7_(injectionVector[62]),
.p_desc366_p_O_FDRacsZ0_7_(injectionVector[63]),
.p_desc367_p_O_FDRacsZ0_7_(injectionVector[64]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_7_(injectionVector[65]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_7_(injectionVector[66]),
.p_desc401_p_O_FDRacsZ0_8_(injectionVector[67]),
.p_desc402_p_O_FDRacsZ0_8_(injectionVector[68]),
.p_desc403_p_O_FDRacsZ0_8_(injectionVector[69]),
.p_desc404_p_O_FDRacsZ0_8_(injectionVector[70]),
.p_desc405_p_O_FDRacsZ0_8_(injectionVector[71]),
.p_desc406_p_O_FDRacsZ0_8_(injectionVector[72]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_8_(injectionVector[73]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_8_(injectionVector[74]),
.p_desc440_p_O_FDRacsZ0_9_(injectionVector[75]),
.p_desc441_p_O_FDRacsZ0_9_(injectionVector[76]),
.p_desc442_p_O_FDRacsZ0_9_(injectionVector[77]),
.p_desc443_p_O_FDRacsZ0_9_(injectionVector[78]),
.p_desc444_p_O_FDRacsZ0_9_(injectionVector[79]),
.p_desc445_p_O_FDRacsZ0_9_(injectionVector[80]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_9_(injectionVector[81]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_9_(injectionVector[82]),
.p_desc479_p_O_FDRacsZ0_10_(injectionVector[83]),
.p_desc480_p_O_FDRacsZ0_10_(injectionVector[84]),
.p_desc481_p_O_FDRacsZ0_10_(injectionVector[85]),
.p_desc482_p_O_FDRacsZ0_10_(injectionVector[86]),
.p_desc483_p_O_FDRacsZ0_10_(injectionVector[87]),
.p_desc484_p_O_FDRacsZ0_10_(injectionVector[88]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_10_(injectionVector[89]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_10_(injectionVector[90]),
.p_desc518_p_O_FDRacsZ0_11_(injectionVector[91]),
.p_desc519_p_O_FDRacsZ0_11_(injectionVector[92]),
.p_desc520_p_O_FDRacsZ0_11_(injectionVector[93]),
.p_desc521_p_O_FDRacsZ0_11_(injectionVector[94]),
.p_desc522_p_O_FDRacsZ0_11_(injectionVector[95]),
.p_desc523_p_O_FDRacsZ0_11_(injectionVector[96]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_11_(injectionVector[97]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_11_(injectionVector[98]),
.p_desc557_p_O_FDRacsZ0_12_(injectionVector[99]),
.p_desc558_p_O_FDRacsZ0_12_(injectionVector[100]),
.p_desc559_p_O_FDRacsZ0_12_(injectionVector[101]),
.p_desc560_p_O_FDRacsZ0_12_(injectionVector[102]),
.p_desc561_p_O_FDRacsZ0_12_(injectionVector[103]),
.p_desc562_p_O_FDRacsZ0_12_(injectionVector[104]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_12_(injectionVector[105]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_12_(injectionVector[106]),
.p_desc596_p_O_FDRacsZ0_13_(injectionVector[107]),
.p_desc597_p_O_FDRacsZ0_13_(injectionVector[108]),
.p_desc598_p_O_FDRacsZ0_13_(injectionVector[109]),
.p_desc599_p_O_FDRacsZ0_13_(injectionVector[110]),
.p_desc600_p_O_FDRacsZ0_13_(injectionVector[111]),
.p_desc601_p_O_FDRacsZ0_13_(injectionVector[112]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_13_(injectionVector[113]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_13_(injectionVector[114]),
.p_desc635_p_O_FDRacsZ0_14_(injectionVector[115]),
.p_desc636_p_O_FDRacsZ0_14_(injectionVector[116]),
.p_desc637_p_O_FDRacsZ0_14_(injectionVector[117]),
.p_desc638_p_O_FDRacsZ0_14_(injectionVector[118]),
.p_desc639_p_O_FDRacsZ0_14_(injectionVector[119]),
.p_desc640_p_O_FDRacsZ0_14_(injectionVector[120]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_14_(injectionVector[121]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_14_(injectionVector[122]),
.p_desc674_p_O_FDRacsZ0_15_(injectionVector[123]),
.p_desc675_p_O_FDRacsZ0_15_(injectionVector[124]),
.p_desc676_p_O_FDRacsZ0_15_(injectionVector[125]),
.p_desc677_p_O_FDRacsZ0_15_(injectionVector[126]),
.p_desc678_p_O_FDRacsZ0_15_(injectionVector[127]),
.p_desc679_p_O_FDRacsZ0_15_(injectionVector[128]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_15_(injectionVector[129]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_15_(injectionVector[130]),
.p_desc713_p_O_FDRacsZ0_16_(injectionVector[131]),
.p_desc714_p_O_FDRacsZ0_16_(injectionVector[132]),
.p_desc715_p_O_FDRacsZ0_16_(injectionVector[133]),
.p_desc716_p_O_FDRacsZ0_16_(injectionVector[134]),
.p_desc717_p_O_FDRacsZ0_16_(injectionVector[135]),
.p_desc718_p_O_FDRacsZ0_16_(injectionVector[136]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_16_(injectionVector[137]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_16_(injectionVector[138]),
.p_desc752_p_O_FDRacsZ0_17_(injectionVector[139]),
.p_desc753_p_O_FDRacsZ0_17_(injectionVector[140]),
.p_desc754_p_O_FDRacsZ0_17_(injectionVector[141]),
.p_desc755_p_O_FDRacsZ0_17_(injectionVector[142]),
.p_desc756_p_O_FDRacsZ0_17_(injectionVector[143]),
.p_desc757_p_O_FDRacsZ0_17_(injectionVector[144]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_17_(injectionVector[145]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_17_(injectionVector[146]),
.p_desc791_p_O_FDRacsZ0_18_(injectionVector[147]),
.p_desc792_p_O_FDRacsZ0_18_(injectionVector[148]),
.p_desc793_p_O_FDRacsZ0_18_(injectionVector[149]),
.p_desc794_p_O_FDRacsZ0_18_(injectionVector[150]),
.p_desc795_p_O_FDRacsZ0_18_(injectionVector[151]),
.p_desc796_p_O_FDRacsZ0_18_(injectionVector[152]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_18_(injectionVector[153]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_18_(injectionVector[154]),
.p_desc830_p_O_FDRacsZ0_19_(injectionVector[155]),
.p_desc831_p_O_FDRacsZ0_19_(injectionVector[156]),
.p_desc832_p_O_FDRacsZ0_19_(injectionVector[157]),
.p_desc833_p_O_FDRacsZ0_19_(injectionVector[158]),
.p_desc834_p_O_FDRacsZ0_19_(injectionVector[159]),
.p_desc835_p_O_FDRacsZ0_19_(injectionVector[160]),
.p_desc836_p_O_FDRacsZ0_19_(injectionVector[161]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_19_(injectionVector[162]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_19_(injectionVector[163]),
.p_desc867_p_O_FDRacsZ0_20_(injectionVector[164]),
.p_desc868_p_O_FDRacsZ0_20_(injectionVector[165]),
.p_desc869_p_O_FDRacsZ0_20_(injectionVector[166]),
.p_desc870_p_O_FDRacsZ0_20_(injectionVector[167]),
.p_desc871_p_O_FDRacsZ0_20_(injectionVector[168]),
.p_desc872_p_O_FDRacsZ0_20_(injectionVector[169]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_20_(injectionVector[170]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_20_(injectionVector[171]),
.p_desc906_p_O_FDRacsZ0_21_(injectionVector[172]),
.p_desc907_p_O_FDRacsZ0_21_(injectionVector[173]),
.p_desc908_p_O_FDRacsZ0_21_(injectionVector[174]),
.p_desc909_p_O_FDRacsZ0_21_(injectionVector[175]),
.p_desc910_p_O_FDRacsZ0_21_(injectionVector[176]),
.p_desc911_p_O_FDRacsZ0_21_(injectionVector[177]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_21_(injectionVector[178]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_21_(injectionVector[179]),
.p_desc945_p_O_FDRacsZ1_(injectionVector[180]),
.p_desc946_p_O_FDRacsZ1_(injectionVector[181]),
.p_desc947_p_O_FDRacsZ1_(injectionVector[182]),
.p_desc948_p_O_FDRacsZ1_(injectionVector[183]),
.p_desc949_p_O_FDRacsZ1_(injectionVector[184]),
.p_desc950_p_O_FDRacsZ1_(injectionVector[185]),
.p_desc951_p_O_FDRacsZ1_(injectionVector[186]),
.p_desc952_p_O_FDRacsZ1_(injectionVector[187]),
.p_desc953_p_O_FDRacsZ1_(injectionVector[188]),
.p_m_axis_outdec_tdata_Z_p_O_FDRacsZ1_(injectionVector[189]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ1_(injectionVector[190]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ1_(injectionVector[191]),
.p_m_axis_outdec_tlast_Z_p_O_FDRacsZ1_(injectionVector[192]),
.p_desc983_p_O_FDRacsZ0_22_(injectionVector[193]),
.p_desc984_p_O_FDRacsZ0_22_(injectionVector[194]),
.p_desc985_p_O_FDRacsZ0_22_(injectionVector[195]),
.p_desc986_p_O_FDRacsZ0_22_(injectionVector[196]),
.p_desc987_p_O_FDRacsZ0_22_(injectionVector[197]),
.p_desc988_p_O_FDRacsZ0_22_(injectionVector[198]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_22_(injectionVector[199]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_22_(injectionVector[200]),
.p_desc1022_p_O_FDRacsZ0_23_(injectionVector[201]),
.p_desc1023_p_O_FDRacsZ0_23_(injectionVector[202]),
.p_desc1024_p_O_FDRacsZ0_23_(injectionVector[203]),
.p_desc1025_p_O_FDRacsZ0_23_(injectionVector[204]),
.p_desc1026_p_O_FDRacsZ0_23_(injectionVector[205]),
.p_desc1027_p_O_FDRacsZ0_23_(injectionVector[206]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_23_(injectionVector[207]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_23_(injectionVector[208]),
.p_desc1061_p_O_FDRacsZ0_24_(injectionVector[209]),
.p_desc1062_p_O_FDRacsZ0_24_(injectionVector[210]),
.p_desc1063_p_O_FDRacsZ0_24_(injectionVector[211]),
.p_desc1064_p_O_FDRacsZ0_24_(injectionVector[212]),
.p_desc1065_p_O_FDRacsZ0_24_(injectionVector[213]),
.p_desc1066_p_O_FDRacsZ0_24_(injectionVector[214]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_24_(injectionVector[215]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_24_(injectionVector[216]),
.p_desc1100_p_O_FDRacsZ0_25_(injectionVector[217]),
.p_desc1101_p_O_FDRacsZ0_25_(injectionVector[218]),
.p_desc1102_p_O_FDRacsZ0_25_(injectionVector[219]),
.p_desc1103_p_O_FDRacsZ0_25_(injectionVector[220]),
.p_desc1104_p_O_FDRacsZ0_25_(injectionVector[221]),
.p_desc1105_p_O_FDRacsZ0_25_(injectionVector[222]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_25_(injectionVector[223]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_25_(injectionVector[224]),
.p_desc1139_p_O_FDRacsZ0_26_(injectionVector[225]),
.p_desc1140_p_O_FDRacsZ0_26_(injectionVector[226]),
.p_desc1141_p_O_FDRacsZ0_26_(injectionVector[227]),
.p_desc1142_p_O_FDRacsZ0_26_(injectionVector[228]),
.p_desc1143_p_O_FDRacsZ0_26_(injectionVector[229]),
.p_desc1144_p_O_FDRacsZ0_26_(injectionVector[230]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_26_(injectionVector[231]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_26_(injectionVector[232]),
.p_desc1178_p_O_FDRacsZ0_27_(injectionVector[233]),
.p_desc1179_p_O_FDRacsZ0_27_(injectionVector[234]),
.p_desc1180_p_O_FDRacsZ0_27_(injectionVector[235]),
.p_desc1181_p_O_FDRacsZ0_27_(injectionVector[236]),
.p_desc1182_p_O_FDRacsZ0_27_(injectionVector[237]),
.p_desc1183_p_O_FDRacsZ0_27_(injectionVector[238]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_27_(injectionVector[239]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_27_(injectionVector[240]),
.p_desc1217_p_O_FDRacsZ0_28_(injectionVector[241]),
.p_desc1218_p_O_FDRacsZ0_28_(injectionVector[242]),
.p_desc1219_p_O_FDRacsZ0_28_(injectionVector[243]),
.p_desc1220_p_O_FDRacsZ0_28_(injectionVector[244]),
.p_desc1221_p_O_FDRacsZ0_28_(injectionVector[245]),
.p_desc1222_p_O_FDRacsZ0_28_(injectionVector[246]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_28_(injectionVector[247]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_28_(injectionVector[248]),
.p_desc1256_p_O_FDRacsZ0_29_(injectionVector[249]),
.p_desc1257_p_O_FDRacsZ0_29_(injectionVector[250]),
.p_desc1258_p_O_FDRacsZ0_29_(injectionVector[251]),
.p_desc1259_p_O_FDRacsZ0_29_(injectionVector[252]),
.p_desc1260_p_O_FDRacsZ0_29_(injectionVector[253]),
.p_desc1261_p_O_FDRacsZ0_29_(injectionVector[254]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_29_(injectionVector[255]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_29_(injectionVector[256]),
.p_desc1295_p_O_FDRacsZ0_30_(injectionVector[257]),
.p_desc1296_p_O_FDRacsZ0_30_(injectionVector[258]),
.p_desc1297_p_O_FDRacsZ0_30_(injectionVector[259]),
.p_desc1298_p_O_FDRacsZ0_30_(injectionVector[260]),
.p_desc1299_p_O_FDRacsZ0_30_(injectionVector[261]),
.p_desc1300_p_O_FDRacsZ0_30_(injectionVector[262]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_30_(injectionVector[263]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_30_(injectionVector[264]),
.p_desc1334_p_O_FDRacsZ0_31_(injectionVector[265]),
.p_desc1335_p_O_FDRacsZ0_31_(injectionVector[266]),
.p_desc1336_p_O_FDRacsZ0_31_(injectionVector[267]),
.p_desc1337_p_O_FDRacsZ0_31_(injectionVector[268]),
.p_desc1338_p_O_FDRacsZ0_31_(injectionVector[269]),
.p_desc1339_p_O_FDRacsZ0_31_(injectionVector[270]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_31_(injectionVector[271]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_31_(injectionVector[272]),
.p_desc1373_p_O_FDRacsZ0_32_(injectionVector[273]),
.p_desc1374_p_O_FDRacsZ0_32_(injectionVector[274]),
.p_desc1375_p_O_FDRacsZ0_32_(injectionVector[275]),
.p_desc1376_p_O_FDRacsZ0_32_(injectionVector[276]),
.p_desc1377_p_O_FDRacsZ0_32_(injectionVector[277]),
.p_desc1378_p_O_FDRacsZ0_32_(injectionVector[278]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_32_(injectionVector[279]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_32_(injectionVector[280]),
.p_desc1412_p_O_FDRacsZ0_33_(injectionVector[281]),
.p_desc1413_p_O_FDRacsZ0_33_(injectionVector[282]),
.p_desc1414_p_O_FDRacsZ0_33_(injectionVector[283]),
.p_desc1415_p_O_FDRacsZ0_33_(injectionVector[284]),
.p_desc1416_p_O_FDRacsZ0_33_(injectionVector[285]),
.p_desc1417_p_O_FDRacsZ0_33_(injectionVector[286]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_33_(injectionVector[287]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_33_(injectionVector[288]),
.p_desc1451_p_O_FDRacsZ0_34_(injectionVector[289]),
.p_desc1452_p_O_FDRacsZ0_34_(injectionVector[290]),
.p_desc1453_p_O_FDRacsZ0_34_(injectionVector[291]),
.p_desc1454_p_O_FDRacsZ0_34_(injectionVector[292]),
.p_desc1455_p_O_FDRacsZ0_34_(injectionVector[293]),
.p_desc1456_p_O_FDRacsZ0_34_(injectionVector[294]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_34_(injectionVector[295]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_34_(injectionVector[296]),
.p_desc1490_p_O_FDRacsZ0_35_(injectionVector[297]),
.p_desc1491_p_O_FDRacsZ0_35_(injectionVector[298]),
.p_desc1492_p_O_FDRacsZ0_35_(injectionVector[299]),
.p_desc1493_p_O_FDRacsZ0_35_(injectionVector[300]),
.p_desc1494_p_O_FDRacsZ0_35_(injectionVector[301]),
.p_desc1495_p_O_FDRacsZ0_35_(injectionVector[302]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_35_(injectionVector[303]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_35_(injectionVector[304]),
.p_desc1529_p_O_FDRacsZ0_36_(injectionVector[305]),
.p_desc1530_p_O_FDRacsZ0_36_(injectionVector[306]),
.p_desc1531_p_O_FDRacsZ0_36_(injectionVector[307]),
.p_desc1532_p_O_FDRacsZ0_36_(injectionVector[308]),
.p_desc1533_p_O_FDRacsZ0_36_(injectionVector[309]),
.p_desc1534_p_O_FDRacsZ0_36_(injectionVector[310]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_36_(injectionVector[311]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_36_(injectionVector[312]),
.p_desc1568_p_O_FDRacsZ0_37_(injectionVector[313]),
.p_desc1569_p_O_FDRacsZ0_37_(injectionVector[314]),
.p_desc1570_p_O_FDRacsZ0_37_(injectionVector[315]),
.p_desc1571_p_O_FDRacsZ0_37_(injectionVector[316]),
.p_desc1572_p_O_FDRacsZ0_37_(injectionVector[317]),
.p_desc1573_p_O_FDRacsZ0_37_(injectionVector[318]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_37_(injectionVector[319]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_37_(injectionVector[320]),
.p_desc1607_p_O_FDRacsZ0_38_(injectionVector[321]),
.p_desc1608_p_O_FDRacsZ0_38_(injectionVector[322]),
.p_desc1609_p_O_FDRacsZ0_38_(injectionVector[323]),
.p_desc1610_p_O_FDRacsZ0_38_(injectionVector[324]),
.p_desc1611_p_O_FDRacsZ0_38_(injectionVector[325]),
.p_desc1612_p_O_FDRacsZ0_38_(injectionVector[326]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_38_(injectionVector[327]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_38_(injectionVector[328]),
.p_desc1646_p_O_FDRacsZ0_39_(injectionVector[329]),
.p_desc1647_p_O_FDRacsZ0_39_(injectionVector[330]),
.p_desc1648_p_O_FDRacsZ0_39_(injectionVector[331]),
.p_desc1649_p_O_FDRacsZ0_39_(injectionVector[332]),
.p_desc1650_p_O_FDRacsZ0_39_(injectionVector[333]),
.p_desc1651_p_O_FDRacsZ0_39_(injectionVector[334]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_39_(injectionVector[335]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_39_(injectionVector[336]),
.p_desc1685_p_O_FDRacsZ0_40_(injectionVector[337]),
.p_desc1686_p_O_FDRacsZ0_40_(injectionVector[338]),
.p_desc1687_p_O_FDRacsZ0_40_(injectionVector[339]),
.p_desc1688_p_O_FDRacsZ0_40_(injectionVector[340]),
.p_desc1689_p_O_FDRacsZ0_40_(injectionVector[341]),
.p_desc1690_p_O_FDRacsZ0_40_(injectionVector[342]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_40_(injectionVector[343]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_40_(injectionVector[344]),
.p_desc1724_p_O_FDRacsZ0_41_(injectionVector[345]),
.p_desc1725_p_O_FDRacsZ0_41_(injectionVector[346]),
.p_desc1726_p_O_FDRacsZ0_41_(injectionVector[347]),
.p_desc1727_p_O_FDRacsZ0_41_(injectionVector[348]),
.p_desc1728_p_O_FDRacsZ0_41_(injectionVector[349]),
.p_desc1729_p_O_FDRacsZ0_41_(injectionVector[350]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_41_(injectionVector[351]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_41_(injectionVector[352]),
.p_desc1763_p_O_FDRacsZ0_42_(injectionVector[353]),
.p_desc1764_p_O_FDRacsZ0_42_(injectionVector[354]),
.p_desc1765_p_O_FDRacsZ0_42_(injectionVector[355]),
.p_desc1766_p_O_FDRacsZ0_42_(injectionVector[356]),
.p_desc1767_p_O_FDRacsZ0_42_(injectionVector[357]),
.p_desc1768_p_O_FDRacsZ0_42_(injectionVector[358]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_42_(injectionVector[359]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_42_(injectionVector[360]),
.p_desc1802_p_O_FDRacsZ0_43_(injectionVector[361]),
.p_desc1803_p_O_FDRacsZ0_43_(injectionVector[362]),
.p_desc1804_p_O_FDRacsZ0_43_(injectionVector[363]),
.p_desc1805_p_O_FDRacsZ0_43_(injectionVector[364]),
.p_desc1806_p_O_FDRacsZ0_43_(injectionVector[365]),
.p_desc1807_p_O_FDRacsZ0_43_(injectionVector[366]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_43_(injectionVector[367]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_43_(injectionVector[368]),
.p_desc1841_p_O_FDRacsZ0_44_(injectionVector[369]),
.p_desc1842_p_O_FDRacsZ0_44_(injectionVector[370]),
.p_desc1843_p_O_FDRacsZ0_44_(injectionVector[371]),
.p_desc1844_p_O_FDRacsZ0_44_(injectionVector[372]),
.p_desc1845_p_O_FDRacsZ0_44_(injectionVector[373]),
.p_desc1846_p_O_FDRacsZ0_44_(injectionVector[374]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_44_(injectionVector[375]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_44_(injectionVector[376]),
.p_desc1880_p_O_FDRacsZ0_45_(injectionVector[377]),
.p_desc1881_p_O_FDRacsZ0_45_(injectionVector[378]),
.p_desc1882_p_O_FDRacsZ0_45_(injectionVector[379]),
.p_desc1883_p_O_FDRacsZ0_45_(injectionVector[380]),
.p_desc1884_p_O_FDRacsZ0_45_(injectionVector[381]),
.p_desc1885_p_O_FDRacsZ0_45_(injectionVector[382]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_45_(injectionVector[383]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_45_(injectionVector[384]),
.p_desc1919_p_O_FDRacsZ0_46_(injectionVector[385]),
.p_desc1920_p_O_FDRacsZ0_46_(injectionVector[386]),
.p_desc1921_p_O_FDRacsZ0_46_(injectionVector[387]),
.p_desc1922_p_O_FDRacsZ0_46_(injectionVector[388]),
.p_desc1923_p_O_FDRacsZ0_46_(injectionVector[389]),
.p_desc1924_p_O_FDRacsZ0_46_(injectionVector[390]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_46_(injectionVector[391]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_46_(injectionVector[392]),
.p_desc1958_p_O_FDRacsZ0_47_(injectionVector[393]),
.p_desc1959_p_O_FDRacsZ0_47_(injectionVector[394]),
.p_desc1960_p_O_FDRacsZ0_47_(injectionVector[395]),
.p_desc1961_p_O_FDRacsZ0_47_(injectionVector[396]),
.p_desc1962_p_O_FDRacsZ0_47_(injectionVector[397]),
.p_desc1963_p_O_FDRacsZ0_47_(injectionVector[398]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_47_(injectionVector[399]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_47_(injectionVector[400]),
.p_desc1997_p_O_FDRacsZ0_48_(injectionVector[401]),
.p_desc1998_p_O_FDRacsZ0_48_(injectionVector[402]),
.p_desc1999_p_O_FDRacsZ0_48_(injectionVector[403]),
.p_desc2000_p_O_FDRacsZ0_48_(injectionVector[404]),
.p_desc2001_p_O_FDRacsZ0_48_(injectionVector[405]),
.p_desc2002_p_O_FDRacsZ0_48_(injectionVector[406]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_48_(injectionVector[407]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_48_(injectionVector[408]),
.p_desc2036_p_O_FDRacsZ0_49_(injectionVector[409]),
.p_desc2037_p_O_FDRacsZ0_49_(injectionVector[410]),
.p_desc2038_p_O_FDRacsZ0_49_(injectionVector[411]),
.p_desc2039_p_O_FDRacsZ0_49_(injectionVector[412]),
.p_desc2040_p_O_FDRacsZ0_49_(injectionVector[413]),
.p_desc2041_p_O_FDRacsZ0_49_(injectionVector[414]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_49_(injectionVector[415]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_49_(injectionVector[416]),
.p_desc2075_p_O_FDRacsZ0_50_(injectionVector[417]),
.p_desc2076_p_O_FDRacsZ0_50_(injectionVector[418]),
.p_desc2077_p_O_FDRacsZ0_50_(injectionVector[419]),
.p_desc2078_p_O_FDRacsZ0_50_(injectionVector[420]),
.p_desc2079_p_O_FDRacsZ0_50_(injectionVector[421]),
.p_desc2080_p_O_FDRacsZ0_50_(injectionVector[422]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_50_(injectionVector[423]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_50_(injectionVector[424]),
.p_desc2114_p_O_FDRacsZ0_51_(injectionVector[425]),
.p_desc2115_p_O_FDRacsZ0_51_(injectionVector[426]),
.p_desc2116_p_O_FDRacsZ0_51_(injectionVector[427]),
.p_desc2117_p_O_FDRacsZ0_51_(injectionVector[428]),
.p_desc2118_p_O_FDRacsZ0_51_(injectionVector[429]),
.p_desc2119_p_O_FDRacsZ0_51_(injectionVector[430]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_51_(injectionVector[431]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_51_(injectionVector[432]),
.p_desc2153_p_O_FDRacsZ0_52_(injectionVector[433]),
.p_desc2154_p_O_FDRacsZ0_52_(injectionVector[434]),
.p_desc2155_p_O_FDRacsZ0_52_(injectionVector[435]),
.p_desc2156_p_O_FDRacsZ0_52_(injectionVector[436]),
.p_desc2157_p_O_FDRacsZ0_52_(injectionVector[437]),
.p_desc2158_p_O_FDRacsZ0_52_(injectionVector[438]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_52_(injectionVector[439]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_52_(injectionVector[440]),
.p_desc2192_p_O_FDRacsZ0_53_(injectionVector[441]),
.p_desc2193_p_O_FDRacsZ0_53_(injectionVector[442]),
.p_desc2194_p_O_FDRacsZ0_53_(injectionVector[443]),
.p_desc2195_p_O_FDRacsZ0_53_(injectionVector[444]),
.p_desc2196_p_O_FDRacsZ0_53_(injectionVector[445]),
.p_desc2197_p_O_FDRacsZ0_53_(injectionVector[446]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_53_(injectionVector[447]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_53_(injectionVector[448]),
.p_desc2231_p_O_FDRacsZ0_54_(injectionVector[449]),
.p_desc2232_p_O_FDRacsZ0_54_(injectionVector[450]),
.p_desc2233_p_O_FDRacsZ0_54_(injectionVector[451]),
.p_desc2234_p_O_FDRacsZ0_54_(injectionVector[452]),
.p_desc2235_p_O_FDRacsZ0_54_(injectionVector[453]),
.p_desc2236_p_O_FDRacsZ0_54_(injectionVector[454]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_54_(injectionVector[455]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_54_(injectionVector[456]),
.p_desc2270_p_O_FDRacsZ0_55_(injectionVector[457]),
.p_desc2271_p_O_FDRacsZ0_55_(injectionVector[458]),
.p_desc2272_p_O_FDRacsZ0_55_(injectionVector[459]),
.p_desc2273_p_O_FDRacsZ0_55_(injectionVector[460]),
.p_desc2274_p_O_FDRacsZ0_55_(injectionVector[461]),
.p_desc2275_p_O_FDRacsZ0_55_(injectionVector[462]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_55_(injectionVector[463]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_55_(injectionVector[464]),
.p_desc2309_p_O_FDRacsZ0_56_(injectionVector[465]),
.p_desc2310_p_O_FDRacsZ0_56_(injectionVector[466]),
.p_desc2311_p_O_FDRacsZ0_56_(injectionVector[467]),
.p_desc2312_p_O_FDRacsZ0_56_(injectionVector[468]),
.p_desc2313_p_O_FDRacsZ0_56_(injectionVector[469]),
.p_desc2314_p_O_FDRacsZ0_56_(injectionVector[470]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_56_(injectionVector[471]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_56_(injectionVector[472]),
.p_desc2348_p_O_FDRacsZ0_57_(injectionVector[473]),
.p_desc2349_p_O_FDRacsZ0_57_(injectionVector[474]),
.p_desc2350_p_O_FDRacsZ0_57_(injectionVector[475]),
.p_desc2351_p_O_FDRacsZ0_57_(injectionVector[476]),
.p_desc2352_p_O_FDRacsZ0_57_(injectionVector[477]),
.p_desc2353_p_O_FDRacsZ0_57_(injectionVector[478]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_57_(injectionVector[479]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_57_(injectionVector[480]),
.p_desc2387_p_O_FDRacsZ0_58_(injectionVector[481]),
.p_desc2388_p_O_FDRacsZ0_58_(injectionVector[482]),
.p_desc2389_p_O_FDRacsZ0_58_(injectionVector[483]),
.p_desc2390_p_O_FDRacsZ0_58_(injectionVector[484]),
.p_desc2391_p_O_FDRacsZ0_58_(injectionVector[485]),
.p_desc2392_p_O_FDRacsZ0_58_(injectionVector[486]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_58_(injectionVector[487]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_58_(injectionVector[488]),
.p_desc2426_p_O_FDRacsZ0_59_(injectionVector[489]),
.p_desc2427_p_O_FDRacsZ0_59_(injectionVector[490]),
.p_desc2428_p_O_FDRacsZ0_59_(injectionVector[491]),
.p_desc2429_p_O_FDRacsZ0_59_(injectionVector[492]),
.p_desc2430_p_O_FDRacsZ0_59_(injectionVector[493]),
.p_desc2431_p_O_FDRacsZ0_59_(injectionVector[494]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_59_(injectionVector[495]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_59_(injectionVector[496]),
.p_desc2465_p_O_FDRacsZ0_60_(injectionVector[497]),
.p_desc2466_p_O_FDRacsZ0_60_(injectionVector[498]),
.p_desc2467_p_O_FDRacsZ0_60_(injectionVector[499]),
.p_desc2468_p_O_FDRacsZ0_60_(injectionVector[500]),
.p_desc2469_p_O_FDRacsZ0_60_(injectionVector[501]),
.p_desc2470_p_O_FDRacsZ0_60_(injectionVector[502]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_60_(injectionVector[503]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_60_(injectionVector[504]),
.p_desc2504_p_O_FDRacsZ0_61_(injectionVector[505]),
.p_desc2505_p_O_FDRacsZ0_61_(injectionVector[506]),
.p_desc2506_p_O_FDRacsZ0_61_(injectionVector[507]),
.p_desc2507_p_O_FDRacsZ0_61_(injectionVector[508]),
.p_desc2508_p_O_FDRacsZ0_61_(injectionVector[509]),
.p_desc2509_p_O_FDRacsZ0_61_(injectionVector[510]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_61_(injectionVector[511]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_61_(injectionVector[512]),
.p_desc2543_p_O_FDRacsZ0_62_(injectionVector[513]),
.p_desc2544_p_O_FDRacsZ0_62_(injectionVector[514]),
.p_desc2545_p_O_FDRacsZ0_62_(injectionVector[515]),
.p_desc2546_p_O_FDRacsZ0_62_(injectionVector[516]),
.p_desc2547_p_O_FDRacsZ0_62_(injectionVector[517]),
.p_desc2548_p_O_FDRacsZ0_62_(injectionVector[518]),
.p_s_axis_inbranch_tlast_d_Z_p_O_FDRacsZ0_62_(injectionVector[519]),
.p_m_axis_outdec_tvalid_int_Z_p_O_FDRacsZ0_62_(injectionVector[520]),
.p_desc2587_p_O_FDRram_ctrl_(injectionVector[521]),
.p_desc2588_p_O_FDRram_ctrl_(injectionVector[522]),
.p_desc2589_p_O_FDRram_ctrl_(injectionVector[523]),
.p_desc2590_p_O_FDRram_ctrl_(injectionVector[524]),
.p_desc2616_p_O_FDRram_ctrl_(injectionVector[525]),
.p_desc2617_p_O_FDRram_ctrl_(injectionVector[526]),
.p_desc2618_p_O_FDRram_ctrl_(injectionVector[527]),
.p_desc2619_p_O_FDRram_ctrl_(injectionVector[528]),
.p_write_window_complete_Z_p_O_FDRram_ctrl_(injectionVector[529]),
.p_write_last_window_complete_Z_p_O_FDRram_ctrl_(injectionVector[530]),
.p_last_of_block_Z_p_O_FDRram_ctrl_(injectionVector[531]),
.p_desc2659_p_O_FDRram_ctrl_(injectionVector[532]),
.p_desc2660_p_O_FDRram_ctrl_(injectionVector[533]),
.p_desc2661_p_O_FDRram_ctrl_(injectionVector[534]),
.p_desc2662_p_O_FDRram_ctrl_(injectionVector[535]),
.p_desc2663_p_O_FDRram_ctrl_(injectionVector[536]),
.p_desc2664_p_O_FDRram_ctrl_(injectionVector[537]),
.p_desc2665_p_O_FDRram_ctrl_(injectionVector[538]),
.p_desc2966_p_O_FDRram_ctrl_(injectionVector[539]),
.p_desc2967_p_O_FDRram_ctrl_(injectionVector[540]),
.p_desc2968_p_O_FDRram_ctrl_(injectionVector[541]),
.p_desc2969_p_O_FDRram_ctrl_(injectionVector[542]),
.p_desc3139_p_O_FDRram_ctrl_(injectionVector[543]),
.p_desc3140_p_O_FDRram_ctrl_(injectionVector[544]),
.p_desc3141_p_O_FDRram_ctrl_(injectionVector[545]),
.p_desc3142_p_O_FDRram_ctrl_(injectionVector[546]),
.p_m_axis_output_tdata_Z_p_O_FDRtrellis_traceback_(injectionVector[547]),
.p_m_axis_output_tvalid_int_Z_p_O_FDRtrellis_traceback_(injectionVector[548]),
.p_m_axis_output_tdata_Z_p_O_FDRtrellis_traceback_1_(injectionVector[549]),
.p_m_axis_output_tvalid_int_Z_p_O_FDRtrellis_traceback_1_(injectionVector[550]),
.p_send_output_Z_p_O_FDRreorder_(injectionVector[551]),
.p_m_axis_output_last_tuser_Z_p_O_FDRreorder_(injectionVector[552]),
.p_last_window_Z_p_O_FDRreorder_(injectionVector[553]),
.p_send_output_fast_Z_p_O_FDRreorder_(injectionVector[554]),
.p_send_output_rep1_Z_p_O_FDRreorder_(injectionVector[555]),
.p_send_output_rep2_Z_p_O_FDRreorder_(injectionVector[556]),
.p_desc3400_p_O_FDRreorder_(injectionVector[557]),
.p_desc3401_p_O_FDRreorder_(injectionVector[558]),
.p_desc3402_p_O_FDRreorder_(injectionVector[559]),
.p_desc3403_p_O_FDRreorder_(injectionVector[560]),
.p_desc3404_p_O_FDRreorder_(injectionVector[561]),
.p_desc3405_p_O_FDRreorder_(injectionVector[562]),
.p_desc3406_p_O_FDRreorder_(injectionVector[563]),
.p_send_output_Z_p_O_FDRreorder_1_(injectionVector[564]),
.p_m_axis_output_last_tuser_Z_p_O_FDRreorder_1_(injectionVector[565]),
.p_last_window_Z_p_O_FDRreorder_1_(injectionVector[566]),
.p_send_output_fast_Z_p_O_FDRreorder_1_(injectionVector[567]),
.p_send_output_rep1_Z_p_O_FDRreorder_1_(injectionVector[568]),
.p_send_output_rep2_Z_p_O_FDRreorder_1_(injectionVector[569]),
.p_desc3605_p_O_FDRreorder_1_(injectionVector[570]),
.p_desc3606_p_O_FDRreorder_1_(injectionVector[571]),
.p_desc3607_p_O_FDRreorder_1_(injectionVector[572]),
.p_desc3608_p_O_FDRreorder_1_(injectionVector[573]),
.p_desc3609_p_O_FDRreorder_1_(injectionVector[574]),
.p_desc3610_p_O_FDRreorder_1_(injectionVector[575]),
.p_desc3611_p_O_FDRreorder_1_(injectionVector[576]),
.p_desc3706_p_O_FDR(injectionVector[577]));
endmodule