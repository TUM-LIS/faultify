module axi4s_buffer_inj (buffer_tdata_i,acs_tvalid,write_ram_fsm,s_axis_input_tdata_0,s_axis_input_tdata_1,s_axis_input_tdata_2,s_axis_input_tdata_3,s_axis_input_tdata_8,s_axis_input_tdata_9,s_axis_input_tdata_10,s_axis_input_tdata_11,buffer_tdata_3,buffer_tdata_2,buffer_tdata_1,buffer_tdata_10,buffer_tdata_9,buffer_tdata_11,buffer_tdata_8,buffer_tdata_0,s_axis_input_tready,aclk,aresetn_i,buffer_tvalid,un27_s_axis_input_tready_int,write_ram_fsm_0_rep1,write_ram_fsm_4_rep1,N_1756_1,s_axis_input_tvalid,s_axis_input_tlast,N_2388_i,buffer_tlast);
output [3:1] buffer_tdata_i ;
input acs_tvalid ;
input [1:1] write_ram_fsm ;
input s_axis_input_tdata_0 ;
input s_axis_input_tdata_1 ;
input s_axis_input_tdata_2 ;
input s_axis_input_tdata_3 ;
input s_axis_input_tdata_8 ;
input s_axis_input_tdata_9 ;
input s_axis_input_tdata_10 ;
input s_axis_input_tdata_11 ;
output buffer_tdata_3 ;
output buffer_tdata_2 ;
output buffer_tdata_1 ;
output buffer_tdata_10 ;
output buffer_tdata_9 ;
output buffer_tdata_11 ;
output buffer_tdata_8 ;
output buffer_tdata_0 ;
output s_axis_input_tready ;
input aclk ;
input aresetn_i ;
output buffer_tvalid ;
input un27_s_axis_input_tready_int ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input s_axis_input_tvalid ;
input s_axis_input_tlast ;
output N_2388_i ;
output buffer_tlast ;
wire s_axis_input_tdata_0 ;
wire s_axis_input_tdata_1 ;
wire s_axis_input_tdata_2 ;
wire s_axis_input_tdata_3 ;
wire s_axis_input_tdata_8 ;
wire s_axis_input_tdata_9 ;
wire s_axis_input_tdata_10 ;
wire s_axis_input_tdata_11 ;
wire buffer_tdata_3 ;
wire buffer_tdata_2 ;
wire buffer_tdata_1 ;
wire buffer_tdata_10 ;
wire buffer_tdata_9 ;
wire buffer_tdata_11 ;
wire buffer_tdata_8 ;
wire buffer_tdata_0 ;
wire s_axis_input_tready ;
wire aclk ;
wire aresetn_i ;
wire buffer_tvalid ;
wire un27_s_axis_input_tready_int ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire s_axis_input_tvalid ;
wire s_axis_input_tlast ;
wire N_2388_i ;
wire buffer_tlast ;
wire [11:0] buffer_data ;
wire [11:0] output_reg_4 ;
wire un3_output_accept_0 ;
wire buffer_full ;
wire buffer_full_1_sqmuxa_i ;
wire un5_input_valid_1_i ;
wire un5_input_valid ;
wire output_valid_reg_RNO ;
wire buffer_last ;
wire output_last_reg_4 ;
wire N_1106 ;
wire N_1105 ;
wire N_1104 ;
wire N_1103 ;
wire N_1102 ;
wire N_1101 ;
wire N_1100 ;
wire N_1099 ;
wire N_1098 ;
wire N_1097 ;
wire N_1096 ;
wire N_1095 ;
wire N_1094 ;
wire N_1093 ;
wire N_1092 ;
wire N_1091 ;
wire N_1090 ;
wire N_1089 ;
wire N_1088 ;
wire N_1087 ;
wire N_1086 ;
wire N_1085 ;
wire N_1084 ;
wire N_1083 ;
wire N_1082 ;
wire N_1081 ;
wire N_1080 ;
wire N_1079 ;
wire N_1078 ;
wire N_1077 ;
wire N_1076 ;
wire N_1075 ;
wire N_1074 ;
wire N_1073 ;
wire N_1072 ;
wire N_1071 ;
wire N_1070 ;
wire N_1069 ;
wire N_1068 ;
wire N_1067 ;
wire N_1066 ;
wire N_1065 ;
wire N_1064 ;
wire N_1063 ;
wire N_1062 ;
wire N_1061 ;
wire N_1060 ;
wire N_1059 ;
wire GND ;
wire VCC ;
// instances
  LUT1 desc0(.I0(buffer_tdata_3),.O(buffer_tdata_i[3:3]));
defparam desc0.INIT=2'h1;
  LUT1 desc1(.I0(buffer_tdata_2),.O(buffer_tdata_i[2:2]));
defparam desc1.INIT=2'h1;
  LUT1 desc2(.I0(buffer_tdata_1),.O(buffer_tdata_i[1:1]));
defparam desc2.INIT=2'h1;
  FDS input_accept_int_Z(.Q(s_axis_input_tready),.D(un3_output_accept_0),.C(aclk),.S(aresetn_i));
  LUT6 desc3(.I0(buffer_full),.I1(buffer_tvalid),.I2(acs_tvalid),.I3(un27_s_axis_input_tready_int),.I4(s_axis_input_tready),.I5(buffer_full_1_sqmuxa_i),.O(un3_output_accept_0));
defparam desc3.INIT=64'h08880888FFFF0000;
  LUT6 output_valid_reg_RNIA2NP4(.I0(write_ram_fsm_0_rep1),.I1(buffer_tvalid),.I2(write_ram_fsm_4_rep1),.I3(acs_tvalid),.I4(write_ram_fsm[1:1]),.I5(N_1756_1),.O(un5_input_valid_1_i));
defparam output_valid_reg_RNIA2NP4.INIT=64'h33FF37FF33FF33FF;
  LUT5 desc4(.I0(s_axis_input_tvalid),.I1(s_axis_input_tready),.I2(buffer_tvalid),.I3(acs_tvalid),.I4(un27_s_axis_input_tready_int),.O(un5_input_valid));
defparam desc4.INIT=32'h80000000;
  LUT5_L output_valid_reg_RNO_cZ(.I0(s_axis_input_tvalid),.I1(buffer_full),.I2(buffer_tvalid),.I3(acs_tvalid),.I4(un27_s_axis_input_tready_int),.LO(output_valid_reg_RNO));
defparam output_valid_reg_RNO_cZ.INIT=32'hFAEAEAEA;
  LUT6_L desc5(.I0(s_axis_input_tlast),.I1(buffer_last),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_last_reg_4));
defparam desc5.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc6(.I0(s_axis_input_tdata_0),.I1(buffer_data[0:0]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[0:0]));
defparam desc6.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc7(.I0(s_axis_input_tdata_1),.I1(buffer_data[1:1]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[1:1]));
defparam desc7.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc8(.I0(s_axis_input_tdata_2),.I1(buffer_data[2:2]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[2:2]));
defparam desc8.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc9(.I0(s_axis_input_tdata_3),.I1(buffer_data[3:3]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[3:3]));
defparam desc9.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc10(.I0(s_axis_input_tdata_8),.I1(buffer_data[8:8]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[8:8]));
defparam desc10.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc11(.I0(s_axis_input_tdata_9),.I1(buffer_data[9:9]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[9:9]));
defparam desc11.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc12(.I0(s_axis_input_tdata_10),.I1(buffer_data[10:10]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[10:10]));
defparam desc12.INIT=64'hAAAACAAACAAACAAA;
  LUT6_L desc13(.I0(s_axis_input_tdata_11),.I1(buffer_data[11:11]),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.LO(output_reg_4[11:11]));
defparam desc13.INIT=64'hAAAACAAACAAACAAA;
  LUT6 buffer_full_1_sqmuxa_i_cZ(.I0(s_axis_input_tvalid),.I1(s_axis_input_tready),.I2(buffer_full),.I3(buffer_tvalid),.I4(acs_tvalid),.I5(un27_s_axis_input_tready_int),.O(buffer_full_1_sqmuxa_i));
defparam buffer_full_1_sqmuxa_i_cZ.INIT=64'h8800F000F000F000;
  LUT4 desc14(.I0(buffer_tdata_10),.I1(buffer_tdata_9),.I2(buffer_tdata_11),.I3(buffer_tdata_8),.O(N_2388_i));
defparam desc14.INIT=16'h0F0E;
  FDR output_valid_reg_Z(.Q(buffer_tvalid),.D(output_valid_reg_RNO),.C(aclk),.R(aresetn_i));
  FDRE buffer_last_Z(.Q(buffer_last),.D(s_axis_input_tlast),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc15(.Q(buffer_data[11:11]),.D(s_axis_input_tdata_11),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc16(.Q(buffer_data[10:10]),.D(s_axis_input_tdata_10),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc17(.Q(buffer_data[9:9]),.D(s_axis_input_tdata_9),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc18(.Q(buffer_data[8:8]),.D(s_axis_input_tdata_8),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc19(.Q(buffer_data[3:3]),.D(s_axis_input_tdata_3),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc20(.Q(buffer_data[2:2]),.D(s_axis_input_tdata_2),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc21(.Q(buffer_data[1:1]),.D(s_axis_input_tdata_1),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE desc22(.Q(buffer_data[0:0]),.D(s_axis_input_tdata_0),.C(aclk),.R(aresetn_i),.CE(un5_input_valid));
  FDRE output_last_reg_Z(.Q(buffer_tlast),.D(output_last_reg_4),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc23(.Q(buffer_tdata_11),.D(output_reg_4[11:11]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc24(.Q(buffer_tdata_10),.D(output_reg_4[10:10]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc25(.Q(buffer_tdata_9),.D(output_reg_4[9:9]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc26(.Q(buffer_tdata_8),.D(output_reg_4[8:8]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc27(.Q(buffer_tdata_3),.D(output_reg_4[3:3]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc28(.Q(buffer_tdata_2),.D(output_reg_4[2:2]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc29(.Q(buffer_tdata_1),.D(output_reg_4[1:1]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE desc30(.Q(buffer_tdata_0),.D(output_reg_4[0:0]),.C(aclk),.R(aresetn_i),.CE(un5_input_valid_1_i));
  FDRE buffer_full_Z(.Q(buffer_full),.D(un5_input_valid),.C(aclk),.R(aresetn_i),.CE(buffer_full_1_sqmuxa_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module branch_distanceZ3_inj (branch_tdata_3_fast,buffer_tdata_0,buffer_tdata_8,buffer_tdata_1,buffer_tdata_9,buffer_tdata_10,buffer_tdata_11,buffer_tdata_3,buffer_tdata_2,buffer_tdata_i,branch_tdata_3,branch_tdata_3_0_rep2,aclk,aresetn_i,un1_output_accept,branch_tdata_3_0_rep1,N_2388_i,p_m_axis_output_tdata_0_rep2_Z_p_O_FDRE,p_m_axis_output_tdata_0_rep1_Z_p_O_FDRE,p_desc31_p_O_FDRE,p_desc32_p_O_FDRE,p_desc33_p_O_FDRE,p_desc34_p_O_FDRE,p_desc35_p_O_FDRE,p_desc36_p_O_FDRE,p_desc37_p_O_FDRE);
output branch_tdata_3_fast ;
input buffer_tdata_0 ;
input buffer_tdata_8 ;
input buffer_tdata_1 ;
input buffer_tdata_9 ;
input buffer_tdata_10 ;
input buffer_tdata_11 ;
input buffer_tdata_3 ;
input buffer_tdata_2 ;
input [3:1] buffer_tdata_i ;
output [5:0] branch_tdata_3 ;
output branch_tdata_3_0_rep2 ;
input aclk ;
input aresetn_i ;
input un1_output_accept ;
output branch_tdata_3_0_rep1 ;
input N_2388_i ;
wire buffer_tdata_0 ;
wire buffer_tdata_8 ;
wire buffer_tdata_1 ;
wire buffer_tdata_9 ;
wire buffer_tdata_10 ;
wire buffer_tdata_11 ;
wire buffer_tdata_3 ;
wire buffer_tdata_2 ;
wire branch_tdata_3_0_rep2 ;
wire aclk ;
wire aresetn_i ;
wire un1_output_accept ;
wire branch_tdata_3_0_rep1 ;
wire N_2388_i ;
wire [5:1] v_branch_result_3 ;
wire GND ;
wire VCC ;
wire v_branch_result_3_axb_0_i ;
wire v_branch_result_3_axb_0_i_rep1 ;
wire v_branch_result_3_axb_0_i_fast ;
wire v_branch_result_3_axb_0_i_rep2 ;
wire v_branch_result_3_axb_0 ;
wire v_branch_result_3_axb_1 ;
wire v_branch_result_3_axb_5 ;
wire v_branch_result_3_axb_2 ;
wire v_branch_result_3_axb_3 ;
wire v_branch_result_3_axb_4 ;
wire v_branch_result_3_cry_4 ;
wire v_branch_result_3_cry_3 ;
wire v_branch_result_3_cry_2 ;
wire v_branch_result_3_cry_1 ;
wire v_branch_result_3_cry_0 ;
wire N_3 ;
wire N_1 ;
input p_m_axis_output_tdata_0_rep2_Z_p_O_FDRE ;
input p_m_axis_output_tdata_0_rep1_Z_p_O_FDRE ;
input p_desc31_p_O_FDRE ;
input p_desc32_p_O_FDRE ;
input p_desc33_p_O_FDRE ;
input p_desc34_p_O_FDRE ;
input p_desc35_p_O_FDRE ;
input p_desc36_p_O_FDRE ;
input p_desc37_p_O_FDRE ;
// instances
  LUT2 v_branch_result_3_axb_0_cZ(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_3_axb_0));
defparam v_branch_result_3_axb_0_cZ.INIT=4'h9;
  p_O_FDRE m_axis_output_tdata_0_rep2_Z(.Q(branch_tdata_3_0_rep2),.D(v_branch_result_3_axb_0_i_rep2),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_0_rep2_Z_p_O_FDRE));
  p_O_FDRE m_axis_output_tdata_0_rep1_Z(.Q(branch_tdata_3_0_rep1),.D(v_branch_result_3_axb_0_i_rep1),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_0_rep1_Z_p_O_FDRE));
  p_O_FDRE desc31(.Q(branch_tdata_3_fast),.D(v_branch_result_3_axb_0_i_fast),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc31_p_O_FDRE));
  LUT3_L v_branch_result_3_axb_1_cZ(.I0(buffer_tdata_1),.I1(buffer_tdata_9),.I2(buffer_tdata_8),.LO(v_branch_result_3_axb_1));
defparam v_branch_result_3_axb_1_cZ.INIT=8'h69;
  LUT5_L v_branch_result_3_axb_5_cZ(.I0(buffer_tdata_10),.I1(buffer_tdata_9),.I2(buffer_tdata_11),.I3(buffer_tdata_3),.I4(buffer_tdata_8),.LO(v_branch_result_3_axb_5));
defparam v_branch_result_3_axb_5_cZ.INIT=32'h0FF00EF1;
  LUT4_L v_branch_result_3_axb_2_cZ(.I0(buffer_tdata_2),.I1(buffer_tdata_10),.I2(buffer_tdata_9),.I3(buffer_tdata_8),.LO(v_branch_result_3_axb_2));
defparam v_branch_result_3_axb_2_cZ.INIT=16'h6669;
  LUT5_L v_branch_result_3_axb_3_cZ(.I0(buffer_tdata_10),.I1(buffer_tdata_9),.I2(buffer_tdata_11),.I3(buffer_tdata_3),.I4(buffer_tdata_8),.LO(v_branch_result_3_axb_3));
defparam v_branch_result_3_axb_3_cZ.INIT=32'h0FF01EE1;
  LUT5_L v_branch_result_3_axb_4_cZ(.I0(buffer_tdata_10),.I1(buffer_tdata_9),.I2(buffer_tdata_11),.I3(buffer_tdata_3),.I4(buffer_tdata_8),.LO(v_branch_result_3_axb_4));
defparam v_branch_result_3_axb_4_cZ.INIT=32'h0FF00EF1;
  XORCY v_branch_result_3_s_5(.LI(v_branch_result_3_axb_5),.CI(v_branch_result_3_cry_4),.O(v_branch_result_3[5:5]));
  XORCY v_branch_result_3_s_4(.LI(v_branch_result_3_axb_4),.CI(v_branch_result_3_cry_3),.O(v_branch_result_3[4:4]));
  MUXCY_L v_branch_result_3_cry_4_cZ(.DI(N_2388_i),.CI(v_branch_result_3_cry_3),.S(v_branch_result_3_axb_4),.LO(v_branch_result_3_cry_4));
  XORCY v_branch_result_3_s_3(.LI(v_branch_result_3_axb_3),.CI(v_branch_result_3_cry_2),.O(v_branch_result_3[3:3]));
  MUXCY_L v_branch_result_3_cry_3_cZ(.DI(buffer_tdata_i[3:3]),.CI(v_branch_result_3_cry_2),.S(v_branch_result_3_axb_3),.LO(v_branch_result_3_cry_3));
  XORCY v_branch_result_3_s_2(.LI(v_branch_result_3_axb_2),.CI(v_branch_result_3_cry_1),.O(v_branch_result_3[2:2]));
  MUXCY_L v_branch_result_3_cry_2_cZ(.DI(buffer_tdata_i[2:2]),.CI(v_branch_result_3_cry_1),.S(v_branch_result_3_axb_2),.LO(v_branch_result_3_cry_2));
  XORCY v_branch_result_3_s_1(.LI(v_branch_result_3_axb_1),.CI(v_branch_result_3_cry_0),.O(v_branch_result_3[1:1]));
  MUXCY_L v_branch_result_3_cry_1_cZ(.DI(buffer_tdata_i[1:1]),.CI(v_branch_result_3_cry_0),.S(v_branch_result_3_axb_1),.LO(v_branch_result_3_cry_1));
  MUXCY_L v_branch_result_3_cry_0_cZ(.DI(buffer_tdata_8),.CI(VCC),.S(v_branch_result_3_axb_0),.LO(v_branch_result_3_cry_0));
  p_O_FDRE desc32(.Q(branch_tdata_3[5:5]),.D(v_branch_result_3[5:5]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc32_p_O_FDRE));
  p_O_FDRE desc33(.Q(branch_tdata_3[4:4]),.D(v_branch_result_3[4:4]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc33_p_O_FDRE));
  p_O_FDRE desc34(.Q(branch_tdata_3[3:3]),.D(v_branch_result_3[3:3]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc34_p_O_FDRE));
  p_O_FDRE desc35(.Q(branch_tdata_3[2:2]),.D(v_branch_result_3[2:2]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc35_p_O_FDRE));
  p_O_FDRE desc36(.Q(branch_tdata_3[1:1]),.D(v_branch_result_3[1:1]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc36_p_O_FDRE));
  p_O_FDRE desc37(.Q(branch_tdata_3[0:0]),.D(v_branch_result_3_axb_0_i),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc37_p_O_FDRE));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT2 v_branch_result_3_axb_0_i_0_fast_lut6_2_o6(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_3_axb_0_i_fast));
defparam v_branch_result_3_axb_0_i_0_fast_lut6_2_o6.INIT=4'h6;
  LUT2 v_branch_result_3_axb_0_i_0_fast_lut6_2_o5(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_3_axb_0_i_rep2));
defparam v_branch_result_3_axb_0_i_0_fast_lut6_2_o5.INIT=4'h6;
  LUT2 v_branch_result_3_axb_0_i_0_lut6_2_o6(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_3_axb_0_i));
defparam v_branch_result_3_axb_0_i_0_lut6_2_o6.INIT=4'h6;
  LUT2 v_branch_result_3_axb_0_i_0_lut6_2_o5(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_3_axb_0_i_rep1));
defparam v_branch_result_3_axb_0_i_0_lut6_2_o5.INIT=4'h6;
endmodule
module branch_distanceZ2_inj (branch_tdata_2_fast,buffer_tdata_0,buffer_tdata_8,buffer_tdata_11,buffer_tdata_3,buffer_tdata_2,buffer_tdata_10,buffer_tdata_1,buffer_tdata_9,branch_tdata_2_5,branch_tdata_2_3,branch_tdata_2_2,branch_tdata_2_1,branch_tdata_2_0,un10_v_branch_result_axb_0_i_rep2,un10_v_branch_result_axb_0_i_fast,un10_v_branch_result_axb_0_i_rep1,branch_tdata_2_0_rep2,aclk,aresetn_i,un1_output_accept,branch_tdata_2_0_rep1,v_branch_result_axb_0_i_fast,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE,p_desc39_p_O_FDRE,p_desc52_p_O_FDRE,p_desc53_p_O_FDRE,p_desc54_p_O_FDRE,p_desc55_p_O_FDRE,p_desc56_p_O_FDRE);
output branch_tdata_2_fast ;
input buffer_tdata_0 ;
input buffer_tdata_8 ;
input buffer_tdata_11 ;
input buffer_tdata_3 ;
input buffer_tdata_2 ;
input buffer_tdata_10 ;
input buffer_tdata_1 ;
input buffer_tdata_9 ;
output branch_tdata_2_5 ;
output branch_tdata_2_3 ;
output branch_tdata_2_2 ;
output branch_tdata_2_1 ;
output branch_tdata_2_0 ;
output un10_v_branch_result_axb_0_i_rep2 ;
output un10_v_branch_result_axb_0_i_fast ;
output un10_v_branch_result_axb_0_i_rep1 ;
output branch_tdata_2_0_rep2 ;
input aclk ;
input aresetn_i ;
input un1_output_accept ;
output branch_tdata_2_0_rep1 ;
input v_branch_result_axb_0_i_fast ;
wire buffer_tdata_0 ;
wire buffer_tdata_8 ;
wire buffer_tdata_11 ;
wire buffer_tdata_3 ;
wire buffer_tdata_2 ;
wire buffer_tdata_10 ;
wire buffer_tdata_1 ;
wire buffer_tdata_9 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_0 ;
wire un10_v_branch_result_axb_0_i_rep2 ;
wire un10_v_branch_result_axb_0_i_fast ;
wire un10_v_branch_result_axb_0_i_rep1 ;
wire branch_tdata_2_0_rep2 ;
wire aclk ;
wire aresetn_i ;
wire un1_output_accept ;
wire branch_tdata_2_0_rep1 ;
wire v_branch_result_axb_0_i_fast ;
wire [31:28] v_branch_result ;
wire GND ;
wire VCC ;
wire v_branch_result_axb_0_i ;
wire v_branch_result_axb_0_i_rep1 ;
wire v_branch_result_axb_0_i_rep2 ;
wire v_branch_result_axb_0 ;
wire v_branch_result_axb_4 ;
wire v_branch_result_axb_3 ;
wire v_branch_result_axb_2 ;
wire v_branch_result_axb_1 ;
wire v_branch_result_cry_3 ;
wire v_branch_result_cry_2 ;
wire v_branch_result_cry_1 ;
wire v_branch_result_cry_0 ;
wire N_2 ;
wire N_1 ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE ;
input p_desc39_p_O_FDRE ;
input p_desc52_p_O_FDRE ;
input p_desc53_p_O_FDRE ;
input p_desc54_p_O_FDRE ;
input p_desc55_p_O_FDRE ;
input p_desc56_p_O_FDRE ;
// instances
  LUT2 desc38(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_axb_0));
defparam desc38.INIT=4'h9;
  p_O_FDRE m_axis_output_tdata_1_0_rep2_Z(.Q(branch_tdata_2_0_rep2),.D(v_branch_result_axb_0_i_rep2),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE));
  p_O_FDRE m_axis_output_tdata_1_0_rep1_Z(.Q(branch_tdata_2_0_rep1),.D(v_branch_result_axb_0_i_rep1),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE));
  p_O_FDRE desc39(.Q(branch_tdata_2_fast),.D(v_branch_result_axb_0_i_fast),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc39_p_O_FDRE));
  LUT2_L desc40(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(v_branch_result_axb_4));
defparam desc40.INIT=4'h9;
  LUT2_L desc41(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(v_branch_result_axb_3));
defparam desc41.INIT=4'h9;
  LUT2_L desc42(.I0(buffer_tdata_2),.I1(buffer_tdata_10),.LO(v_branch_result_axb_2));
defparam desc42.INIT=4'h9;
  LUT2_L desc43(.I0(buffer_tdata_1),.I1(buffer_tdata_9),.LO(v_branch_result_axb_1));
defparam desc43.INIT=4'h9;
  XORCY desc44(.LI(v_branch_result_axb_4),.CI(v_branch_result_cry_3),.O(v_branch_result[31:31]));
  XORCY desc45(.LI(v_branch_result_axb_3),.CI(v_branch_result_cry_2),.O(v_branch_result[30:30]));
  MUXCY_L desc46(.DI(buffer_tdata_11),.CI(v_branch_result_cry_2),.S(v_branch_result_axb_3),.LO(v_branch_result_cry_3));
  XORCY desc47(.LI(v_branch_result_axb_2),.CI(v_branch_result_cry_1),.O(v_branch_result[29:29]));
  MUXCY_L desc48(.DI(buffer_tdata_10),.CI(v_branch_result_cry_1),.S(v_branch_result_axb_2),.LO(v_branch_result_cry_2));
  XORCY desc49(.LI(v_branch_result_axb_1),.CI(v_branch_result_cry_0),.O(v_branch_result[28:28]));
  MUXCY_L desc50(.DI(buffer_tdata_9),.CI(v_branch_result_cry_0),.S(v_branch_result_axb_1),.LO(v_branch_result_cry_1));
  MUXCY_L desc51(.DI(buffer_tdata_8),.CI(VCC),.S(v_branch_result_axb_0),.LO(v_branch_result_cry_0));
  p_O_FDRE desc52(.Q(branch_tdata_2_5),.D(v_branch_result[31:31]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc52_p_O_FDRE));
  p_O_FDRE desc53(.Q(branch_tdata_2_3),.D(v_branch_result[30:30]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc53_p_O_FDRE));
  p_O_FDRE desc54(.Q(branch_tdata_2_2),.D(v_branch_result[29:29]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc54_p_O_FDRE));
  p_O_FDRE desc55(.Q(branch_tdata_2_1),.D(v_branch_result[28:28]),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc55_p_O_FDRE));
  p_O_FDRE desc56(.Q(branch_tdata_2_0),.D(v_branch_result_axb_0_i),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc56_p_O_FDRE));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT2 desc57(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_axb_0_i_rep2));
defparam desc57.INIT=4'h6;
  LUT2 desc58(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un10_v_branch_result_axb_0_i_rep1));
defparam desc58.INIT=4'h6;
  LUT2 desc59(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_axb_0_i_rep1));
defparam desc59.INIT=4'h6;
  LUT2 desc60(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un10_v_branch_result_axb_0_i_fast));
defparam desc60.INIT=4'h6;
  LUT2 desc61(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_axb_0_i));
defparam desc61.INIT=4'h6;
  LUT2 desc62(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un10_v_branch_result_axb_0_i_rep2));
defparam desc62.INIT=4'h6;
endmodule
module branch_distanceZ0_inj (branch_tlast,branch_tdata_0_fast,buffer_tdata_11,buffer_tdata_3,buffer_tdata_2,buffer_tdata_10,buffer_tdata_1,buffer_tdata_9,buffer_tdata_0,buffer_tdata_8,acs_tvalid,write_ram_fsm,branch_tvalid,branch_tdata_0_5,branch_tdata_0_3,branch_tdata_0_2,branch_tdata_0_1,branch_tdata_0_0,aclk,aresetn_i,branch_tdata_0_0_rep2,un1_output_accept,branch_tdata_0_0_rep1,write_ram_fsm_0_rep1,buffer_tvalid,write_ram_fsm_4_rep1,N_1756_1,buffer_tlast,un27_s_axis_input_tready_int,s_axis_inbranch_tlast_d_RNIIAVE1_O5,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE,p_desc63_p_O_FDRE,p_desc78_p_O_FDRE,p_desc79_p_O_FDRE,p_desc80_p_O_FDRE,p_desc81_p_O_FDRE,p_desc82_p_O_FDRE);
output branch_tlast ;
output branch_tdata_0_fast ;
input buffer_tdata_11 ;
input buffer_tdata_3 ;
input buffer_tdata_2 ;
input buffer_tdata_10 ;
input buffer_tdata_1 ;
input buffer_tdata_9 ;
input buffer_tdata_0 ;
input buffer_tdata_8 ;
input acs_tvalid ;
input [1:1] write_ram_fsm ;
output branch_tvalid ;
output branch_tdata_0_5 ;
output branch_tdata_0_3 ;
output branch_tdata_0_2 ;
output branch_tdata_0_1 ;
output branch_tdata_0_0 ;
input aclk ;
input aresetn_i ;
output branch_tdata_0_0_rep2 ;
output un1_output_accept ;
output branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep1 ;
input buffer_tvalid ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input buffer_tlast ;
input un27_s_axis_input_tready_int ;
input s_axis_inbranch_tlast_d_RNIIAVE1_O5 ;
wire buffer_tdata_11 ;
wire buffer_tdata_3 ;
wire buffer_tdata_2 ;
wire buffer_tdata_10 ;
wire buffer_tdata_1 ;
wire buffer_tdata_9 ;
wire buffer_tdata_0 ;
wire buffer_tdata_8 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_0 ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire un1_output_accept ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep1 ;
wire buffer_tvalid ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire buffer_tlast ;
wire un27_s_axis_input_tready_int ;
wire s_axis_inbranch_tlast_d_RNIIAVE1_O5 ;
wire m_axis_output_tlast ;
wire un7_v_branch_result_axb_0 ;
wire un7_v_branch_result_axb_4 ;
wire un7_v_branch_result_axb_3 ;
wire un7_v_branch_result_axb_2 ;
wire un7_v_branch_result_axb_1 ;
wire un7_v_branch_result_cry_3 ;
wire un7_v_branch_result_s_4 ;
wire un7_v_branch_result_cry_2 ;
wire un7_v_branch_result_s_3 ;
wire un7_v_branch_result_cry_1 ;
wire un7_v_branch_result_s_2 ;
wire un7_v_branch_result_cry_0 ;
wire un7_v_branch_result_s_1 ;
wire GND ;
wire VCC ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE ;
input p_desc63_p_O_FDRE ;
input p_desc78_p_O_FDRE ;
input p_desc79_p_O_FDRE ;
input p_desc80_p_O_FDRE ;
input p_desc81_p_O_FDRE ;
input p_desc82_p_O_FDRE ;
// instances
  FDR m_axis_output_tlast_Z(.Q(branch_tlast),.D(m_axis_output_tlast),.C(aclk),.R(aresetn_i));
  p_O_FDRE m_axis_output_tdata_1_0_rep2_Z(.Q(branch_tdata_0_0_rep2),.D(un7_v_branch_result_axb_0),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE));
  p_O_FDRE m_axis_output_tdata_1_0_rep1_Z(.Q(branch_tdata_0_0_rep1),.D(un7_v_branch_result_axb_0),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE));
  p_O_FDRE desc63(.Q(branch_tdata_0_fast),.D(un7_v_branch_result_axb_0),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc63_p_O_FDRE));
  LUT2_L desc64(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(un7_v_branch_result_axb_4));
defparam desc64.INIT=4'h6;
  LUT2_L desc65(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(un7_v_branch_result_axb_3));
defparam desc65.INIT=4'h6;
  LUT2_L desc66(.I0(buffer_tdata_2),.I1(buffer_tdata_10),.LO(un7_v_branch_result_axb_2));
defparam desc66.INIT=4'h6;
  LUT2_L desc67(.I0(buffer_tdata_1),.I1(buffer_tdata_9),.LO(un7_v_branch_result_axb_1));
defparam desc67.INIT=4'h6;
  LUT2 desc68(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un7_v_branch_result_axb_0));
defparam desc68.INIT=4'h6;
  LUT6 desc69(.I0(write_ram_fsm_0_rep1),.I1(buffer_tvalid),.I2(write_ram_fsm_4_rep1),.I3(acs_tvalid),.I4(write_ram_fsm[1:1]),.I5(N_1756_1),.O(un1_output_accept));
defparam desc69.INIT=64'h00CC04CC00CC00CC;
  LUT6_L m_axis_output_tlast_e(.I0(buffer_tlast),.I1(buffer_tvalid),.I2(acs_tvalid),.I3(branch_tlast),.I4(branch_tvalid),.I5(un27_s_axis_input_tready_int),.LO(m_axis_output_tlast));
defparam m_axis_output_tlast_e.INIT=64'hF808FB088888BB88;
  FDR m_axis_output_tvalid_int_Z(.Q(branch_tvalid),.D(s_axis_inbranch_tlast_d_RNIIAVE1_O5),.C(aclk),.R(aresetn_i));
  XORCY desc70(.LI(un7_v_branch_result_axb_4),.CI(un7_v_branch_result_cry_3),.O(un7_v_branch_result_s_4));
  XORCY desc71(.LI(un7_v_branch_result_axb_3),.CI(un7_v_branch_result_cry_2),.O(un7_v_branch_result_s_3));
  MUXCY_L desc72(.DI(buffer_tdata_3),.CI(un7_v_branch_result_cry_2),.S(un7_v_branch_result_axb_3),.LO(un7_v_branch_result_cry_3));
  XORCY desc73(.LI(un7_v_branch_result_axb_2),.CI(un7_v_branch_result_cry_1),.O(un7_v_branch_result_s_2));
  MUXCY_L desc74(.DI(buffer_tdata_2),.CI(un7_v_branch_result_cry_1),.S(un7_v_branch_result_axb_2),.LO(un7_v_branch_result_cry_2));
  XORCY desc75(.LI(un7_v_branch_result_axb_1),.CI(un7_v_branch_result_cry_0),.O(un7_v_branch_result_s_1));
  MUXCY_L desc76(.DI(buffer_tdata_1),.CI(un7_v_branch_result_cry_0),.S(un7_v_branch_result_axb_1),.LO(un7_v_branch_result_cry_1));
  MUXCY_L desc77(.DI(buffer_tdata_0),.CI(GND),.S(un7_v_branch_result_axb_0),.LO(un7_v_branch_result_cry_0));
  p_O_FDRE desc78(.Q(branch_tdata_0_5),.D(un7_v_branch_result_s_4),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc78_p_O_FDRE));
  p_O_FDRE desc79(.Q(branch_tdata_0_3),.D(un7_v_branch_result_s_3),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc79_p_O_FDRE));
  p_O_FDRE desc80(.Q(branch_tdata_0_2),.D(un7_v_branch_result_s_2),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc80_p_O_FDRE));
  p_O_FDRE desc81(.Q(branch_tdata_0_1),.D(un7_v_branch_result_s_1),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc81_p_O_FDRE));
  p_O_FDRE desc82(.Q(branch_tdata_0_0),.D(un7_v_branch_result_axb_0),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc82_p_O_FDRE));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module branch_distanceZ1_inj (branch_tdata_1_fast,buffer_tdata_0,buffer_tdata_8,buffer_tdata_11,buffer_tdata_3,buffer_tdata_1,buffer_tdata_9,buffer_tdata_2,buffer_tdata_10,branch_tdata_1_5,branch_tdata_1_3,branch_tdata_1_2,branch_tdata_1_1,branch_tdata_1_0,v_branch_result_axb_0_i_fast,branch_tdata_1_0_rep2,un10_v_branch_result_axb_0_i_rep2,aclk,aresetn_i,un1_output_accept,branch_tdata_1_0_rep1,un10_v_branch_result_axb_0_i_rep1,un10_v_branch_result_axb_0_i_fast,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE,p_desc83_p_O_FDRE,p_desc84_p_O_FDRE,p_desc85_p_O_FDRE,p_desc86_p_O_FDRE,p_desc87_p_O_FDRE,p_desc88_p_O_FDRE);
output branch_tdata_1_fast ;
input buffer_tdata_0 ;
input buffer_tdata_8 ;
input buffer_tdata_11 ;
input buffer_tdata_3 ;
input buffer_tdata_1 ;
input buffer_tdata_9 ;
input buffer_tdata_2 ;
input buffer_tdata_10 ;
output branch_tdata_1_5 ;
output branch_tdata_1_3 ;
output branch_tdata_1_2 ;
output branch_tdata_1_1 ;
output branch_tdata_1_0 ;
output v_branch_result_axb_0_i_fast ;
output branch_tdata_1_0_rep2 ;
input un10_v_branch_result_axb_0_i_rep2 ;
input aclk ;
input aresetn_i ;
input un1_output_accept ;
output branch_tdata_1_0_rep1 ;
input un10_v_branch_result_axb_0_i_rep1 ;
input un10_v_branch_result_axb_0_i_fast ;
wire buffer_tdata_0 ;
wire buffer_tdata_8 ;
wire buffer_tdata_11 ;
wire buffer_tdata_3 ;
wire buffer_tdata_1 ;
wire buffer_tdata_9 ;
wire buffer_tdata_2 ;
wire buffer_tdata_10 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_0 ;
wire v_branch_result_axb_0_i_fast ;
wire branch_tdata_1_0_rep2 ;
wire un10_v_branch_result_axb_0_i_rep2 ;
wire aclk ;
wire aresetn_i ;
wire un1_output_accept ;
wire branch_tdata_1_0_rep1 ;
wire un10_v_branch_result_axb_0_i_rep1 ;
wire un10_v_branch_result_axb_0_i_fast ;
wire GND ;
wire VCC ;
wire un10_v_branch_result_axb_0_i ;
wire un10_v_branch_result_axb_0 ;
wire un10_v_branch_result_axb_4 ;
wire un10_v_branch_result_axb_1 ;
wire un10_v_branch_result_axb_2 ;
wire un10_v_branch_result_axb_3 ;
wire un10_v_branch_result_cry_3 ;
wire un10_v_branch_result_s_4 ;
wire un10_v_branch_result_cry_2 ;
wire un10_v_branch_result_s_3 ;
wire un10_v_branch_result_cry_1 ;
wire un10_v_branch_result_s_2 ;
wire un10_v_branch_result_cry_0 ;
wire un10_v_branch_result_s_1 ;
wire N_1 ;
wire N_1_0 ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE ;
input p_desc83_p_O_FDRE ;
input p_desc84_p_O_FDRE ;
input p_desc85_p_O_FDRE ;
input p_desc86_p_O_FDRE ;
input p_desc87_p_O_FDRE ;
input p_desc88_p_O_FDRE ;
// instances
  LUT2 un10_v_branch_result_cry_0_RNO(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un10_v_branch_result_axb_0));
defparam un10_v_branch_result_cry_0_RNO.INIT=4'h9;
  p_O_FDRE m_axis_output_tdata_1_0_rep2_Z(.Q(branch_tdata_1_0_rep2),.D(un10_v_branch_result_axb_0_i_rep2),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE));
  p_O_FDRE m_axis_output_tdata_1_0_rep1_Z(.Q(branch_tdata_1_0_rep1),.D(un10_v_branch_result_axb_0_i_rep1),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE));
  p_O_FDRE desc83(.Q(branch_tdata_1_fast),.D(un10_v_branch_result_axb_0_i_fast),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc83_p_O_FDRE));
  LUT2_L un10_v_branch_result_axb_4_cZ(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(un10_v_branch_result_axb_4));
defparam un10_v_branch_result_axb_4_cZ.INIT=4'h9;
  LUT2_L un10_v_branch_result_axb_1_cZ(.I0(buffer_tdata_1),.I1(buffer_tdata_9),.LO(un10_v_branch_result_axb_1));
defparam un10_v_branch_result_axb_1_cZ.INIT=4'h9;
  LUT2_L un10_v_branch_result_axb_2_cZ(.I0(buffer_tdata_2),.I1(buffer_tdata_10),.LO(un10_v_branch_result_axb_2));
defparam un10_v_branch_result_axb_2_cZ.INIT=4'h9;
  LUT2_L un10_v_branch_result_axb_3_cZ(.I0(buffer_tdata_11),.I1(buffer_tdata_3),.LO(un10_v_branch_result_axb_3));
defparam un10_v_branch_result_axb_3_cZ.INIT=4'h9;
  XORCY un10_v_branch_result_s_4_cZ(.LI(un10_v_branch_result_axb_4),.CI(un10_v_branch_result_cry_3),.O(un10_v_branch_result_s_4));
  XORCY un10_v_branch_result_s_3_cZ(.LI(un10_v_branch_result_axb_3),.CI(un10_v_branch_result_cry_2),.O(un10_v_branch_result_s_3));
  MUXCY_L un10_v_branch_result_cry_3_cZ(.DI(buffer_tdata_3),.CI(un10_v_branch_result_cry_2),.S(un10_v_branch_result_axb_3),.LO(un10_v_branch_result_cry_3));
  XORCY un10_v_branch_result_s_2_cZ(.LI(un10_v_branch_result_axb_2),.CI(un10_v_branch_result_cry_1),.O(un10_v_branch_result_s_2));
  MUXCY_L un10_v_branch_result_cry_2_cZ(.DI(buffer_tdata_2),.CI(un10_v_branch_result_cry_1),.S(un10_v_branch_result_axb_2),.LO(un10_v_branch_result_cry_2));
  XORCY un10_v_branch_result_s_1_cZ(.LI(un10_v_branch_result_axb_1),.CI(un10_v_branch_result_cry_0),.O(un10_v_branch_result_s_1));
  MUXCY_L un10_v_branch_result_cry_1_cZ(.DI(buffer_tdata_1),.CI(un10_v_branch_result_cry_0),.S(un10_v_branch_result_axb_1),.LO(un10_v_branch_result_cry_1));
  MUXCY_L un10_v_branch_result_cry_0_cZ(.DI(buffer_tdata_0),.CI(VCC),.S(un10_v_branch_result_axb_0),.LO(un10_v_branch_result_cry_0));
  p_O_FDRE desc84(.Q(branch_tdata_1_5),.D(un10_v_branch_result_s_4),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc84_p_O_FDRE));
  p_O_FDRE desc85(.Q(branch_tdata_1_3),.D(un10_v_branch_result_s_3),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc85_p_O_FDRE));
  p_O_FDRE desc86(.Q(branch_tdata_1_2),.D(un10_v_branch_result_s_2),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc86_p_O_FDRE));
  p_O_FDRE desc87(.Q(branch_tdata_1_1),.D(un10_v_branch_result_s_1),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc87_p_O_FDRE));
  p_O_FDRE desc88(.Q(branch_tdata_1_0),.D(un10_v_branch_result_axb_0_i),.C(aclk),.R(aresetn_i),.CE(un1_output_accept),.E(p_desc88_p_O_FDRE));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT2 un10_v_branch_result_axb_0_i_0_lut6_2_o6(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(un10_v_branch_result_axb_0_i));
defparam un10_v_branch_result_axb_0_i_0_lut6_2_o6.INIT=4'h6;
  LUT2 un10_v_branch_result_axb_0_i_0_lut6_2_o5(.I0(buffer_tdata_0),.I1(buffer_tdata_8),.O(v_branch_result_axb_0_i_fast));
defparam un10_v_branch_result_axb_0_i_0_lut6_2_o5.INIT=4'h6;
endmodule
module acsZ0_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_50,acs_prob_tdata_51,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_57,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,N_1756_1,aresetn,p_desc95_p_O_FD,p_desc96_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc125_p_O_FDRE);
input branch_tlast ;
output [57:57] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_50 ;
input [8:0] acs_prob_tdata_51 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_57 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIT11R_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNISNV71 ;
wire un4_v_high_s_7 ;
wire un4_v_low_s_7 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8 ;
wire un4_v_low_s_8 ;
wire un4_v_high_s_6 ;
wire un4_v_low_s_6 ;
wire un4_v_high_s_5 ;
wire un4_v_low_s_5 ;
wire un4_v_high_s_4 ;
wire un4_v_low_s_4 ;
wire un4_v_high_s_3 ;
wire un4_v_low_s_3 ;
wire un4_v_high_s_2 ;
wire un4_v_low_s_2 ;
wire un4_v_high_s_1 ;
wire un4_v_low_s_1 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire N_2368 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire GND ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire N_1 ;
input p_desc95_p_O_FD ;
input p_desc96_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc125_p_O_FDRE ;
// instances
  FDR desc89(.Q(acs_prob_tdata_57[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  FDR desc90(.Q(acs_prob_tdata_57[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  FDR desc91(.Q(acs_prob_tdata_57[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  FDR desc92(.Q(acs_prob_tdata_57[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  FDR desc93(.Q(acs_prob_tdata_57[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  FDR desc94(.Q(acs_prob_tdata_57[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71));
  p_O_FD desc95(.Q(acs_prob_tdata_57[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc95_p_O_FD));
  p_O_FD desc96(.Q(acs_prob_tdata_57[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc96_p_O_FD));
  LUT6 desc97(.I0(un4_v_high_s_7),.I1(un4_v_low_s_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISNV71),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc97.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc98(.I0(un4_v_high_s_8),.I1(un4_v_low_s_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISNV71),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc98.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc99(.I0(un4_v_high_s_6),.I1(un4_v_low_s_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc99.INIT=32'hACACFF00;
  LUT5 desc100(.I0(un4_v_high_s_5),.I1(un4_v_low_s_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc100.INIT=32'hACACFF00;
  LUT5 desc101(.I0(un4_v_high_s_4),.I1(un4_v_low_s_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc101.INIT=32'hACACFF00;
  LUT5 desc102(.I0(un4_v_high_s_3),.I1(un4_v_low_s_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc102.INIT=32'hACACFF00;
  LUT5 desc103(.I0(un4_v_high_s_2),.I1(un4_v_low_s_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc103.INIT=32'hACACFF00;
  LUT5 desc104(.I0(un4_v_high_s_1),.I1(un4_v_low_s_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_57[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc104.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[57:57]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_51[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_51[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_51[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_51[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_51[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_51[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_51[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_51[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc105(.I0(acs_prob_tdata_50[0:0]),.I1(acs_prob_tdata_51[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc105.INIT=16'h9669;
  LUT2 desc106(.I0(un4_v_high_s_1),.I1(un4_v_low_s_1),.O(v_diff_1_axb_1));
defparam desc106.INIT=4'h9;
  LUT2 desc107(.I0(un4_v_high_s_2),.I1(un4_v_low_s_2),.O(v_diff_1_axb_2));
defparam desc107.INIT=4'h9;
  LUT2 desc108(.I0(un4_v_high_s_3),.I1(un4_v_low_s_3),.O(v_diff_1_axb_3));
defparam desc108.INIT=4'h9;
  LUT2 desc109(.I0(un4_v_high_s_4),.I1(un4_v_low_s_4),.O(v_diff_1_axb_4));
defparam desc109.INIT=4'h9;
  LUT2 desc110(.I0(un4_v_high_s_5),.I1(un4_v_low_s_5),.O(v_diff_1_axb_5));
defparam desc110.INIT=4'h9;
  LUT2 desc111(.I0(un4_v_high_s_6),.I1(un4_v_low_s_6),.O(v_diff_1_axb_6));
defparam desc111.INIT=4'h9;
  LUT2 desc112(.I0(un4_v_high_s_7),.I1(un4_v_low_s_7),.O(v_diff_1_axb_7));
defparam desc112.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_50[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_50[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_50[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_50[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_50[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_50[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_50[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc113(.I0(acs_prob_tdata_50[0:0]),.I1(acs_prob_tdata_51[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2368));
defparam desc113.INIT=32'h3C3C55AA;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_50[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc114(.I0(un4_v_high_s_8),.I1(un4_v_low_s_8),.O(v_diff_1_axb_8));
defparam desc114.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_51[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT6 desc115(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc115.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIALQ41(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIALQ41.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNISNV71_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNISNV71));
defparam s_axis_inbranch_tlast_d_RNISNV71_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_50[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIT11R_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_low_s_8_cZ(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8));
  XORCY un4_v_low_s_7_cZ(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_50[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6_cZ(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_50[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5_cZ(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_50[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4_cZ(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_50[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3_cZ(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_50[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2_cZ(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_50[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1_cZ(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_50[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_50[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc116(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc117(.DI(un4_v_low_s_7),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc118(.DI(un4_v_low_s_6),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc119(.DI(un4_v_low_s_5),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc120(.DI(un4_v_low_s_4),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc121(.DI(un4_v_low_s_3),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc122(.DI(un4_v_low_s_2),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc123(.DI(un4_v_low_s_1),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc124(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8_cZ(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8));
  XORCY un4_v_high_s_7_cZ(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_51[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6_cZ(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_51[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5_cZ(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_51[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4_cZ(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_51[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3_cZ(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_51[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2_cZ(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_51[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1_cZ(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_51[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_51[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  p_O_FDRE desc125(.Q(acs_prob_tdata_57[0:0]),.D(N_2368),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISNV71),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc125_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc126(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIT11R_O6));
defparam desc126.INIT=16'hF4F0;
  LUT2 desc127(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc127.INIT=4'h8;
endmodule
module acsZ0_1_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_25,acs_prob_tdata_24,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_12,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc134_p_O_FD,p_desc135_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc164_p_O_FDRE);
input branch_tlast ;
output [12:12] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_25 ;
input [8:0] acs_prob_tdata_24 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_12 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI2FB11_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIAKN81 ;
wire un4_v_high_s_7_0 ;
wire un4_v_low_s_7_0 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_0 ;
wire un4_v_low_s_8_0 ;
wire un4_v_high_s_6_0 ;
wire un4_v_low_s_6_0 ;
wire un4_v_high_s_5_0 ;
wire un4_v_low_s_5_0 ;
wire un4_v_high_s_4_0 ;
wire un4_v_low_s_4_0 ;
wire un4_v_high_s_3_0 ;
wire un4_v_low_s_3_0 ;
wire un4_v_high_s_2_0 ;
wire un4_v_low_s_2_0 ;
wire un4_v_high_s_1_0 ;
wire un4_v_low_s_1_0 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2348 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc134_p_O_FD ;
input p_desc135_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc164_p_O_FDRE ;
// instances
  FDR desc128(.Q(acs_prob_tdata_12[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  FDR desc129(.Q(acs_prob_tdata_12[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  FDR desc130(.Q(acs_prob_tdata_12[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  FDR desc131(.Q(acs_prob_tdata_12[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  FDR desc132(.Q(acs_prob_tdata_12[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  FDR desc133(.Q(acs_prob_tdata_12[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81));
  p_O_FD desc134(.Q(acs_prob_tdata_12[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc134_p_O_FD));
  p_O_FD desc135(.Q(acs_prob_tdata_12[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc135_p_O_FD));
  LUT6 desc136(.I0(un4_v_high_s_7_0),.I1(un4_v_low_s_7_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAKN81),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc136.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc137(.I0(un4_v_high_s_8_0),.I1(un4_v_low_s_8_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAKN81),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc137.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc138(.I0(un4_v_high_s_6_0),.I1(un4_v_low_s_6_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc138.INIT=32'hACACFF00;
  LUT5 desc139(.I0(un4_v_high_s_5_0),.I1(un4_v_low_s_5_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc139.INIT=32'hACACFF00;
  LUT5 desc140(.I0(un4_v_high_s_4_0),.I1(un4_v_low_s_4_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc140.INIT=32'hACACFF00;
  LUT5 desc141(.I0(un4_v_high_s_3_0),.I1(un4_v_low_s_3_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc141.INIT=32'hACACFF00;
  LUT5 desc142(.I0(un4_v_high_s_2_0),.I1(un4_v_low_s_2_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc142.INIT=32'hACACFF00;
  LUT5 desc143(.I0(un4_v_high_s_1_0),.I1(un4_v_low_s_1_0),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_12[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc143.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[12:12]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc144(.I0(acs_prob_tdata_24[0:0]),.I1(acs_prob_tdata_25[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc144.INIT=16'h9669;
  LUT2 desc145(.I0(un4_v_high_s_1_0),.I1(un4_v_low_s_1_0),.O(v_diff_1_axb_1));
defparam desc145.INIT=4'h9;
  LUT2 desc146(.I0(un4_v_high_s_2_0),.I1(un4_v_low_s_2_0),.O(v_diff_1_axb_2));
defparam desc146.INIT=4'h9;
  LUT2 desc147(.I0(un4_v_high_s_3_0),.I1(un4_v_low_s_3_0),.O(v_diff_1_axb_3));
defparam desc147.INIT=4'h9;
  LUT2 desc148(.I0(un4_v_high_s_4_0),.I1(un4_v_low_s_4_0),.O(v_diff_1_axb_4));
defparam desc148.INIT=4'h9;
  LUT2 desc149(.I0(un4_v_high_s_5_0),.I1(un4_v_low_s_5_0),.O(v_diff_1_axb_5));
defparam desc149.INIT=4'h9;
  LUT2 desc150(.I0(un4_v_high_s_6_0),.I1(un4_v_low_s_6_0),.O(v_diff_1_axb_6));
defparam desc150.INIT=4'h9;
  LUT2 desc151(.I0(un4_v_high_s_7_0),.I1(un4_v_low_s_7_0),.O(v_diff_1_axb_7));
defparam desc151.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_24[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_24[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_24[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_24[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_24[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_24[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_24[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_25[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_25[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_25[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_25[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_25[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_25[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_25[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_25[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc152(.I0(acs_prob_tdata_24[0:0]),.I1(acs_prob_tdata_25[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2348));
defparam desc152.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_25[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_24[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc153(.I0(un4_v_high_s_8_0),.I1(un4_v_low_s_8_0),.O(v_diff_1_axb_8));
defparam desc153.INIT=4'h9;
  LUT6 desc154(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc154.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIOHI51(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIOHI51.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIAKN81_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIAKN81));
defparam s_axis_inbranch_tlast_d_RNIAKN81_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_24[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI2FB11_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_0));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_0));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_25[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_0));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_25[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_0));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_25[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_0));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_25[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_0));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_25[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_0));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_25[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_0));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_25[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_25[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_0));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_0));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_24[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_0));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_24[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_0));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_24[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_0));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_24[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_0));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_24[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_0));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_24[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_0));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_24[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_24[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc155(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc156(.DI(un4_v_low_s_7_0),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc157(.DI(un4_v_low_s_6_0),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc158(.DI(un4_v_low_s_5_0),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc159(.DI(un4_v_low_s_4_0),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc160(.DI(un4_v_low_s_3_0),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc161(.DI(un4_v_low_s_2_0),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc162(.DI(un4_v_low_s_1_0),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc163(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc164(.Q(acs_prob_tdata_12[0:0]),.D(N_2348),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAKN81),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc164_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc165(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI2FB11_O6));
defparam desc165.INIT=16'hF4F0;
  LUT2 desc166(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc166.INIT=4'h8;
endmodule
module acsZ0_2_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_45,acs_prob_tdata_44,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_54,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,N_1756_1,aresetn,p_desc173_p_O_FD,p_desc174_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc203_p_O_FDRE);
input branch_tlast ;
output [54:54] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_45 ;
input [8:0] acs_prob_tdata_44 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_54 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIKV121_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIMEM11 ;
wire un4_v_high_s_7_1 ;
wire un4_v_low_s_7_1 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_1 ;
wire un4_v_low_s_8_1 ;
wire un4_v_high_s_6_1 ;
wire un4_v_low_s_6_1 ;
wire un4_v_high_s_5_1 ;
wire un4_v_low_s_5_1 ;
wire un4_v_high_s_4_1 ;
wire un4_v_low_s_4_1 ;
wire un4_v_high_s_3_1 ;
wire un4_v_low_s_3_1 ;
wire un4_v_high_s_2_1 ;
wire un4_v_low_s_2_1 ;
wire un4_v_high_s_1_1 ;
wire un4_v_low_s_1_1 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2328 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc173_p_O_FD ;
input p_desc174_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc203_p_O_FDRE ;
// instances
  FDR desc167(.Q(acs_prob_tdata_54[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  FDR desc168(.Q(acs_prob_tdata_54[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  FDR desc169(.Q(acs_prob_tdata_54[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  FDR desc170(.Q(acs_prob_tdata_54[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  FDR desc171(.Q(acs_prob_tdata_54[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  FDR desc172(.Q(acs_prob_tdata_54[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11));
  p_O_FD desc173(.Q(acs_prob_tdata_54[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc173_p_O_FD));
  p_O_FD desc174(.Q(acs_prob_tdata_54[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc174_p_O_FD));
  LUT6 desc175(.I0(un4_v_high_s_7_1),.I1(un4_v_low_s_7_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMEM11),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc175.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc176(.I0(un4_v_high_s_8_1),.I1(un4_v_low_s_8_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMEM11),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc176.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc177(.I0(un4_v_high_s_6_1),.I1(un4_v_low_s_6_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc177.INIT=32'hACACFF00;
  LUT5 desc178(.I0(un4_v_high_s_5_1),.I1(un4_v_low_s_5_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc178.INIT=32'hACACFF00;
  LUT5 desc179(.I0(un4_v_high_s_4_1),.I1(un4_v_low_s_4_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc179.INIT=32'hACACFF00;
  LUT5 desc180(.I0(un4_v_high_s_3_1),.I1(un4_v_low_s_3_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc180.INIT=32'hACACFF00;
  LUT5 desc181(.I0(un4_v_high_s_2_1),.I1(un4_v_low_s_2_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc181.INIT=32'hACACFF00;
  LUT5 desc182(.I0(un4_v_high_s_1_1),.I1(un4_v_low_s_1_1),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_54[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc182.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[54:54]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc183(.I0(acs_prob_tdata_44[0:0]),.I1(acs_prob_tdata_45[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc183.INIT=16'h9669;
  LUT2 desc184(.I0(un4_v_high_s_1_1),.I1(un4_v_low_s_1_1),.O(v_diff_1_axb_1));
defparam desc184.INIT=4'h9;
  LUT2 desc185(.I0(un4_v_high_s_2_1),.I1(un4_v_low_s_2_1),.O(v_diff_1_axb_2));
defparam desc185.INIT=4'h9;
  LUT2 desc186(.I0(un4_v_high_s_3_1),.I1(un4_v_low_s_3_1),.O(v_diff_1_axb_3));
defparam desc186.INIT=4'h9;
  LUT2 desc187(.I0(un4_v_high_s_4_1),.I1(un4_v_low_s_4_1),.O(v_diff_1_axb_4));
defparam desc187.INIT=4'h9;
  LUT2 desc188(.I0(un4_v_high_s_5_1),.I1(un4_v_low_s_5_1),.O(v_diff_1_axb_5));
defparam desc188.INIT=4'h9;
  LUT2 desc189(.I0(un4_v_high_s_6_1),.I1(un4_v_low_s_6_1),.O(v_diff_1_axb_6));
defparam desc189.INIT=4'h9;
  LUT2 desc190(.I0(un4_v_high_s_7_1),.I1(un4_v_low_s_7_1),.O(v_diff_1_axb_7));
defparam desc190.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_44[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_44[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_44[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_44[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_44[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_44[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_44[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_45[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_45[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_45[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_45[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_45[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_45[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_45[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_45[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc191(.I0(acs_prob_tdata_44[0:0]),.I1(acs_prob_tdata_45[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2328));
defparam desc191.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_45[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_44[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc192(.I0(un4_v_high_s_8_1),.I1(un4_v_low_s_8_1),.O(v_diff_1_axb_8));
defparam desc192.INIT=4'h9;
  LUT6 desc193(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc193.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI4CHU(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI4CHU.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIMEM11_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIMEM11));
defparam s_axis_inbranch_tlast_d_RNIMEM11_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_44[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIKV121_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_1));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_1));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_45[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_1));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_45[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_1));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_45[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_1));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_45[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_1));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_45[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_1));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_45[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_1));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_45[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_45[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_1));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_1));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_44[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_1));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_44[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_1));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_44[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_1));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_44[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_1));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_44[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_1));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_44[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_1));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_44[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_44[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc194(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc195(.DI(un4_v_low_s_7_1),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc196(.DI(un4_v_low_s_6_1),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc197(.DI(un4_v_low_s_5_1),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc198(.DI(un4_v_low_s_4_1),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc199(.DI(un4_v_low_s_3_1),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc200(.DI(un4_v_low_s_2_1),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc201(.DI(un4_v_low_s_1_1),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc202(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc203(.Q(acs_prob_tdata_54[0:0]),.D(N_2328),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMEM11),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc203_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc204(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIKV121_O6));
defparam desc204.INIT=16'hF4F0;
  LUT2 desc205(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc205.INIT=4'h8;
endmodule
module acsZ0_3_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_21,acs_prob_tdata_20,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_42,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc212_p_O_FD,p_desc213_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc242_p_O_FDRE);
input branch_tlast ;
output [42:42] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_21 ;
input [8:0] acs_prob_tdata_20 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_42 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIBQC91_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIG3A81 ;
wire un4_v_high_s_7_2 ;
wire un4_v_low_s_7_2 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_2 ;
wire un4_v_low_s_8_2 ;
wire un4_v_high_s_6_2 ;
wire un4_v_low_s_6_2 ;
wire un4_v_high_s_5_2 ;
wire un4_v_low_s_5_2 ;
wire un4_v_high_s_4_2 ;
wire un4_v_low_s_4_2 ;
wire un4_v_high_s_3_2 ;
wire un4_v_low_s_3_2 ;
wire un4_v_high_s_2_2 ;
wire un4_v_low_s_2_2 ;
wire un4_v_high_s_1_2 ;
wire un4_v_low_s_1_2 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2308 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc212_p_O_FD ;
input p_desc213_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc242_p_O_FDRE ;
// instances
  FDR desc206(.Q(acs_prob_tdata_42[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  FDR desc207(.Q(acs_prob_tdata_42[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  FDR desc208(.Q(acs_prob_tdata_42[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  FDR desc209(.Q(acs_prob_tdata_42[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  FDR desc210(.Q(acs_prob_tdata_42[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  FDR desc211(.Q(acs_prob_tdata_42[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81));
  p_O_FD desc212(.Q(acs_prob_tdata_42[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc212_p_O_FD));
  p_O_FD desc213(.Q(acs_prob_tdata_42[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc213_p_O_FD));
  LUT6 desc214(.I0(un4_v_high_s_7_2),.I1(un4_v_low_s_7_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG3A81),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc214.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc215(.I0(un4_v_high_s_8_2),.I1(un4_v_low_s_8_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG3A81),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc215.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc216(.I0(un4_v_high_s_6_2),.I1(un4_v_low_s_6_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc216.INIT=32'hACACFF00;
  LUT5 desc217(.I0(un4_v_high_s_5_2),.I1(un4_v_low_s_5_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc217.INIT=32'hACACFF00;
  LUT5 desc218(.I0(un4_v_high_s_4_2),.I1(un4_v_low_s_4_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc218.INIT=32'hACACFF00;
  LUT5 desc219(.I0(un4_v_high_s_3_2),.I1(un4_v_low_s_3_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc219.INIT=32'hACACFF00;
  LUT5 desc220(.I0(un4_v_high_s_2_2),.I1(un4_v_low_s_2_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc220.INIT=32'hACACFF00;
  LUT5 desc221(.I0(un4_v_high_s_1_2),.I1(un4_v_low_s_1_2),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_42[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc221.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[42:42]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc222(.I0(acs_prob_tdata_20[0:0]),.I1(acs_prob_tdata_21[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc222.INIT=16'h9669;
  LUT2 desc223(.I0(un4_v_high_s_1_2),.I1(un4_v_low_s_1_2),.O(v_diff_1_axb_1));
defparam desc223.INIT=4'h9;
  LUT2 desc224(.I0(un4_v_high_s_2_2),.I1(un4_v_low_s_2_2),.O(v_diff_1_axb_2));
defparam desc224.INIT=4'h9;
  LUT2 desc225(.I0(un4_v_high_s_3_2),.I1(un4_v_low_s_3_2),.O(v_diff_1_axb_3));
defparam desc225.INIT=4'h9;
  LUT2 desc226(.I0(un4_v_high_s_4_2),.I1(un4_v_low_s_4_2),.O(v_diff_1_axb_4));
defparam desc226.INIT=4'h9;
  LUT2 desc227(.I0(un4_v_high_s_5_2),.I1(un4_v_low_s_5_2),.O(v_diff_1_axb_5));
defparam desc227.INIT=4'h9;
  LUT2 desc228(.I0(un4_v_high_s_6_2),.I1(un4_v_low_s_6_2),.O(v_diff_1_axb_6));
defparam desc228.INIT=4'h9;
  LUT2 desc229(.I0(un4_v_high_s_7_2),.I1(un4_v_low_s_7_2),.O(v_diff_1_axb_7));
defparam desc229.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_20[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_20[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_20[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_20[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_20[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_20[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_20[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_21[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_21[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_21[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_21[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_21[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_21[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_21[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_21[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc230(.I0(acs_prob_tdata_20[0:0]),.I1(acs_prob_tdata_21[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2308));
defparam desc230.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_21[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_20[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc231(.I0(un4_v_high_s_8_2),.I1(un4_v_low_s_8_2),.O(v_diff_1_axb_8));
defparam desc231.INIT=4'h9;
  LUT6 desc232(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc232.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIU0551(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIU0551.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIG3A81_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIG3A81));
defparam s_axis_inbranch_tlast_d_RNIG3A81_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_20[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIBQC91_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_2));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_2));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_21[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_2));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_21[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_2));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_21[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_2));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_21[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_2));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_21[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_2));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_21[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_2));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_21[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_21[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_2));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_2));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_20[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_2));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_20[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_2));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_20[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_2));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_20[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_2));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_20[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_2));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_20[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_2));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_20[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_20[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc233(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc234(.DI(un4_v_low_s_7_2),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc235(.DI(un4_v_low_s_6_2),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc236(.DI(un4_v_low_s_5_2),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc237(.DI(un4_v_low_s_4_2),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc238(.DI(un4_v_low_s_3_2),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc239(.DI(un4_v_low_s_2_2),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc240(.DI(un4_v_low_s_1_2),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc241(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc242(.Q(acs_prob_tdata_42[0:0]),.D(N_2308),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG3A81),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc242_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc243(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIBQC91_O6));
defparam desc243.INIT=16'hF4F0;
  LUT2 desc244(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc244.INIT=4'h8;
endmodule
module acsZ0_4_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_49,acs_prob_tdata_48,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_24,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc251_p_O_FD,p_desc252_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc281_p_O_FDRE);
input branch_tlast ;
output [24:24] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_49 ;
input [8:0] acs_prob_tdata_48 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_24 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIBK0A1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIGV3I1 ;
wire un4_v_high_s_7_3 ;
wire un4_v_low_s_7_3 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_3 ;
wire un4_v_low_s_8_3 ;
wire un4_v_high_s_6_3 ;
wire un4_v_low_s_6_3 ;
wire un4_v_high_s_5_3 ;
wire un4_v_low_s_5_3 ;
wire un4_v_high_s_4_3 ;
wire un4_v_low_s_4_3 ;
wire un4_v_high_s_3_3 ;
wire un4_v_low_s_3_3 ;
wire un4_v_high_s_2_3 ;
wire un4_v_low_s_2_3 ;
wire un4_v_high_s_1_3 ;
wire un4_v_low_s_1_3 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2288 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc251_p_O_FD ;
input p_desc252_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc281_p_O_FDRE ;
// instances
  FDR desc245(.Q(acs_prob_tdata_24[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  FDR desc246(.Q(acs_prob_tdata_24[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  FDR desc247(.Q(acs_prob_tdata_24[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  FDR desc248(.Q(acs_prob_tdata_24[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  FDR desc249(.Q(acs_prob_tdata_24[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  FDR desc250(.Q(acs_prob_tdata_24[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1));
  p_O_FD desc251(.Q(acs_prob_tdata_24[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc251_p_O_FD));
  p_O_FD desc252(.Q(acs_prob_tdata_24[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc252_p_O_FD));
  LUT6 desc253(.I0(un4_v_high_s_7_3),.I1(un4_v_low_s_7_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGV3I1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc253.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc254(.I0(un4_v_high_s_8_3),.I1(un4_v_low_s_8_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGV3I1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc254.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc255(.I0(un4_v_high_s_6_3),.I1(un4_v_low_s_6_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc255.INIT=32'hACACFF00;
  LUT5 desc256(.I0(un4_v_high_s_5_3),.I1(un4_v_low_s_5_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc256.INIT=32'hACACFF00;
  LUT5 desc257(.I0(un4_v_high_s_4_3),.I1(un4_v_low_s_4_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc257.INIT=32'hACACFF00;
  LUT5 desc258(.I0(un4_v_high_s_3_3),.I1(un4_v_low_s_3_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc258.INIT=32'hACACFF00;
  LUT5 desc259(.I0(un4_v_high_s_2_3),.I1(un4_v_low_s_2_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc259.INIT=32'hACACFF00;
  LUT5 desc260(.I0(un4_v_high_s_1_3),.I1(un4_v_low_s_1_3),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_24[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc260.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[24:24]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc261(.I0(acs_prob_tdata_48[0:0]),.I1(acs_prob_tdata_49[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc261.INIT=16'h9669;
  LUT2 desc262(.I0(un4_v_high_s_1_3),.I1(un4_v_low_s_1_3),.O(v_diff_1_axb_1));
defparam desc262.INIT=4'h9;
  LUT2 desc263(.I0(un4_v_high_s_2_3),.I1(un4_v_low_s_2_3),.O(v_diff_1_axb_2));
defparam desc263.INIT=4'h9;
  LUT2 desc264(.I0(un4_v_high_s_3_3),.I1(un4_v_low_s_3_3),.O(v_diff_1_axb_3));
defparam desc264.INIT=4'h9;
  LUT2 desc265(.I0(un4_v_high_s_4_3),.I1(un4_v_low_s_4_3),.O(v_diff_1_axb_4));
defparam desc265.INIT=4'h9;
  LUT2 desc266(.I0(un4_v_high_s_5_3),.I1(un4_v_low_s_5_3),.O(v_diff_1_axb_5));
defparam desc266.INIT=4'h9;
  LUT2 desc267(.I0(un4_v_high_s_6_3),.I1(un4_v_low_s_6_3),.O(v_diff_1_axb_6));
defparam desc267.INIT=4'h9;
  LUT2 desc268(.I0(un4_v_high_s_7_3),.I1(un4_v_low_s_7_3),.O(v_diff_1_axb_7));
defparam desc268.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_48[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_48[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_48[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_48[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_48[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_48[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_48[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_49[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_49[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_49[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_49[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_49[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_49[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_49[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_49[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc269(.I0(acs_prob_tdata_48[0:0]),.I1(acs_prob_tdata_49[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2288));
defparam desc269.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_49[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_48[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc270(.I0(un4_v_high_s_8_3),.I1(un4_v_low_s_8_3),.O(v_diff_1_axb_8));
defparam desc270.INIT=4'h9;
  LUT6 desc271(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc271.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIUSUE1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIUSUE1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIGV3I1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIGV3I1));
defparam s_axis_inbranch_tlast_d_RNIGV3I1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_48[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIBK0A1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_3));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_3));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_49[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_3));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_49[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_3));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_49[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_3));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_49[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_3));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_49[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_3));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_49[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_3));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_49[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_49[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_3));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_3));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_48[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_3));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_48[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_3));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_48[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_3));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_48[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_3));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_48[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_3));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_48[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_3));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_48[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_48[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc272(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc273(.DI(un4_v_low_s_7_3),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc274(.DI(un4_v_low_s_6_3),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc275(.DI(un4_v_low_s_5_3),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc276(.DI(un4_v_low_s_4_3),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc277(.DI(un4_v_low_s_3_3),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc278(.DI(un4_v_low_s_2_3),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc279(.DI(un4_v_low_s_1_3),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc280(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc281(.Q(acs_prob_tdata_24[0:0]),.D(N_2288),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGV3I1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc281_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc282(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIBK0A1_O6));
defparam desc282.INIT=16'hF4F0;
  LUT2 desc283(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc283.INIT=4'h8;
endmodule
module acsZ0_5_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_51,acs_prob_tdata_50,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_25,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc290_p_O_FD,p_desc291_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc320_p_O_FDRE);
input branch_tlast ;
output [25:25] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_51 ;
input [8:0] acs_prob_tdata_50 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_25 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIEA0T_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNII2741 ;
wire un4_v_high_s_7_4 ;
wire un4_v_low_s_7_4 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_4 ;
wire un4_v_low_s_8_4 ;
wire un4_v_high_s_6_4 ;
wire un4_v_low_s_6_4 ;
wire un4_v_high_s_5_4 ;
wire un4_v_low_s_5_4 ;
wire un4_v_high_s_4_4 ;
wire un4_v_low_s_4_4 ;
wire un4_v_high_s_3_4 ;
wire un4_v_low_s_3_4 ;
wire un4_v_high_s_2_4 ;
wire un4_v_low_s_2_4 ;
wire un4_v_high_s_1_4 ;
wire un4_v_low_s_1_4 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2268 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc290_p_O_FD ;
input p_desc291_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc320_p_O_FDRE ;
// instances
  FDR desc284(.Q(acs_prob_tdata_25[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  FDR desc285(.Q(acs_prob_tdata_25[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  FDR desc286(.Q(acs_prob_tdata_25[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  FDR desc287(.Q(acs_prob_tdata_25[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  FDR desc288(.Q(acs_prob_tdata_25[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  FDR desc289(.Q(acs_prob_tdata_25[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741));
  p_O_FD desc290(.Q(acs_prob_tdata_25[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc290_p_O_FD));
  p_O_FD desc291(.Q(acs_prob_tdata_25[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc291_p_O_FD));
  LUT6 desc292(.I0(un4_v_high_s_7_4),.I1(un4_v_low_s_7_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII2741),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc292.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc293(.I0(un4_v_high_s_8_4),.I1(un4_v_low_s_8_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII2741),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc293.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc294(.I0(un4_v_high_s_6_4),.I1(un4_v_low_s_6_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc294.INIT=32'hACACFF00;
  LUT5 desc295(.I0(un4_v_high_s_5_4),.I1(un4_v_low_s_5_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc295.INIT=32'hACACFF00;
  LUT5 desc296(.I0(un4_v_high_s_4_4),.I1(un4_v_low_s_4_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc296.INIT=32'hACACFF00;
  LUT5 desc297(.I0(un4_v_high_s_3_4),.I1(un4_v_low_s_3_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc297.INIT=32'hACACFF00;
  LUT5 desc298(.I0(un4_v_high_s_2_4),.I1(un4_v_low_s_2_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc298.INIT=32'hACACFF00;
  LUT5 desc299(.I0(un4_v_high_s_1_4),.I1(un4_v_low_s_1_4),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_25[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc299.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[25:25]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc300(.I0(acs_prob_tdata_50[0:0]),.I1(acs_prob_tdata_51[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc300.INIT=16'h9669;
  LUT2 desc301(.I0(un4_v_high_s_1_4),.I1(un4_v_low_s_1_4),.O(v_diff_1_axb_1));
defparam desc301.INIT=4'h9;
  LUT2 desc302(.I0(un4_v_high_s_2_4),.I1(un4_v_low_s_2_4),.O(v_diff_1_axb_2));
defparam desc302.INIT=4'h9;
  LUT2 desc303(.I0(un4_v_high_s_3_4),.I1(un4_v_low_s_3_4),.O(v_diff_1_axb_3));
defparam desc303.INIT=4'h9;
  LUT2 desc304(.I0(un4_v_high_s_4_4),.I1(un4_v_low_s_4_4),.O(v_diff_1_axb_4));
defparam desc304.INIT=4'h9;
  LUT2 desc305(.I0(un4_v_high_s_5_4),.I1(un4_v_low_s_5_4),.O(v_diff_1_axb_5));
defparam desc305.INIT=4'h9;
  LUT2 desc306(.I0(un4_v_high_s_6_4),.I1(un4_v_low_s_6_4),.O(v_diff_1_axb_6));
defparam desc306.INIT=4'h9;
  LUT2 desc307(.I0(un4_v_high_s_7_4),.I1(un4_v_low_s_7_4),.O(v_diff_1_axb_7));
defparam desc307.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_50[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_50[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_50[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_50[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_50[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_50[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_50[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_51[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_51[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_51[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_51[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_51[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_51[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_51[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_51[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc308(.I0(acs_prob_tdata_50[0:0]),.I1(acs_prob_tdata_51[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2268));
defparam desc308.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_51[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_50[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc309(.I0(un4_v_high_s_8_4),.I1(un4_v_low_s_8_4),.O(v_diff_1_axb_8));
defparam desc309.INIT=4'h9;
  LUT6 desc310(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc310.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI00211(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI00211.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNII2741_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNII2741));
defparam s_axis_inbranch_tlast_d_RNII2741_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_50[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIEA0T_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_4));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_4));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_51[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_4));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_51[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_4));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_51[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_4));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_51[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_4));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_51[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_4));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_51[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_4));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_51[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_51[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_4));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_4));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_50[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_4));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_50[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_4));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_50[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_4));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_50[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_4));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_50[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_4));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_50[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_4));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_50[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_50[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc311(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc312(.DI(un4_v_low_s_7_4),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc313(.DI(un4_v_low_s_6_4),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc314(.DI(un4_v_low_s_5_4),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc315(.DI(un4_v_low_s_4_4),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc316(.DI(un4_v_low_s_3_4),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc317(.DI(un4_v_low_s_2_4),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc318(.DI(un4_v_low_s_1_4),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc319(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc320(.Q(acs_prob_tdata_25[0:0]),.D(N_2268),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII2741),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc320_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc321(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIEA0T_O6));
defparam desc321.INIT=16'hF4F0;
  LUT2 desc322(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc322.INIT=4'h8;
endmodule
module acsZ0_6_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_33,acs_prob_tdata_32,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_16,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc329_p_O_FD,p_desc330_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc359_p_O_FDRE);
input branch_tlast ;
output [16:16] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_33 ;
input [8:0] acs_prob_tdata_32 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_16 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIE7AD1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNII04H1 ;
wire un4_v_high_s_7_5 ;
wire un4_v_low_s_7_5 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_5 ;
wire un4_v_low_s_8_5 ;
wire un4_v_high_s_6_5 ;
wire un4_v_low_s_6_5 ;
wire un4_v_high_s_5_5 ;
wire un4_v_low_s_5_5 ;
wire un4_v_high_s_4_5 ;
wire un4_v_low_s_4_5 ;
wire un4_v_high_s_3_5 ;
wire un4_v_low_s_3_5 ;
wire un4_v_high_s_2_5 ;
wire un4_v_low_s_2_5 ;
wire un4_v_high_s_1_5 ;
wire un4_v_low_s_1_5 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_2248 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc329_p_O_FD ;
input p_desc330_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc359_p_O_FDRE ;
// instances
  FDR desc323(.Q(acs_prob_tdata_16[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  FDR desc324(.Q(acs_prob_tdata_16[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  FDR desc325(.Q(acs_prob_tdata_16[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  FDR desc326(.Q(acs_prob_tdata_16[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  FDR desc327(.Q(acs_prob_tdata_16[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  FDR desc328(.Q(acs_prob_tdata_16[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1));
  p_O_FD desc329(.Q(acs_prob_tdata_16[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc329_p_O_FD));
  p_O_FD desc330(.Q(acs_prob_tdata_16[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc330_p_O_FD));
  LUT6 desc331(.I0(un4_v_high_s_7_5),.I1(un4_v_low_s_7_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII04H1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc331.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc332(.I0(un4_v_high_s_8_5),.I1(un4_v_low_s_8_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII04H1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc332.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc333(.I0(un4_v_high_s_6_5),.I1(un4_v_low_s_6_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc333.INIT=32'hACACFF00;
  LUT5 desc334(.I0(un4_v_high_s_5_5),.I1(un4_v_low_s_5_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc334.INIT=32'hACACFF00;
  LUT5 desc335(.I0(un4_v_high_s_4_5),.I1(un4_v_low_s_4_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc335.INIT=32'hACACFF00;
  LUT5 desc336(.I0(un4_v_high_s_3_5),.I1(un4_v_low_s_3_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc336.INIT=32'hACACFF00;
  LUT5 desc337(.I0(un4_v_high_s_2_5),.I1(un4_v_low_s_2_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc337.INIT=32'hACACFF00;
  LUT5 desc338(.I0(un4_v_high_s_1_5),.I1(un4_v_low_s_1_5),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_16[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc338.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[16:16]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_32[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_32[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_32[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_32[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_32[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_32[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_32[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_33[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_33[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_33[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_33[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_33[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_33[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_33[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_33[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc339(.I0(acs_prob_tdata_32[0:0]),.I1(acs_prob_tdata_33[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc339.INIT=16'h9669;
  LUT2 desc340(.I0(un4_v_high_s_1_5),.I1(un4_v_low_s_1_5),.O(v_diff_1_axb_1));
defparam desc340.INIT=4'h9;
  LUT2 desc341(.I0(un4_v_high_s_2_5),.I1(un4_v_low_s_2_5),.O(v_diff_1_axb_2));
defparam desc341.INIT=4'h9;
  LUT2 desc342(.I0(un4_v_high_s_3_5),.I1(un4_v_low_s_3_5),.O(v_diff_1_axb_3));
defparam desc342.INIT=4'h9;
  LUT2 desc343(.I0(un4_v_high_s_4_5),.I1(un4_v_low_s_4_5),.O(v_diff_1_axb_4));
defparam desc343.INIT=4'h9;
  LUT2 desc344(.I0(un4_v_high_s_5_5),.I1(un4_v_low_s_5_5),.O(v_diff_1_axb_5));
defparam desc344.INIT=4'h9;
  LUT2 desc345(.I0(un4_v_high_s_6_5),.I1(un4_v_low_s_6_5),.O(v_diff_1_axb_6));
defparam desc345.INIT=4'h9;
  LUT2 desc346(.I0(un4_v_high_s_7_5),.I1(un4_v_low_s_7_5),.O(v_diff_1_axb_7));
defparam desc346.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc347(.I0(acs_prob_tdata_32[0:0]),.I1(acs_prob_tdata_33[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2248));
defparam desc347.INIT=32'h3C3C55AA;
  LUT2 desc348(.I0(un4_v_high_s_8_5),.I1(un4_v_low_s_8_5),.O(v_diff_1_axb_8));
defparam desc348.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_33[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_32[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc349(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc349.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI0UUD1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI0UUD1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNII04H1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNII04H1));
defparam s_axis_inbranch_tlast_d_RNII04H1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_32[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIE7AD1_O6),.C(aclk),.R(aresetn_i));
  XORCY desc350(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc351(.DI(un4_v_low_s_7_5),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc352(.DI(un4_v_low_s_6_5),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc353(.DI(un4_v_low_s_5_5),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc354(.DI(un4_v_low_s_4_5),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc355(.DI(un4_v_low_s_3_5),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc356(.DI(un4_v_low_s_2_5),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc357(.DI(un4_v_low_s_1_5),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc358(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_5));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_5));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_33[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_5));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_33[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_5));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_33[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_5));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_33[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_5));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_33[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_5));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_33[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_5));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_33[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_33[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_5));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_5));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_32[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_5));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_32[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_5));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_32[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_5));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_32[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_5));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_32[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_5));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_32[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_5));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_32[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_32[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc359(.Q(acs_prob_tdata_16[0:0]),.D(N_2248),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII04H1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc359_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc360(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIE7AD1_O6));
defparam desc360.INIT=16'hF4F0;
  LUT2 desc361(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc361.INIT=4'h8;
endmodule
module acsZ0_7_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_3,acs_prob_tdata_2,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_1,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_4_rep1,N_1756_1,aresetn,p_desc368_p_O_FD,p_desc369_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc398_p_O_FDRE);
input branch_tlast ;
output [1:1] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_3 ;
input [8:0] acs_prob_tdata_2 ;
input [1:0] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_1 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNICHF11_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI6TE71 ;
wire un4_v_high_s_7_6 ;
wire un4_v_low_s_7_6 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_6 ;
wire un4_v_low_s_8_6 ;
wire un4_v_high_s_6_6 ;
wire un4_v_low_s_6_6 ;
wire un4_v_high_s_5_6 ;
wire un4_v_low_s_5_6 ;
wire un4_v_high_s_4_6 ;
wire un4_v_low_s_4_6 ;
wire un4_v_high_s_3_6 ;
wire un4_v_low_s_3_6 ;
wire un4_v_high_s_2_6 ;
wire un4_v_low_s_2_6 ;
wire un4_v_high_s_1_6 ;
wire un4_v_low_s_1_6 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_2228 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc368_p_O_FD ;
input p_desc369_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc398_p_O_FDRE ;
// instances
  FDR desc362(.Q(acs_prob_tdata_1[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  FDR desc363(.Q(acs_prob_tdata_1[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  FDR desc364(.Q(acs_prob_tdata_1[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  FDR desc365(.Q(acs_prob_tdata_1[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  FDR desc366(.Q(acs_prob_tdata_1[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  FDR desc367(.Q(acs_prob_tdata_1[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71));
  p_O_FD desc368(.Q(acs_prob_tdata_1[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc368_p_O_FD));
  p_O_FD desc369(.Q(acs_prob_tdata_1[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc369_p_O_FD));
  LUT6 desc370(.I0(un4_v_high_s_7_6),.I1(un4_v_low_s_7_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI6TE71),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc370.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc371(.I0(un4_v_high_s_8_6),.I1(un4_v_low_s_8_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI6TE71),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc371.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc372(.I0(un4_v_high_s_6_6),.I1(un4_v_low_s_6_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc372.INIT=32'hACACFF00;
  LUT5 desc373(.I0(un4_v_high_s_5_6),.I1(un4_v_low_s_5_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc373.INIT=32'hACACFF00;
  LUT5 desc374(.I0(un4_v_high_s_4_6),.I1(un4_v_low_s_4_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc374.INIT=32'hACACFF00;
  LUT5 desc375(.I0(un4_v_high_s_3_6),.I1(un4_v_low_s_3_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc375.INIT=32'hACACFF00;
  LUT5 desc376(.I0(un4_v_high_s_2_6),.I1(un4_v_low_s_2_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc376.INIT=32'hACACFF00;
  LUT5 desc377(.I0(un4_v_high_s_1_6),.I1(un4_v_low_s_1_6),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_1[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc377.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[1:1]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_2[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_2[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_2[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_2[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_2[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_2[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_2[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_3[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_3[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_3[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_3[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_3[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_3[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_3[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_3[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc378(.I0(acs_prob_tdata_2[0:0]),.I1(acs_prob_tdata_3[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc378.INIT=16'h9669;
  LUT2 desc379(.I0(un4_v_high_s_1_6),.I1(un4_v_low_s_1_6),.O(v_diff_1_axb_1));
defparam desc379.INIT=4'h9;
  LUT2 desc380(.I0(un4_v_high_s_2_6),.I1(un4_v_low_s_2_6),.O(v_diff_1_axb_2));
defparam desc380.INIT=4'h9;
  LUT2 desc381(.I0(un4_v_high_s_3_6),.I1(un4_v_low_s_3_6),.O(v_diff_1_axb_3));
defparam desc381.INIT=4'h9;
  LUT2 desc382(.I0(un4_v_high_s_4_6),.I1(un4_v_low_s_4_6),.O(v_diff_1_axb_4));
defparam desc382.INIT=4'h9;
  LUT2 desc383(.I0(un4_v_high_s_5_6),.I1(un4_v_low_s_5_6),.O(v_diff_1_axb_5));
defparam desc383.INIT=4'h9;
  LUT2 desc384(.I0(un4_v_high_s_6_6),.I1(un4_v_low_s_6_6),.O(v_diff_1_axb_6));
defparam desc384.INIT=4'h9;
  LUT2 desc385(.I0(un4_v_high_s_7_6),.I1(un4_v_low_s_7_6),.O(v_diff_1_axb_7));
defparam desc385.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc386(.I0(acs_prob_tdata_2[0:0]),.I1(acs_prob_tdata_3[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2228));
defparam desc386.INIT=32'h33CC5A5A;
  LUT2 desc387(.I0(un4_v_high_s_8_6),.I1(un4_v_low_s_8_6),.O(v_diff_1_axb_8));
defparam desc387.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_3[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_2[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc388(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4_rep1),.I2(write_ram_fsm[0:0]),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc388.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIKQ941(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIKQ941.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI6TE71_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI6TE71));
defparam s_axis_inbranch_tlast_d_RNI6TE71_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_2[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNICHF11_O6),.C(aclk),.R(aresetn_i));
  XORCY desc389(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc390(.DI(un4_v_low_s_7_6),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc391(.DI(un4_v_low_s_6_6),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc392(.DI(un4_v_low_s_5_6),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc393(.DI(un4_v_low_s_4_6),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc394(.DI(un4_v_low_s_3_6),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc395(.DI(un4_v_low_s_2_6),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc396(.DI(un4_v_low_s_1_6),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc397(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_6));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_6));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_3[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_6));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_3[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_6));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_3[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_6));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_3[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_6));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_3[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_6));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_3[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_6));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_3[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_3[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_6));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_6));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_2[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_6));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_2[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_6));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_2[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_6));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_2[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_6));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_2[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_6));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_2[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_6));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_2[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_2[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc398(.Q(acs_prob_tdata_1[0:0]),.D(N_2228),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6TE71),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc398_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc399(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNICHF11_O6));
defparam desc399.INIT=16'hF4F0;
  LUT2 desc400(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc400.INIT=4'h8;
endmodule
module acsZ0_8_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_3,acs_prob_tdata_2,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_33,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc407_p_O_FD,p_desc408_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc437_p_O_FDRE);
input branch_tlast ;
output [33:33] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_3 ;
input [8:0] acs_prob_tdata_2 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_33 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIBNMP_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIG1751 ;
wire un4_v_high_s_7_7 ;
wire un4_v_low_s_7_7 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_7 ;
wire un4_v_low_s_8_7 ;
wire un4_v_high_s_6_7 ;
wire un4_v_low_s_6_7 ;
wire un4_v_high_s_5_7 ;
wire un4_v_low_s_5_7 ;
wire un4_v_high_s_4_7 ;
wire un4_v_low_s_4_7 ;
wire un4_v_high_s_3_7 ;
wire un4_v_low_s_3_7 ;
wire un4_v_high_s_2_7 ;
wire un4_v_low_s_2_7 ;
wire un4_v_high_s_1_7 ;
wire un4_v_low_s_1_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2208 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc407_p_O_FD ;
input p_desc408_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc437_p_O_FDRE ;
// instances
  FDR desc401(.Q(acs_prob_tdata_33[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  FDR desc402(.Q(acs_prob_tdata_33[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  FDR desc403(.Q(acs_prob_tdata_33[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  FDR desc404(.Q(acs_prob_tdata_33[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  FDR desc405(.Q(acs_prob_tdata_33[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  FDR desc406(.Q(acs_prob_tdata_33[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751));
  p_O_FD desc407(.Q(acs_prob_tdata_33[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc407_p_O_FD));
  p_O_FD desc408(.Q(acs_prob_tdata_33[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc408_p_O_FD));
  LUT6 desc409(.I0(un4_v_high_s_7_7),.I1(un4_v_low_s_7_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG1751),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc409.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc410(.I0(un4_v_high_s_8_7),.I1(un4_v_low_s_8_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG1751),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc410.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc411(.I0(un4_v_high_s_6_7),.I1(un4_v_low_s_6_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc411.INIT=32'hACACFF00;
  LUT5 desc412(.I0(un4_v_high_s_5_7),.I1(un4_v_low_s_5_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc412.INIT=32'hACACFF00;
  LUT5 desc413(.I0(un4_v_high_s_4_7),.I1(un4_v_low_s_4_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc413.INIT=32'hACACFF00;
  LUT5 desc414(.I0(un4_v_high_s_3_7),.I1(un4_v_low_s_3_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc414.INIT=32'hACACFF00;
  LUT5 desc415(.I0(un4_v_high_s_2_7),.I1(un4_v_low_s_2_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc415.INIT=32'hACACFF00;
  LUT5 desc416(.I0(un4_v_high_s_1_7),.I1(un4_v_low_s_1_7),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_33[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc416.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[33:33]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc417(.I0(acs_prob_tdata_2[0:0]),.I1(acs_prob_tdata_3[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc417.INIT=16'h9669;
  LUT2 desc418(.I0(un4_v_high_s_1_7),.I1(un4_v_low_s_1_7),.O(v_diff_1_axb_1));
defparam desc418.INIT=4'h9;
  LUT2 desc419(.I0(un4_v_high_s_2_7),.I1(un4_v_low_s_2_7),.O(v_diff_1_axb_2));
defparam desc419.INIT=4'h9;
  LUT2 desc420(.I0(un4_v_high_s_3_7),.I1(un4_v_low_s_3_7),.O(v_diff_1_axb_3));
defparam desc420.INIT=4'h9;
  LUT2 desc421(.I0(un4_v_high_s_4_7),.I1(un4_v_low_s_4_7),.O(v_diff_1_axb_4));
defparam desc421.INIT=4'h9;
  LUT2 desc422(.I0(un4_v_high_s_5_7),.I1(un4_v_low_s_5_7),.O(v_diff_1_axb_5));
defparam desc422.INIT=4'h9;
  LUT2 desc423(.I0(un4_v_high_s_6_7),.I1(un4_v_low_s_6_7),.O(v_diff_1_axb_6));
defparam desc423.INIT=4'h9;
  LUT2 desc424(.I0(un4_v_high_s_7_7),.I1(un4_v_low_s_7_7),.O(v_diff_1_axb_7));
defparam desc424.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_2[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_2[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_2[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_2[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_2[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_2[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_2[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_3[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_3[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_3[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_3[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_3[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_3[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_3[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_3[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc425(.I0(acs_prob_tdata_2[0:0]),.I1(acs_prob_tdata_3[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2208));
defparam desc425.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_3[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_2[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc426(.I0(un4_v_high_s_8_7),.I1(un4_v_low_s_8_7),.O(v_diff_1_axb_8));
defparam desc426.INIT=4'h9;
  LUT6 desc427(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc427.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIUU121(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIUU121.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIG1751_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIG1751));
defparam s_axis_inbranch_tlast_d_RNIG1751_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_2[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIBNMP_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_7));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_7));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_3[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_7));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_3[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_7));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_3[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_7));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_3[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_7));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_3[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_7));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_3[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_7));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_3[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_3[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_7));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_7));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_2[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_7));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_2[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_7));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_2[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_7));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_2[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_7));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_2[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_7));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_2[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_7));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_2[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_2[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc428(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc429(.DI(un4_v_low_s_7_7),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc430(.DI(un4_v_low_s_6_7),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc431(.DI(un4_v_low_s_5_7),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc432(.DI(un4_v_low_s_4_7),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc433(.DI(un4_v_low_s_3_7),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc434(.DI(un4_v_low_s_2_7),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc435(.DI(un4_v_low_s_1_7),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc436(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc437(.Q(acs_prob_tdata_33[0:0]),.D(N_2208),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG1751),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc437_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc438(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIBNMP_O6));
defparam desc438.INIT=16'hF4F0;
  LUT2 desc439(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc439.INIT=4'h8;
endmodule
module acsZ0_9_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_37,acs_prob_tdata_36,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_18,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc446_p_O_FD,p_desc447_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc476_p_O_FDRE);
input branch_tlast ;
output [18:18] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_37 ;
input [8:0] acs_prob_tdata_36 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_18 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIKJ931_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIM6A51 ;
wire un4_v_high_s_7_8 ;
wire un4_v_low_s_7_8 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_8 ;
wire un4_v_low_s_8_8 ;
wire un4_v_high_s_6_8 ;
wire un4_v_low_s_6_8 ;
wire un4_v_high_s_5_8 ;
wire un4_v_low_s_5_8 ;
wire un4_v_high_s_4_8 ;
wire un4_v_low_s_4_8 ;
wire un4_v_high_s_3_8 ;
wire un4_v_low_s_3_8 ;
wire un4_v_high_s_2_8 ;
wire un4_v_low_s_2_8 ;
wire un4_v_high_s_1_8 ;
wire un4_v_low_s_1_8 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2188 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc446_p_O_FD ;
input p_desc447_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc476_p_O_FDRE ;
// instances
  FDR desc440(.Q(acs_prob_tdata_18[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  FDR desc441(.Q(acs_prob_tdata_18[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  FDR desc442(.Q(acs_prob_tdata_18[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  FDR desc443(.Q(acs_prob_tdata_18[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  FDR desc444(.Q(acs_prob_tdata_18[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  FDR desc445(.Q(acs_prob_tdata_18[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51));
  p_O_FD desc446(.Q(acs_prob_tdata_18[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc446_p_O_FD));
  p_O_FD desc447(.Q(acs_prob_tdata_18[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc447_p_O_FD));
  LUT6 desc448(.I0(un4_v_high_s_7_8),.I1(un4_v_low_s_7_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIM6A51),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc448.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc449(.I0(un4_v_high_s_8_8),.I1(un4_v_low_s_8_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIM6A51),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc449.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc450(.I0(un4_v_high_s_6_8),.I1(un4_v_low_s_6_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc450.INIT=32'hACACFF00;
  LUT5 desc451(.I0(un4_v_high_s_5_8),.I1(un4_v_low_s_5_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc451.INIT=32'hACACFF00;
  LUT5 desc452(.I0(un4_v_high_s_4_8),.I1(un4_v_low_s_4_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc452.INIT=32'hACACFF00;
  LUT5 desc453(.I0(un4_v_high_s_3_8),.I1(un4_v_low_s_3_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc453.INIT=32'hACACFF00;
  LUT5 desc454(.I0(un4_v_high_s_2_8),.I1(un4_v_low_s_2_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc454.INIT=32'hACACFF00;
  LUT5 desc455(.I0(un4_v_high_s_1_8),.I1(un4_v_low_s_1_8),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_18[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc455.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[18:18]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc456(.I0(acs_prob_tdata_36[0:0]),.I1(acs_prob_tdata_37[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc456.INIT=16'h9669;
  LUT2 desc457(.I0(un4_v_high_s_1_8),.I1(un4_v_low_s_1_8),.O(v_diff_1_axb_1));
defparam desc457.INIT=4'h9;
  LUT2 desc458(.I0(un4_v_high_s_2_8),.I1(un4_v_low_s_2_8),.O(v_diff_1_axb_2));
defparam desc458.INIT=4'h9;
  LUT2 desc459(.I0(un4_v_high_s_3_8),.I1(un4_v_low_s_3_8),.O(v_diff_1_axb_3));
defparam desc459.INIT=4'h9;
  LUT2 desc460(.I0(un4_v_high_s_4_8),.I1(un4_v_low_s_4_8),.O(v_diff_1_axb_4));
defparam desc460.INIT=4'h9;
  LUT2 desc461(.I0(un4_v_high_s_5_8),.I1(un4_v_low_s_5_8),.O(v_diff_1_axb_5));
defparam desc461.INIT=4'h9;
  LUT2 desc462(.I0(un4_v_high_s_6_8),.I1(un4_v_low_s_6_8),.O(v_diff_1_axb_6));
defparam desc462.INIT=4'h9;
  LUT2 desc463(.I0(un4_v_high_s_7_8),.I1(un4_v_low_s_7_8),.O(v_diff_1_axb_7));
defparam desc463.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_36[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_36[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_36[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_36[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_36[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_36[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_36[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_37[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_37[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_37[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_37[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_37[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_37[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_37[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_37[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc464(.I0(acs_prob_tdata_36[0:0]),.I1(acs_prob_tdata_37[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2188));
defparam desc464.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_37[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_36[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc465(.I0(un4_v_high_s_8_8),.I1(un4_v_low_s_8_8),.O(v_diff_1_axb_8));
defparam desc465.INIT=4'h9;
  LUT6 desc466(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc466.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI44521(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI44521.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIM6A51_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIM6A51));
defparam s_axis_inbranch_tlast_d_RNIM6A51_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_36[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIKJ931_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_8));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_8));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_37[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_8));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_37[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_8));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_37[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_8));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_37[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_8));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_37[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_8));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_37[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_8));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_37[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_37[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_8));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_8));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_36[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_8));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_36[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_8));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_36[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_8));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_36[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_8));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_36[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_8));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_36[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_8));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_36[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_36[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc467(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc468(.DI(un4_v_low_s_7_8),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc469(.DI(un4_v_low_s_6_8),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc470(.DI(un4_v_low_s_5_8),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc471(.DI(un4_v_low_s_4_8),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc472(.DI(un4_v_low_s_3_8),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc473(.DI(un4_v_low_s_2_8),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc474(.DI(un4_v_low_s_1_8),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc475(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc476(.Q(acs_prob_tdata_18[0:0]),.D(N_2188),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM6A51),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc476_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc477(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIKJ931_O6));
defparam desc477.INIT=16'hF4F0;
  LUT2 desc478(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc478.INIT=4'h8;
endmodule
module acsZ0_10_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_7,acs_prob_tdata_6,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_3,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_4_rep1,N_1756_1,aresetn,p_desc485_p_O_FD,p_desc486_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc515_p_O_FDRE);
input branch_tlast ;
output [3:3] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_7 ;
input [8:0] acs_prob_tdata_6 ;
input [1:0] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_3 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIITE71_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIA3LB1 ;
wire un4_v_high_s_7_9 ;
wire un4_v_low_s_7_9 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_9 ;
wire un4_v_low_s_8_9 ;
wire un4_v_high_s_6_9 ;
wire un4_v_low_s_6_9 ;
wire un4_v_high_s_5_9 ;
wire un4_v_low_s_5_9 ;
wire un4_v_high_s_4_9 ;
wire un4_v_low_s_4_9 ;
wire un4_v_high_s_3_9 ;
wire un4_v_low_s_3_9 ;
wire un4_v_high_s_2_9 ;
wire un4_v_low_s_2_9 ;
wire un4_v_high_s_1_9 ;
wire un4_v_low_s_1_9 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2168 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc485_p_O_FD ;
input p_desc486_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc515_p_O_FDRE ;
// instances
  FDR desc479(.Q(acs_prob_tdata_3[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  FDR desc480(.Q(acs_prob_tdata_3[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  FDR desc481(.Q(acs_prob_tdata_3[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  FDR desc482(.Q(acs_prob_tdata_3[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  FDR desc483(.Q(acs_prob_tdata_3[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  FDR desc484(.Q(acs_prob_tdata_3[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1));
  p_O_FD desc485(.Q(acs_prob_tdata_3[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc485_p_O_FD));
  p_O_FD desc486(.Q(acs_prob_tdata_3[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc486_p_O_FD));
  LUT6 desc487(.I0(un4_v_high_s_7_9),.I1(un4_v_low_s_7_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIA3LB1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc487.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc488(.I0(un4_v_high_s_8_9),.I1(un4_v_low_s_8_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIA3LB1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc488.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc489(.I0(un4_v_high_s_6_9),.I1(un4_v_low_s_6_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc489.INIT=32'hACACFF00;
  LUT5 desc490(.I0(un4_v_high_s_5_9),.I1(un4_v_low_s_5_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc490.INIT=32'hACACFF00;
  LUT5 desc491(.I0(un4_v_high_s_4_9),.I1(un4_v_low_s_4_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc491.INIT=32'hACACFF00;
  LUT5 desc492(.I0(un4_v_high_s_3_9),.I1(un4_v_low_s_3_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc492.INIT=32'hACACFF00;
  LUT5 desc493(.I0(un4_v_high_s_2_9),.I1(un4_v_low_s_2_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc493.INIT=32'hACACFF00;
  LUT5 desc494(.I0(un4_v_high_s_1_9),.I1(un4_v_low_s_1_9),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_3[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc494.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[3:3]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc495(.I0(acs_prob_tdata_6[0:0]),.I1(acs_prob_tdata_7[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc495.INIT=16'h9669;
  LUT2 desc496(.I0(un4_v_high_s_1_9),.I1(un4_v_low_s_1_9),.O(v_diff_1_axb_1));
defparam desc496.INIT=4'h9;
  LUT2 desc497(.I0(un4_v_high_s_2_9),.I1(un4_v_low_s_2_9),.O(v_diff_1_axb_2));
defparam desc497.INIT=4'h9;
  LUT2 desc498(.I0(un4_v_high_s_3_9),.I1(un4_v_low_s_3_9),.O(v_diff_1_axb_3));
defparam desc498.INIT=4'h9;
  LUT2 desc499(.I0(un4_v_high_s_4_9),.I1(un4_v_low_s_4_9),.O(v_diff_1_axb_4));
defparam desc499.INIT=4'h9;
  LUT2 desc500(.I0(un4_v_high_s_5_9),.I1(un4_v_low_s_5_9),.O(v_diff_1_axb_5));
defparam desc500.INIT=4'h9;
  LUT2 desc501(.I0(un4_v_high_s_6_9),.I1(un4_v_low_s_6_9),.O(v_diff_1_axb_6));
defparam desc501.INIT=4'h9;
  LUT2 desc502(.I0(un4_v_high_s_7_9),.I1(un4_v_low_s_7_9),.O(v_diff_1_axb_7));
defparam desc502.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_6[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_6[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_6[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_6[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_6[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_6[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_6[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_7[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_7[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_7[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_7[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_7[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_7[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_7[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_7[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc503(.I0(acs_prob_tdata_6[0:0]),.I1(acs_prob_tdata_7[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2168));
defparam desc503.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_7[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_6[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc504(.I0(un4_v_high_s_8_9),.I1(un4_v_low_s_8_9),.O(v_diff_1_axb_8));
defparam desc504.INIT=4'h9;
  LUT6 desc505(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4_rep1),.I2(write_ram_fsm[0:0]),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc505.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIO0G81(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIO0G81.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIA3LB1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIA3LB1));
defparam s_axis_inbranch_tlast_d_RNIA3LB1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_6[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIITE71_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_9));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_9));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_7[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_9));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_7[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_9));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_7[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_9));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_7[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_9));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_7[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_9));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_7[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_9));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_7[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_7[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_9));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_9));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_6[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_9));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_6[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_9));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_6[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_9));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_6[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_9));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_6[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_9));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_6[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_9));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_6[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_6[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc506(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc507(.DI(un4_v_low_s_7_9),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc508(.DI(un4_v_low_s_6_9),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc509(.DI(un4_v_low_s_5_9),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc510(.DI(un4_v_low_s_4_9),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc511(.DI(un4_v_low_s_3_9),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc512(.DI(un4_v_low_s_2_9),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc513(.DI(un4_v_low_s_1_9),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc514(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc515(.Q(acs_prob_tdata_3[0:0]),.D(N_2168),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIA3LB1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc515_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc516(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIITE71_O6));
defparam desc516.INIT=16'hF4F0;
  LUT2 desc517(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc517.INIT=4'h8;
endmodule
module acsZ0_11_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_61,acs_prob_tdata_60,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_62,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,N_1756_1,aresetn,p_desc524_p_O_FD,p_desc525_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc554_p_O_FDRE);
input branch_tlast ;
output [62:62] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_61 ;
input [8:0] acs_prob_tdata_60 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_62 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIHCOU_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIKDM21 ;
wire un4_v_high_s_7_10 ;
wire un4_v_low_s_7_10 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_10 ;
wire un4_v_low_s_8_10 ;
wire un4_v_high_s_6_10 ;
wire un4_v_low_s_6_10 ;
wire un4_v_high_s_5_10 ;
wire un4_v_low_s_5_10 ;
wire un4_v_high_s_4_10 ;
wire un4_v_low_s_4_10 ;
wire un4_v_high_s_3_10 ;
wire un4_v_low_s_3_10 ;
wire un4_v_high_s_2_10 ;
wire un4_v_low_s_2_10 ;
wire un4_v_high_s_1_10 ;
wire un4_v_low_s_1_10 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2148 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc524_p_O_FD ;
input p_desc525_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc554_p_O_FDRE ;
// instances
  FDR desc518(.Q(acs_prob_tdata_62[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  FDR desc519(.Q(acs_prob_tdata_62[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  FDR desc520(.Q(acs_prob_tdata_62[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  FDR desc521(.Q(acs_prob_tdata_62[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  FDR desc522(.Q(acs_prob_tdata_62[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  FDR desc523(.Q(acs_prob_tdata_62[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21));
  p_O_FD desc524(.Q(acs_prob_tdata_62[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc524_p_O_FD));
  p_O_FD desc525(.Q(acs_prob_tdata_62[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc525_p_O_FD));
  LUT6 desc526(.I0(un4_v_high_s_7_10),.I1(un4_v_low_s_7_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKDM21),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc526.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc527(.I0(un4_v_high_s_8_10),.I1(un4_v_low_s_8_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKDM21),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc527.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc528(.I0(un4_v_high_s_6_10),.I1(un4_v_low_s_6_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc528.INIT=32'hACACFF00;
  LUT5 desc529(.I0(un4_v_high_s_5_10),.I1(un4_v_low_s_5_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc529.INIT=32'hACACFF00;
  LUT5 desc530(.I0(un4_v_high_s_4_10),.I1(un4_v_low_s_4_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc530.INIT=32'hACACFF00;
  LUT5 desc531(.I0(un4_v_high_s_3_10),.I1(un4_v_low_s_3_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc531.INIT=32'hACACFF00;
  LUT5 desc532(.I0(un4_v_high_s_2_10),.I1(un4_v_low_s_2_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc532.INIT=32'hACACFF00;
  LUT5 desc533(.I0(un4_v_high_s_1_10),.I1(un4_v_low_s_1_10),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_62[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc533.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[62:62]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc534(.I0(acs_prob_tdata_60[0:0]),.I1(acs_prob_tdata_61[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc534.INIT=16'h9669;
  LUT2 desc535(.I0(un4_v_high_s_1_10),.I1(un4_v_low_s_1_10),.O(v_diff_1_axb_1));
defparam desc535.INIT=4'h9;
  LUT2 desc536(.I0(un4_v_high_s_2_10),.I1(un4_v_low_s_2_10),.O(v_diff_1_axb_2));
defparam desc536.INIT=4'h9;
  LUT2 desc537(.I0(un4_v_high_s_3_10),.I1(un4_v_low_s_3_10),.O(v_diff_1_axb_3));
defparam desc537.INIT=4'h9;
  LUT2 desc538(.I0(un4_v_high_s_4_10),.I1(un4_v_low_s_4_10),.O(v_diff_1_axb_4));
defparam desc538.INIT=4'h9;
  LUT2 desc539(.I0(un4_v_high_s_5_10),.I1(un4_v_low_s_5_10),.O(v_diff_1_axb_5));
defparam desc539.INIT=4'h9;
  LUT2 desc540(.I0(un4_v_high_s_6_10),.I1(un4_v_low_s_6_10),.O(v_diff_1_axb_6));
defparam desc540.INIT=4'h9;
  LUT2 desc541(.I0(un4_v_high_s_7_10),.I1(un4_v_low_s_7_10),.O(v_diff_1_axb_7));
defparam desc541.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_60[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_60[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_60[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_60[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_60[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_60[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_60[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_61[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_61[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_61[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_61[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_61[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_61[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_61[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_61[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc542(.I0(acs_prob_tdata_60[0:0]),.I1(acs_prob_tdata_61[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2148));
defparam desc542.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_61[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_60[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc543(.I0(un4_v_high_s_8_10),.I1(un4_v_low_s_8_10),.O(v_diff_1_axb_8));
defparam desc543.INIT=4'h9;
  LUT6 desc544(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc544.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI2BHV(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI2BHV.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIKDM21_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIKDM21));
defparam s_axis_inbranch_tlast_d_RNIKDM21_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_60[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIHCOU_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_10));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_10));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_61[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_10));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_61[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_10));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_61[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_10));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_61[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_10));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_61[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_10));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_61[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_10));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_61[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_61[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_10));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_10));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_60[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_10));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_60[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_10));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_60[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_10));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_60[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_10));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_60[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_10));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_60[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_10));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_60[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_60[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc545(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc546(.DI(un4_v_low_s_7_10),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc547(.DI(un4_v_low_s_6_10),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc548(.DI(un4_v_low_s_5_10),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc549(.DI(un4_v_low_s_4_10),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc550(.DI(un4_v_low_s_3_10),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc551(.DI(un4_v_low_s_2_10),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc552(.DI(un4_v_low_s_1_10),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc553(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc554(.Q(acs_prob_tdata_62[0:0]),.D(N_2148),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKDM21),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc554_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc555(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIHCOU_O6));
defparam desc555.INIT=16'hF4F0;
  LUT2 desc556(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc556.INIT=4'h8;
endmodule
module acsZ0_12_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_31,acs_prob_tdata_30,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_47,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,N_1756_1,aresetn,p_desc563_p_O_FD,p_desc564_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc593_p_O_FDRE);
input branch_tlast ;
output [47:47] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_31 ;
input [8:0] acs_prob_tdata_30 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_47 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIQ8BO_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIQIP21 ;
wire un4_v_high_s_7_11 ;
wire un4_v_low_s_7_11 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_11 ;
wire un4_v_low_s_8_11 ;
wire un4_v_high_s_6_11 ;
wire un4_v_low_s_6_11 ;
wire un4_v_high_s_5_11 ;
wire un4_v_low_s_5_11 ;
wire un4_v_high_s_4_11 ;
wire un4_v_low_s_4_11 ;
wire un4_v_high_s_3_11 ;
wire un4_v_low_s_3_11 ;
wire un4_v_high_s_2_11 ;
wire un4_v_low_s_2_11 ;
wire un4_v_high_s_1_11 ;
wire un4_v_low_s_1_11 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2128 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc563_p_O_FD ;
input p_desc564_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc593_p_O_FDRE ;
// instances
  FDR desc557(.Q(acs_prob_tdata_47[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  FDR desc558(.Q(acs_prob_tdata_47[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  FDR desc559(.Q(acs_prob_tdata_47[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  FDR desc560(.Q(acs_prob_tdata_47[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  FDR desc561(.Q(acs_prob_tdata_47[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  FDR desc562(.Q(acs_prob_tdata_47[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21));
  p_O_FD desc563(.Q(acs_prob_tdata_47[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc563_p_O_FD));
  p_O_FD desc564(.Q(acs_prob_tdata_47[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc564_p_O_FD));
  LUT6 desc565(.I0(un4_v_high_s_7_11),.I1(un4_v_low_s_7_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQIP21),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc565.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc566(.I0(un4_v_high_s_8_11),.I1(un4_v_low_s_8_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQIP21),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc566.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc567(.I0(un4_v_high_s_6_11),.I1(un4_v_low_s_6_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc567.INIT=32'hACACFF00;
  LUT5 desc568(.I0(un4_v_high_s_5_11),.I1(un4_v_low_s_5_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc568.INIT=32'hACACFF00;
  LUT5 desc569(.I0(un4_v_high_s_4_11),.I1(un4_v_low_s_4_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc569.INIT=32'hACACFF00;
  LUT5 desc570(.I0(un4_v_high_s_3_11),.I1(un4_v_low_s_3_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc570.INIT=32'hACACFF00;
  LUT5 desc571(.I0(un4_v_high_s_2_11),.I1(un4_v_low_s_2_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc571.INIT=32'hACACFF00;
  LUT5 desc572(.I0(un4_v_high_s_1_11),.I1(un4_v_low_s_1_11),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_47[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc572.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[47:47]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc573(.I0(acs_prob_tdata_30[0:0]),.I1(acs_prob_tdata_31[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc573.INIT=16'h9669;
  LUT2 desc574(.I0(un4_v_high_s_1_11),.I1(un4_v_low_s_1_11),.O(v_diff_1_axb_1));
defparam desc574.INIT=4'h9;
  LUT2 desc575(.I0(un4_v_high_s_2_11),.I1(un4_v_low_s_2_11),.O(v_diff_1_axb_2));
defparam desc575.INIT=4'h9;
  LUT2 desc576(.I0(un4_v_high_s_3_11),.I1(un4_v_low_s_3_11),.O(v_diff_1_axb_3));
defparam desc576.INIT=4'h9;
  LUT2 desc577(.I0(un4_v_high_s_4_11),.I1(un4_v_low_s_4_11),.O(v_diff_1_axb_4));
defparam desc577.INIT=4'h9;
  LUT2 desc578(.I0(un4_v_high_s_5_11),.I1(un4_v_low_s_5_11),.O(v_diff_1_axb_5));
defparam desc578.INIT=4'h9;
  LUT2 desc579(.I0(un4_v_high_s_6_11),.I1(un4_v_low_s_6_11),.O(v_diff_1_axb_6));
defparam desc579.INIT=4'h9;
  LUT2 desc580(.I0(un4_v_high_s_7_11),.I1(un4_v_low_s_7_11),.O(v_diff_1_axb_7));
defparam desc580.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_30[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_30[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_30[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_30[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_30[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_30[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_30[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_31[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_31[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_31[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_31[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_31[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_31[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_31[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_31[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc581(.I0(acs_prob_tdata_30[0:0]),.I1(acs_prob_tdata_31[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2128));
defparam desc581.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_31[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_30[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc582(.I0(un4_v_high_s_8_11),.I1(un4_v_low_s_8_11),.O(v_diff_1_axb_8));
defparam desc582.INIT=4'h9;
  LUT6 desc583(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc583.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI8GKV(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI8GKV.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIQIP21_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIQIP21));
defparam s_axis_inbranch_tlast_d_RNIQIP21_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_30[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIQ8BO_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_11));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_11));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_31[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_11));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_31[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_11));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_31[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_11));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_31[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_11));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_31[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_11));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_31[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_11));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_31[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_31[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_11));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_11));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_30[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_11));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_30[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_11));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_30[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_11));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_30[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_11));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_30[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_11));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_30[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_11));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_30[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_30[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc584(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc585(.DI(un4_v_low_s_7_11),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc586(.DI(un4_v_low_s_6_11),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc587(.DI(un4_v_low_s_5_11),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc588(.DI(un4_v_low_s_4_11),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc589(.DI(un4_v_low_s_3_11),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc590(.DI(un4_v_low_s_2_11),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc591(.DI(un4_v_low_s_1_11),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc592(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc593(.Q(acs_prob_tdata_47[0:0]),.D(N_2128),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQIP21),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc593_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc594(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIQ8BO_O6));
defparam desc594.INIT=16'hF4F0;
  LUT2 desc595(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc595.INIT=4'h8;
endmodule
module acsZ0_13_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_11,acs_prob_tdata_10,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_5,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc602_p_O_FD,p_desc603_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc632_p_O_FDRE);
input branch_tlast ;
output [5:5] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_11 ;
input [8:0] acs_prob_tdata_10 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_5 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIO9ED1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIE9RF1 ;
wire un4_v_high_s_7_12 ;
wire un4_v_low_s_7_12 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_12 ;
wire un4_v_low_s_8_12 ;
wire un4_v_high_s_6_12 ;
wire un4_v_low_s_6_12 ;
wire un4_v_high_s_5_12 ;
wire un4_v_low_s_5_12 ;
wire un4_v_high_s_4_12 ;
wire un4_v_low_s_4_12 ;
wire un4_v_high_s_3_12 ;
wire un4_v_low_s_3_12 ;
wire un4_v_high_s_2_12 ;
wire un4_v_low_s_2_12 ;
wire un4_v_high_s_1_12 ;
wire un4_v_low_s_1_12 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_2108 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc602_p_O_FD ;
input p_desc603_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc632_p_O_FDRE ;
// instances
  FDR desc596(.Q(acs_prob_tdata_5[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  FDR desc597(.Q(acs_prob_tdata_5[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  FDR desc598(.Q(acs_prob_tdata_5[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  FDR desc599(.Q(acs_prob_tdata_5[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  FDR desc600(.Q(acs_prob_tdata_5[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  FDR desc601(.Q(acs_prob_tdata_5[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1));
  p_O_FD desc602(.Q(acs_prob_tdata_5[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc602_p_O_FD));
  p_O_FD desc603(.Q(acs_prob_tdata_5[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc603_p_O_FD));
  LUT6 desc604(.I0(un4_v_high_s_7_12),.I1(un4_v_low_s_7_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE9RF1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc604.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc605(.I0(un4_v_high_s_8_12),.I1(un4_v_low_s_8_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE9RF1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc605.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc606(.I0(un4_v_high_s_6_12),.I1(un4_v_low_s_6_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc606.INIT=32'hACACFF00;
  LUT5 desc607(.I0(un4_v_high_s_5_12),.I1(un4_v_low_s_5_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc607.INIT=32'hACACFF00;
  LUT5 desc608(.I0(un4_v_high_s_4_12),.I1(un4_v_low_s_4_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc608.INIT=32'hACACFF00;
  LUT5 desc609(.I0(un4_v_high_s_3_12),.I1(un4_v_low_s_3_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc609.INIT=32'hACACFF00;
  LUT5 desc610(.I0(un4_v_high_s_2_12),.I1(un4_v_low_s_2_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc610.INIT=32'hACACFF00;
  LUT5 desc611(.I0(un4_v_high_s_1_12),.I1(un4_v_low_s_1_12),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_5[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc611.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[5:5]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_10[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_10[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_10[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_10[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_10[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_10[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_10[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_11[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_11[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_11[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_11[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_11[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_11[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_11[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_11[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc612(.I0(acs_prob_tdata_10[0:0]),.I1(acs_prob_tdata_11[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc612.INIT=16'h9669;
  LUT2 desc613(.I0(un4_v_high_s_1_12),.I1(un4_v_low_s_1_12),.O(v_diff_1_axb_1));
defparam desc613.INIT=4'h9;
  LUT2 desc614(.I0(un4_v_high_s_2_12),.I1(un4_v_low_s_2_12),.O(v_diff_1_axb_2));
defparam desc614.INIT=4'h9;
  LUT2 desc615(.I0(un4_v_high_s_3_12),.I1(un4_v_low_s_3_12),.O(v_diff_1_axb_3));
defparam desc615.INIT=4'h9;
  LUT2 desc616(.I0(un4_v_high_s_4_12),.I1(un4_v_low_s_4_12),.O(v_diff_1_axb_4));
defparam desc616.INIT=4'h9;
  LUT2 desc617(.I0(un4_v_high_s_5_12),.I1(un4_v_low_s_5_12),.O(v_diff_1_axb_5));
defparam desc617.INIT=4'h9;
  LUT2 desc618(.I0(un4_v_high_s_6_12),.I1(un4_v_low_s_6_12),.O(v_diff_1_axb_6));
defparam desc618.INIT=4'h9;
  LUT2 desc619(.I0(un4_v_high_s_7_12),.I1(un4_v_low_s_7_12),.O(v_diff_1_axb_7));
defparam desc619.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc620(.I0(acs_prob_tdata_10[0:0]),.I1(acs_prob_tdata_11[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2108));
defparam desc620.INIT=32'h3C3C55AA;
  LUT2 desc621(.I0(un4_v_high_s_8_12),.I1(un4_v_low_s_8_12),.O(v_diff_1_axb_8));
defparam desc621.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_11[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_10[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc622(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc622.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIS6MC1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIS6MC1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIE9RF1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIE9RF1));
defparam s_axis_inbranch_tlast_d_RNIE9RF1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_10[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIO9ED1_O6),.C(aclk),.R(aresetn_i));
  XORCY desc623(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc624(.DI(un4_v_low_s_7_12),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc625(.DI(un4_v_low_s_6_12),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc626(.DI(un4_v_low_s_5_12),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc627(.DI(un4_v_low_s_4_12),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc628(.DI(un4_v_low_s_3_12),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc629(.DI(un4_v_low_s_2_12),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc630(.DI(un4_v_low_s_1_12),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc631(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_12));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_12));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_11[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_12));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_11[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_12));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_11[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_12));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_11[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_12));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_11[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_12));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_11[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_12));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_11[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_11[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_12));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_12));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_10[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_12));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_10[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_12));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_10[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_12));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_10[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_12));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_10[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_12));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_10[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_12));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_10[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_10[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc632(.Q(acs_prob_tdata_5[0:0]),.D(N_2108),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE9RF1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc632_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc633(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIO9ED1_O6));
defparam desc633.INIT=16'hF4F0;
  LUT2 desc634(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc634.INIT=4'h8;
endmodule
module acsZ0_14_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_11,acs_prob_tdata_10,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_37,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc641_p_O_FD,p_desc642_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc671_p_O_FDRE);
input branch_tlast ;
output [37:37] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_11 ;
input [8:0] acs_prob_tdata_10 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_37 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNINFL51_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIODJD1 ;
wire un4_v_high_s_7_13 ;
wire un4_v_low_s_7_13 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_13 ;
wire un4_v_low_s_8_13 ;
wire un4_v_high_s_6_13 ;
wire un4_v_low_s_6_13 ;
wire un4_v_high_s_5_13 ;
wire un4_v_low_s_5_13 ;
wire un4_v_high_s_4_13 ;
wire un4_v_low_s_4_13 ;
wire un4_v_high_s_3_13 ;
wire un4_v_low_s_3_13 ;
wire un4_v_high_s_2_13 ;
wire un4_v_low_s_2_13 ;
wire un4_v_high_s_1_13 ;
wire un4_v_low_s_1_13 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_2088 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc641_p_O_FD ;
input p_desc642_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc671_p_O_FDRE ;
// instances
  FDR desc635(.Q(acs_prob_tdata_37[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  FDR desc636(.Q(acs_prob_tdata_37[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  FDR desc637(.Q(acs_prob_tdata_37[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  FDR desc638(.Q(acs_prob_tdata_37[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  FDR desc639(.Q(acs_prob_tdata_37[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  FDR desc640(.Q(acs_prob_tdata_37[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1));
  p_O_FD desc641(.Q(acs_prob_tdata_37[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc641_p_O_FD));
  p_O_FD desc642(.Q(acs_prob_tdata_37[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc642_p_O_FD));
  LUT6 desc643(.I0(un4_v_high_s_7_13),.I1(un4_v_low_s_7_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIODJD1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc643.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc644(.I0(un4_v_high_s_8_13),.I1(un4_v_low_s_8_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIODJD1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc644.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc645(.I0(un4_v_high_s_6_13),.I1(un4_v_low_s_6_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc645.INIT=32'hACACFF00;
  LUT5 desc646(.I0(un4_v_high_s_5_13),.I1(un4_v_low_s_5_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc646.INIT=32'hACACFF00;
  LUT5 desc647(.I0(un4_v_high_s_4_13),.I1(un4_v_low_s_4_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc647.INIT=32'hACACFF00;
  LUT5 desc648(.I0(un4_v_high_s_3_13),.I1(un4_v_low_s_3_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc648.INIT=32'hACACFF00;
  LUT5 desc649(.I0(un4_v_high_s_2_13),.I1(un4_v_low_s_2_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc649.INIT=32'hACACFF00;
  LUT5 desc650(.I0(un4_v_high_s_1_13),.I1(un4_v_low_s_1_13),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_37[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc650.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[37:37]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_10[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_10[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_10[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_10[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_10[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_10[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_10[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_11[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_11[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_11[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_11[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_11[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_11[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_11[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_11[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc651(.I0(acs_prob_tdata_10[0:0]),.I1(acs_prob_tdata_11[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc651.INIT=16'h9669;
  LUT2 desc652(.I0(un4_v_high_s_1_13),.I1(un4_v_low_s_1_13),.O(v_diff_1_axb_1));
defparam desc652.INIT=4'h9;
  LUT2 desc653(.I0(un4_v_high_s_2_13),.I1(un4_v_low_s_2_13),.O(v_diff_1_axb_2));
defparam desc653.INIT=4'h9;
  LUT2 desc654(.I0(un4_v_high_s_3_13),.I1(un4_v_low_s_3_13),.O(v_diff_1_axb_3));
defparam desc654.INIT=4'h9;
  LUT2 desc655(.I0(un4_v_high_s_4_13),.I1(un4_v_low_s_4_13),.O(v_diff_1_axb_4));
defparam desc655.INIT=4'h9;
  LUT2 desc656(.I0(un4_v_high_s_5_13),.I1(un4_v_low_s_5_13),.O(v_diff_1_axb_5));
defparam desc656.INIT=4'h9;
  LUT2 desc657(.I0(un4_v_high_s_6_13),.I1(un4_v_low_s_6_13),.O(v_diff_1_axb_6));
defparam desc657.INIT=4'h9;
  LUT2 desc658(.I0(un4_v_high_s_7_13),.I1(un4_v_low_s_7_13),.O(v_diff_1_axb_7));
defparam desc658.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc659(.I0(acs_prob_tdata_10[0:0]),.I1(acs_prob_tdata_11[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_2088));
defparam desc659.INIT=32'h33CC5A5A;
  LUT2 desc660(.I0(un4_v_high_s_8_13),.I1(un4_v_low_s_8_13),.O(v_diff_1_axb_8));
defparam desc660.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_11[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_10[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc661(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc661.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI6BEA1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI6BEA1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIODJD1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIODJD1));
defparam s_axis_inbranch_tlast_d_RNIODJD1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_10[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNINFL51_O6),.C(aclk),.R(aresetn_i));
  XORCY desc662(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc663(.DI(un4_v_low_s_7_13),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc664(.DI(un4_v_low_s_6_13),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc665(.DI(un4_v_low_s_5_13),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc666(.DI(un4_v_low_s_4_13),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc667(.DI(un4_v_low_s_3_13),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc668(.DI(un4_v_low_s_2_13),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc669(.DI(un4_v_low_s_1_13),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc670(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_13));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_13));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_11[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_13));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_11[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_13));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_11[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_13));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_11[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_13));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_11[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_13));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_11[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_13));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_11[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_11[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_13));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_13));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_10[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_13));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_10[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_13));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_10[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_13));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_10[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_13));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_10[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_13));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_10[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_13));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_10[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_10[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc671(.Q(acs_prob_tdata_37[0:0]),.D(N_2088),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIODJD1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc671_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc672(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNINFL51_O6));
defparam desc672.INIT=16'hF4F0;
  LUT2 desc673(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc673.INIT=4'h8;
endmodule
module acsZ0_15_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_34,acs_prob_tdata_35,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_49,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_3_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,N_1756_1,aresetn,p_desc680_p_O_FD,p_desc681_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc710_p_O_FDRE);
input branch_tlast ;
output [49:49] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_34 ;
input [8:0] acs_prob_tdata_35 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_49 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_3_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_3_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI0LAU_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIUOV61 ;
wire un4_v_high_s_7_14 ;
wire un4_v_low_s_7_14 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_14 ;
wire un4_v_low_s_8_14 ;
wire un4_v_high_s_6_14 ;
wire un4_v_low_s_6_14 ;
wire un4_v_high_s_5_14 ;
wire un4_v_low_s_5_14 ;
wire un4_v_high_s_4_14 ;
wire un4_v_low_s_4_14 ;
wire un4_v_high_s_3_14 ;
wire un4_v_low_s_3_14 ;
wire un4_v_high_s_2_14 ;
wire un4_v_low_s_2_14 ;
wire un4_v_high_s_1_14 ;
wire un4_v_low_s_1_14 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire N_2068 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire GND ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire N_1 ;
input p_desc680_p_O_FD ;
input p_desc681_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc710_p_O_FDRE ;
// instances
  FDR desc674(.Q(acs_prob_tdata_49[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  FDR desc675(.Q(acs_prob_tdata_49[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  FDR desc676(.Q(acs_prob_tdata_49[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  FDR desc677(.Q(acs_prob_tdata_49[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  FDR desc678(.Q(acs_prob_tdata_49[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  FDR desc679(.Q(acs_prob_tdata_49[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61));
  p_O_FD desc680(.Q(acs_prob_tdata_49[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc680_p_O_FD));
  p_O_FD desc681(.Q(acs_prob_tdata_49[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc681_p_O_FD));
  LUT6 desc682(.I0(un4_v_high_s_7_14),.I1(un4_v_low_s_7_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIUOV61),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc682.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc683(.I0(un4_v_high_s_8_14),.I1(un4_v_low_s_8_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIUOV61),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc683.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc684(.I0(un4_v_high_s_6_14),.I1(un4_v_low_s_6_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc684.INIT=32'hACACFF00;
  LUT5 desc685(.I0(un4_v_high_s_5_14),.I1(un4_v_low_s_5_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc685.INIT=32'hACACFF00;
  LUT5 desc686(.I0(un4_v_high_s_4_14),.I1(un4_v_low_s_4_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc686.INIT=32'hACACFF00;
  LUT5 desc687(.I0(un4_v_high_s_3_14),.I1(un4_v_low_s_3_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc687.INIT=32'hACACFF00;
  LUT5 desc688(.I0(un4_v_high_s_2_14),.I1(un4_v_low_s_2_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc688.INIT=32'hACACFF00;
  LUT5 desc689(.I0(un4_v_high_s_1_14),.I1(un4_v_low_s_1_14),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_49[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc689.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[49:49]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_35[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_35[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_35[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_35[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_35[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_35[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_35[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_35[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc690(.I0(acs_prob_tdata_34[0:0]),.I1(acs_prob_tdata_35[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc690.INIT=16'h9669;
  LUT2 desc691(.I0(un4_v_high_s_1_14),.I1(un4_v_low_s_1_14),.O(v_diff_1_axb_1));
defparam desc691.INIT=4'h9;
  LUT2 desc692(.I0(un4_v_high_s_2_14),.I1(un4_v_low_s_2_14),.O(v_diff_1_axb_2));
defparam desc692.INIT=4'h9;
  LUT2 desc693(.I0(un4_v_high_s_3_14),.I1(un4_v_low_s_3_14),.O(v_diff_1_axb_3));
defparam desc693.INIT=4'h9;
  LUT2 desc694(.I0(un4_v_high_s_4_14),.I1(un4_v_low_s_4_14),.O(v_diff_1_axb_4));
defparam desc694.INIT=4'h9;
  LUT2 desc695(.I0(un4_v_high_s_5_14),.I1(un4_v_low_s_5_14),.O(v_diff_1_axb_5));
defparam desc695.INIT=4'h9;
  LUT2 desc696(.I0(un4_v_high_s_6_14),.I1(un4_v_low_s_6_14),.O(v_diff_1_axb_6));
defparam desc696.INIT=4'h9;
  LUT2 desc697(.I0(un4_v_high_s_7_14),.I1(un4_v_low_s_7_14),.O(v_diff_1_axb_7));
defparam desc697.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_34[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_34[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_34[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_34[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_34[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_34[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_34[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc698(.I0(acs_prob_tdata_34[0:0]),.I1(acs_prob_tdata_35[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2068));
defparam desc698.INIT=32'h33CC5A5A;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_34[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc699(.I0(un4_v_high_s_8_14),.I1(un4_v_low_s_8_14),.O(v_diff_1_axb_8));
defparam desc699.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_35[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT6 desc700(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc700.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNICMQ31(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNICMQ31.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIUOV61_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIUOV61));
defparam s_axis_inbranch_tlast_d_RNIUOV61_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_34[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI0LAU_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_14));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_14));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_34[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_14));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_34[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_14));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_34[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_14));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_34[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_14));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_34[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_14));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_34[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_14));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_34[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_34[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc701(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc702(.DI(un4_v_low_s_7_14),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc703(.DI(un4_v_low_s_6_14),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc704(.DI(un4_v_low_s_5_14),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc705(.DI(un4_v_low_s_4_14),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc706(.DI(un4_v_low_s_3_14),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc707(.DI(un4_v_low_s_2_14),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc708(.DI(un4_v_low_s_1_14),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc709(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_14));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_14));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_35[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_14));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_35[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_14));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_35[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_14));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_35[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_14));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_35[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_14));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_35[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_14));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_35[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_35[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  p_O_FDRE desc710(.Q(acs_prob_tdata_49[0:0]),.D(N_2068),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUOV61),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc710_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc711(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI0LAU_O6));
defparam desc711.INIT=16'hF4F0;
  LUT2 desc712(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc712.INIT=4'h8;
endmodule
module acsZ0_16_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_5,acs_prob_tdata_4,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_34,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc719_p_O_FD,p_desc720_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc749_p_O_FDRE);
input branch_tlast ;
output [34:34] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_5 ;
input [8:0] acs_prob_tdata_4 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_34 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIEDMS_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNII4A71 ;
wire un4_v_high_s_7_15 ;
wire un4_v_low_s_7_15 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_15 ;
wire un4_v_low_s_8_15 ;
wire un4_v_high_s_6_15 ;
wire un4_v_low_s_6_15 ;
wire un4_v_high_s_5_15 ;
wire un4_v_low_s_5_15 ;
wire un4_v_high_s_4_15 ;
wire un4_v_low_s_4_15 ;
wire un4_v_high_s_3_15 ;
wire un4_v_low_s_3_15 ;
wire un4_v_high_s_2_15 ;
wire un4_v_low_s_2_15 ;
wire un4_v_high_s_1_15 ;
wire un4_v_low_s_1_15 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2048 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc719_p_O_FD ;
input p_desc720_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc749_p_O_FDRE ;
// instances
  FDR desc713(.Q(acs_prob_tdata_34[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  FDR desc714(.Q(acs_prob_tdata_34[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  FDR desc715(.Q(acs_prob_tdata_34[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  FDR desc716(.Q(acs_prob_tdata_34[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  FDR desc717(.Q(acs_prob_tdata_34[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  FDR desc718(.Q(acs_prob_tdata_34[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71));
  p_O_FD desc719(.Q(acs_prob_tdata_34[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc719_p_O_FD));
  p_O_FD desc720(.Q(acs_prob_tdata_34[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc720_p_O_FD));
  LUT6 desc721(.I0(un4_v_high_s_7_15),.I1(un4_v_low_s_7_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII4A71),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc721.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc722(.I0(un4_v_high_s_8_15),.I1(un4_v_low_s_8_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII4A71),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc722.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc723(.I0(un4_v_high_s_6_15),.I1(un4_v_low_s_6_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc723.INIT=32'hACACFF00;
  LUT5 desc724(.I0(un4_v_high_s_5_15),.I1(un4_v_low_s_5_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc724.INIT=32'hACACFF00;
  LUT5 desc725(.I0(un4_v_high_s_4_15),.I1(un4_v_low_s_4_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc725.INIT=32'hACACFF00;
  LUT5 desc726(.I0(un4_v_high_s_3_15),.I1(un4_v_low_s_3_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc726.INIT=32'hACACFF00;
  LUT5 desc727(.I0(un4_v_high_s_2_15),.I1(un4_v_low_s_2_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc727.INIT=32'hACACFF00;
  LUT5 desc728(.I0(un4_v_high_s_1_15),.I1(un4_v_low_s_1_15),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_34[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc728.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[34:34]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc729(.I0(acs_prob_tdata_4[0:0]),.I1(acs_prob_tdata_5[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc729.INIT=16'h9669;
  LUT2 desc730(.I0(un4_v_high_s_1_15),.I1(un4_v_low_s_1_15),.O(v_diff_1_axb_1));
defparam desc730.INIT=4'h9;
  LUT2 desc731(.I0(un4_v_high_s_2_15),.I1(un4_v_low_s_2_15),.O(v_diff_1_axb_2));
defparam desc731.INIT=4'h9;
  LUT2 desc732(.I0(un4_v_high_s_3_15),.I1(un4_v_low_s_3_15),.O(v_diff_1_axb_3));
defparam desc732.INIT=4'h9;
  LUT2 desc733(.I0(un4_v_high_s_4_15),.I1(un4_v_low_s_4_15),.O(v_diff_1_axb_4));
defparam desc733.INIT=4'h9;
  LUT2 desc734(.I0(un4_v_high_s_5_15),.I1(un4_v_low_s_5_15),.O(v_diff_1_axb_5));
defparam desc734.INIT=4'h9;
  LUT2 desc735(.I0(un4_v_high_s_6_15),.I1(un4_v_low_s_6_15),.O(v_diff_1_axb_6));
defparam desc735.INIT=4'h9;
  LUT2 desc736(.I0(un4_v_high_s_7_15),.I1(un4_v_low_s_7_15),.O(v_diff_1_axb_7));
defparam desc736.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_4[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_4[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_4[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_4[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_4[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_4[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_4[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_5[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_5[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_5[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_5[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_5[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_5[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_5[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_5[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc737(.I0(acs_prob_tdata_4[0:0]),.I1(acs_prob_tdata_5[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2048));
defparam desc737.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_5[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_4[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc738(.I0(un4_v_high_s_8_15),.I1(un4_v_low_s_8_15),.O(v_diff_1_axb_8));
defparam desc738.INIT=4'h9;
  LUT6 desc739(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc739.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI02541(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI02541.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNII4A71_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNII4A71));
defparam s_axis_inbranch_tlast_d_RNII4A71_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_4[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIEDMS_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_15));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_15));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_5[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_15));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_5[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_15));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_5[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_15));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_5[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_15));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_5[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_15));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_5[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_15));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_5[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_5[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_15));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_15));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_4[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_15));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_4[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_15));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_4[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_15));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_4[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_15));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_4[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_15));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_4[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_15));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_4[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_4[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc740(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc741(.DI(un4_v_low_s_7_15),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc742(.DI(un4_v_low_s_6_15),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc743(.DI(un4_v_low_s_5_15),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc744(.DI(un4_v_low_s_4_15),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc745(.DI(un4_v_low_s_3_15),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc746(.DI(un4_v_low_s_2_15),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc747(.DI(un4_v_low_s_1_15),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc748(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc749(.Q(acs_prob_tdata_34[0:0]),.D(N_2048),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII4A71),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc749_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc750(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIEDMS_O6));
defparam desc750.INIT=16'hF4F0;
  LUT2 desc751(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc751.INIT=4'h8;
endmodule
module acsZ0_17_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_39,acs_prob_tdata_38,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_19,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc758_p_O_FD,p_desc759_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc788_p_O_FDRE);
input branch_tlast ;
output [19:19] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_39 ;
input [8:0] acs_prob_tdata_38 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_19 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIN9961_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIO9D71 ;
wire un4_v_high_s_7_16 ;
wire un4_v_low_s_7_16 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_16 ;
wire un4_v_low_s_8_16 ;
wire un4_v_high_s_6_16 ;
wire un4_v_low_s_6_16 ;
wire un4_v_high_s_5_16 ;
wire un4_v_low_s_5_16 ;
wire un4_v_high_s_4_16 ;
wire un4_v_low_s_4_16 ;
wire un4_v_high_s_3_16 ;
wire un4_v_low_s_3_16 ;
wire un4_v_high_s_2_16 ;
wire un4_v_low_s_2_16 ;
wire un4_v_high_s_1_16 ;
wire un4_v_low_s_1_16 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2028 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc758_p_O_FD ;
input p_desc759_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc788_p_O_FDRE ;
// instances
  FDR desc752(.Q(acs_prob_tdata_19[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  FDR desc753(.Q(acs_prob_tdata_19[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  FDR desc754(.Q(acs_prob_tdata_19[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  FDR desc755(.Q(acs_prob_tdata_19[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  FDR desc756(.Q(acs_prob_tdata_19[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  FDR desc757(.Q(acs_prob_tdata_19[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71));
  p_O_FD desc758(.Q(acs_prob_tdata_19[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc758_p_O_FD));
  p_O_FD desc759(.Q(acs_prob_tdata_19[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc759_p_O_FD));
  LUT6 desc760(.I0(un4_v_high_s_7_16),.I1(un4_v_low_s_7_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIO9D71),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc760.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc761(.I0(un4_v_high_s_8_16),.I1(un4_v_low_s_8_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIO9D71),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc761.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc762(.I0(un4_v_high_s_6_16),.I1(un4_v_low_s_6_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc762.INIT=32'hACACFF00;
  LUT5 desc763(.I0(un4_v_high_s_5_16),.I1(un4_v_low_s_5_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc763.INIT=32'hACACFF00;
  LUT5 desc764(.I0(un4_v_high_s_4_16),.I1(un4_v_low_s_4_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc764.INIT=32'hACACFF00;
  LUT5 desc765(.I0(un4_v_high_s_3_16),.I1(un4_v_low_s_3_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc765.INIT=32'hACACFF00;
  LUT5 desc766(.I0(un4_v_high_s_2_16),.I1(un4_v_low_s_2_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc766.INIT=32'hACACFF00;
  LUT5 desc767(.I0(un4_v_high_s_1_16),.I1(un4_v_low_s_1_16),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_19[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc767.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[19:19]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc768(.I0(acs_prob_tdata_38[0:0]),.I1(acs_prob_tdata_39[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc768.INIT=16'h9669;
  LUT2 desc769(.I0(un4_v_high_s_1_16),.I1(un4_v_low_s_1_16),.O(v_diff_1_axb_1));
defparam desc769.INIT=4'h9;
  LUT2 desc770(.I0(un4_v_high_s_2_16),.I1(un4_v_low_s_2_16),.O(v_diff_1_axb_2));
defparam desc770.INIT=4'h9;
  LUT2 desc771(.I0(un4_v_high_s_3_16),.I1(un4_v_low_s_3_16),.O(v_diff_1_axb_3));
defparam desc771.INIT=4'h9;
  LUT2 desc772(.I0(un4_v_high_s_4_16),.I1(un4_v_low_s_4_16),.O(v_diff_1_axb_4));
defparam desc772.INIT=4'h9;
  LUT2 desc773(.I0(un4_v_high_s_5_16),.I1(un4_v_low_s_5_16),.O(v_diff_1_axb_5));
defparam desc773.INIT=4'h9;
  LUT2 desc774(.I0(un4_v_high_s_6_16),.I1(un4_v_low_s_6_16),.O(v_diff_1_axb_6));
defparam desc774.INIT=4'h9;
  LUT2 desc775(.I0(un4_v_high_s_7_16),.I1(un4_v_low_s_7_16),.O(v_diff_1_axb_7));
defparam desc775.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_38[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_38[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_38[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_38[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_38[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_38[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_38[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_39[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_39[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_39[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_39[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_39[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_39[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_39[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_39[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc776(.I0(acs_prob_tdata_38[0:0]),.I1(acs_prob_tdata_39[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2028));
defparam desc776.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_39[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_38[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc777(.I0(un4_v_high_s_8_16),.I1(un4_v_low_s_8_16),.O(v_diff_1_axb_8));
defparam desc777.INIT=4'h9;
  LUT6 desc778(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc778.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI67841(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI67841.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIO9D71_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIO9D71));
defparam s_axis_inbranch_tlast_d_RNIO9D71_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_38[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIN9961_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_16));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_16));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_39[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_16));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_39[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_16));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_39[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_16));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_39[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_16));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_39[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_16));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_39[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_16));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_39[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_39[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_16));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_16));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_38[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_16));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_38[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_16));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_38[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_16));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_38[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_16));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_38[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_16));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_38[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_16));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_38[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_38[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc779(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc780(.DI(un4_v_low_s_7_16),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc781(.DI(un4_v_low_s_6_16),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc782(.DI(un4_v_low_s_5_16),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc783(.DI(un4_v_low_s_4_16),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc784(.DI(un4_v_low_s_3_16),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc785(.DI(un4_v_low_s_2_16),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc786(.DI(un4_v_low_s_1_16),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc787(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc788(.Q(acs_prob_tdata_19[0:0]),.D(N_2028),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIO9D71),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc788_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc789(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIN9961_O6));
defparam desc789.INIT=16'hF4F0;
  LUT2 desc790(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc790.INIT=4'h8;
endmodule
module acsZ0_18_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_9,acs_prob_tdata_8,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_4,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_4_rep1,N_1756_1,aresetn,p_desc797_p_O_FD,p_desc798_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc827_p_O_FDRE);
input branch_tlast ;
output [4:4] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_9 ;
input [8:0] acs_prob_tdata_8 ;
input [1:0] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_4 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNILJEA1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIC6OD1 ;
wire un4_v_high_s_7_17 ;
wire un4_v_low_s_7_17 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_17 ;
wire un4_v_low_s_8_17 ;
wire un4_v_high_s_6_17 ;
wire un4_v_low_s_6_17 ;
wire un4_v_high_s_5_17 ;
wire un4_v_low_s_5_17 ;
wire un4_v_high_s_4_17 ;
wire un4_v_low_s_4_17 ;
wire un4_v_high_s_3_17 ;
wire un4_v_low_s_3_17 ;
wire un4_v_high_s_2_17 ;
wire un4_v_low_s_2_17 ;
wire un4_v_high_s_1_17 ;
wire un4_v_low_s_1_17 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_2008 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc797_p_O_FD ;
input p_desc798_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc827_p_O_FDRE ;
// instances
  FDR desc791(.Q(acs_prob_tdata_4[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  FDR desc792(.Q(acs_prob_tdata_4[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  FDR desc793(.Q(acs_prob_tdata_4[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  FDR desc794(.Q(acs_prob_tdata_4[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  FDR desc795(.Q(acs_prob_tdata_4[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  FDR desc796(.Q(acs_prob_tdata_4[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1));
  p_O_FD desc797(.Q(acs_prob_tdata_4[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc797_p_O_FD));
  p_O_FD desc798(.Q(acs_prob_tdata_4[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc798_p_O_FD));
  LUT6 desc799(.I0(un4_v_high_s_7_17),.I1(un4_v_low_s_7_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIC6OD1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc799.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc800(.I0(un4_v_high_s_8_17),.I1(un4_v_low_s_8_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIC6OD1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc800.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc801(.I0(un4_v_high_s_6_17),.I1(un4_v_low_s_6_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc801.INIT=32'hACACFF00;
  LUT5 desc802(.I0(un4_v_high_s_5_17),.I1(un4_v_low_s_5_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc802.INIT=32'hACACFF00;
  LUT5 desc803(.I0(un4_v_high_s_4_17),.I1(un4_v_low_s_4_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc803.INIT=32'hACACFF00;
  LUT5 desc804(.I0(un4_v_high_s_3_17),.I1(un4_v_low_s_3_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc804.INIT=32'hACACFF00;
  LUT5 desc805(.I0(un4_v_high_s_2_17),.I1(un4_v_low_s_2_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc805.INIT=32'hACACFF00;
  LUT5 desc806(.I0(un4_v_high_s_1_17),.I1(un4_v_low_s_1_17),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_4[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc806.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[4:4]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc807(.I0(acs_prob_tdata_8[0:0]),.I1(acs_prob_tdata_9[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc807.INIT=16'h9669;
  LUT2 desc808(.I0(un4_v_high_s_1_17),.I1(un4_v_low_s_1_17),.O(v_diff_1_axb_1));
defparam desc808.INIT=4'h9;
  LUT2 desc809(.I0(un4_v_high_s_2_17),.I1(un4_v_low_s_2_17),.O(v_diff_1_axb_2));
defparam desc809.INIT=4'h9;
  LUT2 desc810(.I0(un4_v_high_s_3_17),.I1(un4_v_low_s_3_17),.O(v_diff_1_axb_3));
defparam desc810.INIT=4'h9;
  LUT2 desc811(.I0(un4_v_high_s_4_17),.I1(un4_v_low_s_4_17),.O(v_diff_1_axb_4));
defparam desc811.INIT=4'h9;
  LUT2 desc812(.I0(un4_v_high_s_5_17),.I1(un4_v_low_s_5_17),.O(v_diff_1_axb_5));
defparam desc812.INIT=4'h9;
  LUT2 desc813(.I0(un4_v_high_s_6_17),.I1(un4_v_low_s_6_17),.O(v_diff_1_axb_6));
defparam desc813.INIT=4'h9;
  LUT2 desc814(.I0(un4_v_high_s_7_17),.I1(un4_v_low_s_7_17),.O(v_diff_1_axb_7));
defparam desc814.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_8[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_8[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_8[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_8[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_8[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_8[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_8[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_9[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_9[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_9[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_9[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_9[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_9[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_9[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_9[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc815(.I0(acs_prob_tdata_8[0:0]),.I1(acs_prob_tdata_9[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_2008));
defparam desc815.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_9[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_8[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc816(.I0(un4_v_high_s_8_17),.I1(un4_v_low_s_8_17),.O(v_diff_1_axb_8));
defparam desc816.INIT=4'h9;
  LUT6 desc817(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4_rep1),.I2(write_ram_fsm[0:0]),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc817.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIQ3JA1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQ3JA1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIC6OD1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIC6OD1));
defparam s_axis_inbranch_tlast_d_RNIC6OD1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_8[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNILJEA1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_17));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_17));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_9[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_17));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_9[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_17));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_9[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_17));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_9[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_17));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_9[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_17));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_9[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_17));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_9[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_9[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_17));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_17));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_8[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_17));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_8[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_17));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_8[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_17));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_8[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_17));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_8[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_17));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_8[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_17));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_8[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_8[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc818(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc819(.DI(un4_v_low_s_7_17),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc820(.DI(un4_v_low_s_6_17),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc821(.DI(un4_v_low_s_5_17),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc822(.DI(un4_v_low_s_4_17),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc823(.DI(un4_v_low_s_3_17),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc824(.DI(un4_v_low_s_2_17),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc825(.DI(un4_v_low_s_1_17),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc826(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc827(.Q(acs_prob_tdata_4[0:0]),.D(N_2008),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIC6OD1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc827_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc828(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNILJEA1_O6));
defparam desc828.INIT=16'hF4F0;
  LUT2 desc829(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc829.INIT=4'h8;
endmodule
module acsZ0_19_inj (branch_tvalid,acs_prob_tdata_63,acs_dec_tdata,branch_tdata_0_0,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_3,acs_prob_tdata_62,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tlast,branch_tdata_0_fast,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,N_1756_1,aresetn,p_m_axis_outdec_tdata_Z_p_O_FDRE);
input branch_tvalid ;
output [8:0] acs_prob_tdata_63 ;
output [63:63] acs_dec_tdata ;
input branch_tdata_0_0 ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_62 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tlast ;
input branch_tdata_0_fast ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_0 ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [8:0] m_axis_outprob_tdata_8_0 ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire s_axis_inbranch_tlast_d_RNIQ65C1_O5 ;
wire s_axis_inbranch_tlast_d_RNIMGP41 ;
wire un4_v_high_s_8_18 ;
wire un4_v_low_s_8_18 ;
wire un4_v_high_s_7_18 ;
wire un4_v_low_s_7_18 ;
wire un4_v_high_s_6_18 ;
wire un4_v_low_s_6_18 ;
wire un4_v_high_s_5_18 ;
wire un4_v_low_s_5_18 ;
wire un4_v_high_s_4_18 ;
wire un4_v_low_s_4_18 ;
wire un4_v_high_s_3_18 ;
wire un4_v_low_s_3_18 ;
wire un4_v_high_s_2_18 ;
wire un4_v_low_s_2_18 ;
wire un4_v_high_s_1_18 ;
wire un4_v_low_s_1_18 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire s_axis_inbranch_tlast_d_0 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
// instances
  FDR desc830(.Q(acs_prob_tdata_63[0:0]),.D(m_axis_outprob_tdata_8_0[0:0]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc831(.Q(acs_prob_tdata_63[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc832(.Q(acs_prob_tdata_63[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc833(.Q(acs_prob_tdata_63[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc834(.Q(acs_prob_tdata_63[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc835(.Q(acs_prob_tdata_63[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDR desc836(.Q(acs_prob_tdata_63[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMGP41));
  FDS desc837(.Q(acs_prob_tdata_63[7:7]),.D(m_axis_outprob_tdata_8_0[7:7]),.C(aclk),.S(s_axis_inbranch_tlast_d_RNIMGP41));
  FDS desc838(.Q(acs_prob_tdata_63[8:8]),.D(m_axis_outprob_tdata_8_0[8:8]),.C(aclk),.S(s_axis_inbranch_tlast_d_RNIMGP41));
  LUT5 desc839(.I0(un4_v_high_s_8_18),.I1(un4_v_low_s_8_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[8:8]));
defparam desc839.INIT=32'hACACFF00;
  LUT5 desc840(.I0(un4_v_high_s_7_18),.I1(un4_v_low_s_7_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[7:7]));
defparam desc840.INIT=32'hACACFF00;
  LUT5 desc841(.I0(un4_v_high_s_6_18),.I1(un4_v_low_s_6_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc841.INIT=32'hACACFF00;
  LUT5 desc842(.I0(un4_v_high_s_5_18),.I1(un4_v_low_s_5_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc842.INIT=32'hACACFF00;
  LUT5 desc843(.I0(un4_v_high_s_4_18),.I1(un4_v_low_s_4_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc843.INIT=32'hACACFF00;
  LUT5 desc844(.I0(un4_v_high_s_3_18),.I1(un4_v_low_s_3_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc844.INIT=32'hACACFF00;
  LUT5 desc845(.I0(un4_v_high_s_2_18),.I1(un4_v_low_s_2_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc845.INIT=32'hACACFF00;
  LUT5 desc846(.I0(un4_v_high_s_1_18),.I1(un4_v_low_s_1_18),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_63[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc846.INIT=32'hACACFF00;
  LUT6 desc847(.I0(acs_prob_tdata_62[0:0]),.I1(acs_prob_tdata_63[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.I5(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[0:0]));
defparam desc847.INIT=64'h33CC5A5ACCCCCCCC;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[63:63]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc848(.I0(acs_prob_tdata_62[0:0]),.I1(acs_prob_tdata_63[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc848.INIT=16'h9669;
  LUT2 desc849(.I0(un4_v_high_s_1_18),.I1(un4_v_low_s_1_18),.O(v_diff_1_axb_1));
defparam desc849.INIT=4'h9;
  LUT2 desc850(.I0(un4_v_high_s_2_18),.I1(un4_v_low_s_2_18),.O(v_diff_1_axb_2));
defparam desc850.INIT=4'h9;
  LUT2 desc851(.I0(un4_v_high_s_3_18),.I1(un4_v_low_s_3_18),.O(v_diff_1_axb_3));
defparam desc851.INIT=4'h9;
  LUT2 desc852(.I0(un4_v_high_s_4_18),.I1(un4_v_low_s_4_18),.O(v_diff_1_axb_4));
defparam desc852.INIT=4'h9;
  LUT2 desc853(.I0(un4_v_high_s_5_18),.I1(un4_v_low_s_5_18),.O(v_diff_1_axb_5));
defparam desc853.INIT=4'h9;
  LUT2 desc854(.I0(un4_v_high_s_6_18),.I1(un4_v_low_s_6_18),.O(v_diff_1_axb_6));
defparam desc854.INIT=4'h9;
  LUT2 desc855(.I0(un4_v_high_s_7_18),.I1(un4_v_low_s_7_18),.O(v_diff_1_axb_7));
defparam desc855.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_62[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_62[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_62[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_62[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_62[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_62[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_62[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_63[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_63[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_63[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_63[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_63[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_63[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_63[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_63[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_63[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_62[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc856(.I0(un4_v_high_s_8_18),.I1(un4_v_low_s_8_18),.O(v_diff_1_axb_8));
defparam desc856.INIT=4'h9;
  LUT6 desc857(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc857.INIT=64'h5557000055550000;
  LUT2_L s_axis_inbranch_tlast_d_e(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.LO(s_axis_inbranch_tlast_d_0));
defparam s_axis_inbranch_tlast_d_e.INIT=4'h8;
  LUT5 s_axis_inbranch_tlast_d_RNIMGP41_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIMGP41));
defparam s_axis_inbranch_tlast_d_RNIMGP41_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_62[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(s_axis_inbranch_tlast_d_RNIQ65C1_O5),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_18));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_18));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_63[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_18));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_63[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_18));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_63[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_18));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_63[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_18));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_63[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_18));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_63[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_18));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_63[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_63[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_18));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_18));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_62[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_18));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_62[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_18));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_62[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_18));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_62[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_18));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_62[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_18));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_62[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_18));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_62[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_62[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc858(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc859(.DI(un4_v_low_s_7_18),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc860(.DI(un4_v_low_s_6_18),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc861(.DI(un4_v_low_s_5_18),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc862(.DI(un4_v_low_s_4_18),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc863(.DI(un4_v_low_s_3_18),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc864(.DI(un4_v_low_s_2_18),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc865(.DI(un4_v_low_s_1_18),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc866(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 s_axis_inbranch_tlast_d_RNIQ65C1_o6(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQ65C1_o6.INIT=16'hBAFA;
  LUT4 s_axis_inbranch_tlast_d_RNIQ65C1_o5(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIQ65C1_O5));
defparam s_axis_inbranch_tlast_d_RNIQ65C1_o5.INIT=16'hF4F0;
endmodule
module acsZ0_20_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_59,acs_prob_tdata_58,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_61,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,N_1756_1,aresetn,p_desc873_p_O_FD,p_desc874_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc903_p_O_FDRE);
input branch_tlast ;
output [61:61] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_59 ;
input [8:0] acs_prob_tdata_58 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_61 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIEMOR_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIIAJ01 ;
wire un4_v_high_s_7_19 ;
wire un4_v_low_s_7_19 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_19 ;
wire un4_v_low_s_8_19 ;
wire un4_v_high_s_6_19 ;
wire un4_v_low_s_6_19 ;
wire un4_v_high_s_5_19 ;
wire un4_v_low_s_5_19 ;
wire un4_v_high_s_4_19 ;
wire un4_v_low_s_4_19 ;
wire un4_v_high_s_3_19 ;
wire un4_v_low_s_3_19 ;
wire un4_v_high_s_2_19 ;
wire un4_v_low_s_2_19 ;
wire un4_v_high_s_1_19 ;
wire un4_v_low_s_1_19 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1968 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc873_p_O_FD ;
input p_desc874_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc903_p_O_FDRE ;
// instances
  FDR desc867(.Q(acs_prob_tdata_61[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  FDR desc868(.Q(acs_prob_tdata_61[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  FDR desc869(.Q(acs_prob_tdata_61[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  FDR desc870(.Q(acs_prob_tdata_61[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  FDR desc871(.Q(acs_prob_tdata_61[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  FDR desc872(.Q(acs_prob_tdata_61[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01));
  p_O_FD desc873(.Q(acs_prob_tdata_61[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc873_p_O_FD));
  p_O_FD desc874(.Q(acs_prob_tdata_61[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc874_p_O_FD));
  LUT6 desc875(.I0(un4_v_high_s_7_19),.I1(un4_v_low_s_7_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIIAJ01),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc875.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc876(.I0(un4_v_high_s_8_19),.I1(un4_v_low_s_8_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIIAJ01),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc876.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc877(.I0(un4_v_high_s_6_19),.I1(un4_v_low_s_6_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc877.INIT=32'hACACFF00;
  LUT5 desc878(.I0(un4_v_high_s_5_19),.I1(un4_v_low_s_5_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc878.INIT=32'hACACFF00;
  LUT5 desc879(.I0(un4_v_high_s_4_19),.I1(un4_v_low_s_4_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc879.INIT=32'hACACFF00;
  LUT5 desc880(.I0(un4_v_high_s_3_19),.I1(un4_v_low_s_3_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc880.INIT=32'hACACFF00;
  LUT5 desc881(.I0(un4_v_high_s_2_19),.I1(un4_v_low_s_2_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc881.INIT=32'hACACFF00;
  LUT5 desc882(.I0(un4_v_high_s_1_19),.I1(un4_v_low_s_1_19),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_61[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc882.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[61:61]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc883(.I0(acs_prob_tdata_58[0:0]),.I1(acs_prob_tdata_59[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc883.INIT=16'h9669;
  LUT2 desc884(.I0(un4_v_high_s_1_19),.I1(un4_v_low_s_1_19),.O(v_diff_1_axb_1));
defparam desc884.INIT=4'h9;
  LUT2 desc885(.I0(un4_v_high_s_2_19),.I1(un4_v_low_s_2_19),.O(v_diff_1_axb_2));
defparam desc885.INIT=4'h9;
  LUT2 desc886(.I0(un4_v_high_s_3_19),.I1(un4_v_low_s_3_19),.O(v_diff_1_axb_3));
defparam desc886.INIT=4'h9;
  LUT2 desc887(.I0(un4_v_high_s_4_19),.I1(un4_v_low_s_4_19),.O(v_diff_1_axb_4));
defparam desc887.INIT=4'h9;
  LUT2 desc888(.I0(un4_v_high_s_5_19),.I1(un4_v_low_s_5_19),.O(v_diff_1_axb_5));
defparam desc888.INIT=4'h9;
  LUT2 desc889(.I0(un4_v_high_s_6_19),.I1(un4_v_low_s_6_19),.O(v_diff_1_axb_6));
defparam desc889.INIT=4'h9;
  LUT2 desc890(.I0(un4_v_high_s_7_19),.I1(un4_v_low_s_7_19),.O(v_diff_1_axb_7));
defparam desc890.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_58[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_58[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_58[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_58[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_58[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_58[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_58[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_59[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_59[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_59[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_59[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_59[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_59[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_59[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_59[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc891(.I0(acs_prob_tdata_58[0:0]),.I1(acs_prob_tdata_59[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1968));
defparam desc891.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_59[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_58[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc892(.I0(un4_v_high_s_8_19),.I1(un4_v_low_s_8_19),.O(v_diff_1_axb_8));
defparam desc892.INIT=4'h9;
  LUT6 desc893(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc893.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI08ET(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI08ET.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIIAJ01_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIIAJ01));
defparam s_axis_inbranch_tlast_d_RNIIAJ01_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_58[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIEMOR_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_19));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_19));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_59[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_19));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_59[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_19));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_59[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_19));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_59[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_19));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_59[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_19));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_59[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_19));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_59[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_59[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_19));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_19));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_58[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_19));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_58[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_19));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_58[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_19));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_58[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_19));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_58[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_19));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_58[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_19));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_58[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_58[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc894(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc895(.DI(un4_v_low_s_7_19),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc896(.DI(un4_v_low_s_6_19),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc897(.DI(un4_v_low_s_5_19),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc898(.DI(un4_v_low_s_4_19),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc899(.DI(un4_v_low_s_3_19),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc900(.DI(un4_v_low_s_2_19),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc901(.DI(un4_v_low_s_1_19),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc902(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc903(.Q(acs_prob_tdata_61[0:0]),.D(N_1968),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIAJ01),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc903_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc904(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIEMOR_O6));
defparam desc904.INIT=16'hF4F0;
  LUT2 desc905(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc905.INIT=4'h8;
endmodule
module acsZ0_21_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_1,acs_prob_tdata_0,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_32,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc912_p_O_FD,p_desc913_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc942_p_O_FDRE);
input branch_tlast ;
output [32:32] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_1 ;
input [8:0] acs_prob_tdata_0 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_32 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI81NM_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIEU331 ;
wire un4_v_high_s_7_20 ;
wire un4_v_low_s_7_20 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_20 ;
wire un4_v_low_s_8_20 ;
wire un4_v_high_s_6_20 ;
wire un4_v_low_s_6_20 ;
wire un4_v_high_s_5_20 ;
wire un4_v_low_s_5_20 ;
wire un4_v_high_s_4_20 ;
wire un4_v_low_s_4_20 ;
wire un4_v_high_s_3_20 ;
wire un4_v_low_s_3_20 ;
wire un4_v_high_s_2_20 ;
wire un4_v_low_s_2_20 ;
wire un4_v_high_s_1_20 ;
wire un4_v_low_s_1_20 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1948 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc912_p_O_FD ;
input p_desc913_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc942_p_O_FDRE ;
// instances
  FDR desc906(.Q(acs_prob_tdata_32[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  FDR desc907(.Q(acs_prob_tdata_32[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  FDR desc908(.Q(acs_prob_tdata_32[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  FDR desc909(.Q(acs_prob_tdata_32[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  FDR desc910(.Q(acs_prob_tdata_32[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  FDR desc911(.Q(acs_prob_tdata_32[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331));
  p_O_FD desc912(.Q(acs_prob_tdata_32[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc912_p_O_FD));
  p_O_FD desc913(.Q(acs_prob_tdata_32[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc913_p_O_FD));
  LUT6 desc914(.I0(un4_v_high_s_7_20),.I1(un4_v_low_s_7_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIEU331),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc914.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc915(.I0(un4_v_high_s_8_20),.I1(un4_v_low_s_8_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIEU331),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc915.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc916(.I0(un4_v_high_s_6_20),.I1(un4_v_low_s_6_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc916.INIT=32'hACACFF00;
  LUT5 desc917(.I0(un4_v_high_s_5_20),.I1(un4_v_low_s_5_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc917.INIT=32'hACACFF00;
  LUT5 desc918(.I0(un4_v_high_s_4_20),.I1(un4_v_low_s_4_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc918.INIT=32'hACACFF00;
  LUT5 desc919(.I0(un4_v_high_s_3_20),.I1(un4_v_low_s_3_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc919.INIT=32'hACACFF00;
  LUT5 desc920(.I0(un4_v_high_s_2_20),.I1(un4_v_low_s_2_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc920.INIT=32'hACACFF00;
  LUT5 desc921(.I0(un4_v_high_s_1_20),.I1(un4_v_low_s_1_20),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_32[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc921.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[32:32]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_0[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_0[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_0[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_0[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_0[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_0[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_0[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_1[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_1[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_1[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_1[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_1[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_1[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_1[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_1[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc922(.I0(acs_prob_tdata_0[0:0]),.I1(acs_prob_tdata_1[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc922.INIT=16'h9669;
  LUT2 desc923(.I0(un4_v_high_s_1_20),.I1(un4_v_low_s_1_20),.O(v_diff_1_axb_1));
defparam desc923.INIT=4'h9;
  LUT2 desc924(.I0(un4_v_high_s_2_20),.I1(un4_v_low_s_2_20),.O(v_diff_1_axb_2));
defparam desc924.INIT=4'h9;
  LUT2 desc925(.I0(un4_v_high_s_3_20),.I1(un4_v_low_s_3_20),.O(v_diff_1_axb_3));
defparam desc925.INIT=4'h9;
  LUT2 desc926(.I0(un4_v_high_s_4_20),.I1(un4_v_low_s_4_20),.O(v_diff_1_axb_4));
defparam desc926.INIT=4'h9;
  LUT2 desc927(.I0(un4_v_high_s_5_20),.I1(un4_v_low_s_5_20),.O(v_diff_1_axb_5));
defparam desc927.INIT=4'h9;
  LUT2 desc928(.I0(un4_v_high_s_6_20),.I1(un4_v_low_s_6_20),.O(v_diff_1_axb_6));
defparam desc928.INIT=4'h9;
  LUT2 desc929(.I0(un4_v_high_s_7_20),.I1(un4_v_low_s_7_20),.O(v_diff_1_axb_7));
defparam desc929.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc930(.I0(acs_prob_tdata_0[0:0]),.I1(acs_prob_tdata_1[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1948));
defparam desc930.INIT=32'h3C3C55AA;
  LUT2 desc931(.I0(un4_v_high_s_8_20),.I1(un4_v_low_s_8_20),.O(v_diff_1_axb_8));
defparam desc931.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_1[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_0[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc932(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc932.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNISRUV(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNISRUV.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIEU331_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIEU331));
defparam s_axis_inbranch_tlast_d_RNIEU331_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_0[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI81NM_O6),.C(aclk),.R(aresetn_i));
  XORCY desc933(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc934(.DI(un4_v_low_s_7_20),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc935(.DI(un4_v_low_s_6_20),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc936(.DI(un4_v_low_s_5_20),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc937(.DI(un4_v_low_s_4_20),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc938(.DI(un4_v_low_s_3_20),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc939(.DI(un4_v_low_s_2_20),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc940(.DI(un4_v_low_s_1_20),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc941(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_20));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_20));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_1[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_20));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_1[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_20));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_1[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_20));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_1[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_20));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_1[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_20));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_1[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_20));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_1[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_1[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_20));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_20));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_0[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_20));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_0[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_20));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_0[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_20));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_0[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_20));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_0[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_20));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_0[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_20));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_0[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_0[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc942(.Q(acs_prob_tdata_32[0:0]),.D(N_1948),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEU331),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc942_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc943(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI81NM_O6));
defparam desc943.INIT=16'hF4F0;
  LUT2 desc944(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc944.INIT=4'h8;
endmodule
module acsZ1_inj (acs_tvalid,branch_tlast,branch_tvalid,acs_prob_tdata_0,acs_dec_tdata,branch_tdata_0_0,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_3,acs_prob_tdata_1,write_ram_fsm,branch_tdata_0_fast,acs_tlast,un27_s_axis_input_tready_int,un1_output_accept,s_axis_inbranch_tlast_d_RNIIAVE1_O5,aclk,aresetn_i,branch_tdata_3_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep1,N_1756_1,un1_s_axis_input_tvalid,aresetn);
output acs_tvalid ;
input branch_tlast ;
input branch_tvalid ;
output [8:0] acs_prob_tdata_0 ;
output acs_dec_tdata ;
input branch_tdata_0_0 ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_1 ;
input [1:1] write_ram_fsm ;
input branch_tdata_0_fast ;
output acs_tlast ;
input un27_s_axis_input_tready_int ;
input un1_output_accept ;
output s_axis_inbranch_tlast_d_RNIIAVE1_O5 ;
input aclk ;
input aresetn_i ;
input branch_tdata_3_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
output un1_s_axis_input_tvalid ;
input aresetn ;
wire branch_tdata_0_0 ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire un27_s_axis_input_tready_int ;
wire un1_output_accept ;
wire s_axis_inbranch_tlast_d_RNIIAVE1_O5 ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_3_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire un1_s_axis_input_tvalid ;
wire aresetn ;
wire [8:0] m_axis_outprob_tdata_17_0 ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire VCC ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_e_lut6_2_O5 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire s_axis_inbranch_tlast_d_RNI4QB51 ;
wire m_axis_outprob_tdata_0_sqmuxa_set ;
wire un4_v_high_s_8_21 ;
wire un4_v_low_s_8_21 ;
wire un4_v_high_s_7_21 ;
wire un4_v_low_s_7_21 ;
wire un4_v_high_s_6_21 ;
wire un4_v_low_s_6_21 ;
wire un4_v_high_s_5_21 ;
wire un4_v_low_s_5_21 ;
wire un4_v_high_s_4_21 ;
wire un4_v_low_s_4_21 ;
wire un4_v_high_s_3_21 ;
wire un4_v_low_s_3_21 ;
wire un4_v_high_s_2_21 ;
wire un4_v_low_s_2_21 ;
wire un4_v_high_s_1_21 ;
wire un4_v_low_s_1_21 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
// instances
  FDR desc945(.Q(acs_prob_tdata_0[0:0]),.D(m_axis_outprob_tdata_17_0[0:0]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc946(.Q(acs_prob_tdata_0[1:1]),.D(m_axis_outprob_tdata_17_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc947(.Q(acs_prob_tdata_0[2:2]),.D(m_axis_outprob_tdata_17_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc948(.Q(acs_prob_tdata_0[3:3]),.D(m_axis_outprob_tdata_17_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc949(.Q(acs_prob_tdata_0[4:4]),.D(m_axis_outprob_tdata_17_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc950(.Q(acs_prob_tdata_0[5:5]),.D(m_axis_outprob_tdata_17_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc951(.Q(acs_prob_tdata_0[6:6]),.D(m_axis_outprob_tdata_17_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc952(.Q(acs_prob_tdata_0[7:7]),.D(m_axis_outprob_tdata_17_0[7:7]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR desc953(.Q(acs_prob_tdata_0[8:8]),.D(m_axis_outprob_tdata_17_0[8:8]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI4QB51));
  FDR m_axis_outdec_tdata_Z(.Q(acs_dec_tdata),.D(m_axis_outprob_tdata_0_sqmuxa_set),.C(aclk),.R(aresetn_i));
  LUT5 desc954(.I0(un4_v_high_s_8_21),.I1(un4_v_low_s_8_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[8:8]));
defparam desc954.INIT=32'hACACFF00;
  LUT5 desc955(.I0(un4_v_high_s_7_21),.I1(un4_v_low_s_7_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[7:7]));
defparam desc955.INIT=32'hACACFF00;
  LUT5 desc956(.I0(un4_v_high_s_6_21),.I1(un4_v_low_s_6_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[6:6]));
defparam desc956.INIT=32'hACACFF00;
  LUT5 desc957(.I0(un4_v_high_s_5_21),.I1(un4_v_low_s_5_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[5:5]));
defparam desc957.INIT=32'hACACFF00;
  LUT5 desc958(.I0(un4_v_high_s_4_21),.I1(un4_v_low_s_4_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[4:4]));
defparam desc958.INIT=32'hACACFF00;
  LUT5 desc959(.I0(un4_v_high_s_3_21),.I1(un4_v_low_s_3_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[3:3]));
defparam desc959.INIT=32'hACACFF00;
  LUT5 desc960(.I0(un4_v_high_s_2_21),.I1(un4_v_low_s_2_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[2:2]));
defparam desc960.INIT=32'hACACFF00;
  LUT5 desc961(.I0(un4_v_high_s_1_21),.I1(un4_v_low_s_1_21),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_0[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[1:1]));
defparam desc961.INIT=32'hACACFF00;
  LUT6 desc962(.I0(acs_prob_tdata_0[0:0]),.I1(acs_prob_tdata_1[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.I5(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_17_0[0:0]));
defparam desc962.INIT=64'h33CC5A5AAAAAAAAA;
  LUT5 m_axis_outdec_tdata_RNO(.I0(acs_dec_tdata),.I1(acs_tvalid),.I2(v_diff_1[8:8]),.I3(un27_s_axis_input_tready_int),.I4(branch_tvalid),.O(m_axis_outprob_tdata_0_sqmuxa_set));
defparam m_axis_outdec_tdata_RNO.INIT=32'hB8F0AAAA;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_0[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_0[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_0[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_0[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_0[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_0[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_0[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_1[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_1[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_1[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_1[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_1[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_1[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_1[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_1[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc963(.I0(acs_prob_tdata_0[0:0]),.I1(acs_prob_tdata_1[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc963.INIT=16'h9669;
  LUT2 desc964(.I0(un4_v_high_s_1_21),.I1(un4_v_low_s_1_21),.O(v_diff_1_axb_1));
defparam desc964.INIT=4'h9;
  LUT2 desc965(.I0(un4_v_high_s_2_21),.I1(un4_v_low_s_2_21),.O(v_diff_1_axb_2));
defparam desc965.INIT=4'h9;
  LUT2 desc966(.I0(un4_v_high_s_3_21),.I1(un4_v_low_s_3_21),.O(v_diff_1_axb_3));
defparam desc966.INIT=4'h9;
  LUT2 desc967(.I0(un4_v_high_s_4_21),.I1(un4_v_low_s_4_21),.O(v_diff_1_axb_4));
defparam desc967.INIT=4'h9;
  LUT2 desc968(.I0(un4_v_high_s_5_21),.I1(un4_v_low_s_5_21),.O(v_diff_1_axb_5));
defparam desc968.INIT=4'h9;
  LUT2 desc969(.I0(un4_v_high_s_6_21),.I1(un4_v_low_s_6_21),.O(v_diff_1_axb_6));
defparam desc969.INIT=4'h9;
  LUT2 desc970(.I0(un4_v_high_s_7_21),.I1(un4_v_low_s_7_21),.O(v_diff_1_axb_7));
defparam desc970.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT2 desc971(.I0(un4_v_high_s_8_21),.I1(un4_v_low_s_8_21),.O(v_diff_1_axb_8));
defparam desc971.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_1[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_0[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT5 desc972(.I0(write_ram_fsm_0_rep1),.I1(write_ram_fsm_4_rep1),.I2(acs_tvalid),.I3(write_ram_fsm[1:1]),.I4(N_1756_1),.O(un1_s_axis_input_tvalid));
defparam desc972.INIT=32'h00100000;
  LUT5 s_axis_inbranch_tlast_d_RNI4QB51_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(acs_tvalid),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI4QB51));
defparam s_axis_inbranch_tlast_d_RNI4QB51_cZ.INIT=32'hD5DD55DD;
  LUT2 desc973(.I0(acs_prob_tdata_0[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam desc973.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(acs_tvalid),.D(s_axis_inbranch_tlast_d_e_lut6_2_O5),.C(aclk),.R(aresetn_i));
  XORCY desc974(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc975(.DI(un4_v_low_s_7_21),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc976(.DI(un4_v_low_s_6_21),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc977(.DI(un4_v_low_s_5_21),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc978(.DI(un4_v_low_s_4_21),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc979(.DI(un4_v_low_s_3_21),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc980(.DI(un4_v_low_s_2_21),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc981(.DI(un4_v_low_s_1_21),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc982(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_21));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_21));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_1[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_21));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_1[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_21));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_1[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_21));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_1[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_21));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_1[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_21));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_1[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_21));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_1[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_1[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_21));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_21));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_0[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_21));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_0[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_21));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_0[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_21));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_0[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_21));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_0[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_21));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_0[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_21));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_0[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_0[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  FDR m_axis_outdec_tlast_Z(.Q(acs_tlast),.D(branch_tlast),.C(aclk),.R(aresetn_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 s_axis_inbranch_tlast_d_RNIIAVE1_o6(.I0(s_axis_inbranch_tlast_d),.I1(acs_tvalid),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIIAVE1_o6.INIT=16'hBAFA;
  LUT4 s_axis_inbranch_tlast_d_RNIIAVE1_o5(.I0(acs_tvalid),.I1(branch_tvalid),.I2(un1_output_accept),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIIAVE1_O5));
defparam s_axis_inbranch_tlast_d_RNIIAVE1_o5.INIT=16'hF8F0;
  LUT4 s_axis_inbranch_tlast_d_e_lut6_2_o6(.I0(acs_tvalid),.I1(branch_tlast),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_0));
defparam s_axis_inbranch_tlast_d_e_lut6_2_o6.INIT=16'h40C0;
  LUT4 s_axis_inbranch_tlast_d_e_lut6_2_o5(.I0(s_axis_inbranch_tlast_d),.I1(acs_tvalid),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_e_lut6_2_O5));
defparam s_axis_inbranch_tlast_d_e_lut6_2_o5.INIT=16'h74F0;
endmodule
module acsZ0_22_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_29,acs_prob_tdata_28,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_46,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,N_1756_1,aresetn,p_desc989_p_O_FD,p_desc990_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1019_p_O_FDRE);
input branch_tlast ;
output [46:46] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_29 ;
input [8:0] acs_prob_tdata_28 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_46 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNINIBL_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIOFM01 ;
wire un4_v_high_s_7_22 ;
wire un4_v_low_s_7_22 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_22 ;
wire un4_v_low_s_8_22 ;
wire un4_v_high_s_6_22 ;
wire un4_v_low_s_6_22 ;
wire un4_v_high_s_5_22 ;
wire un4_v_low_s_5_22 ;
wire un4_v_high_s_4_22 ;
wire un4_v_low_s_4_22 ;
wire un4_v_high_s_3_22 ;
wire un4_v_low_s_3_22 ;
wire un4_v_high_s_2_22 ;
wire un4_v_low_s_2_22 ;
wire un4_v_high_s_1_22 ;
wire un4_v_low_s_1_22 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1908 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc989_p_O_FD ;
input p_desc990_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1019_p_O_FDRE ;
// instances
  FDR desc983(.Q(acs_prob_tdata_46[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  FDR desc984(.Q(acs_prob_tdata_46[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  FDR desc985(.Q(acs_prob_tdata_46[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  FDR desc986(.Q(acs_prob_tdata_46[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  FDR desc987(.Q(acs_prob_tdata_46[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  FDR desc988(.Q(acs_prob_tdata_46[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01));
  p_O_FD desc989(.Q(acs_prob_tdata_46[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc989_p_O_FD));
  p_O_FD desc990(.Q(acs_prob_tdata_46[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc990_p_O_FD));
  LUT6 desc991(.I0(un4_v_high_s_7_22),.I1(un4_v_low_s_7_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOFM01),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc991.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc992(.I0(un4_v_high_s_8_22),.I1(un4_v_low_s_8_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOFM01),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc992.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc993(.I0(un4_v_high_s_6_22),.I1(un4_v_low_s_6_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc993.INIT=32'hACACFF00;
  LUT5 desc994(.I0(un4_v_high_s_5_22),.I1(un4_v_low_s_5_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc994.INIT=32'hACACFF00;
  LUT5 desc995(.I0(un4_v_high_s_4_22),.I1(un4_v_low_s_4_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc995.INIT=32'hACACFF00;
  LUT5 desc996(.I0(un4_v_high_s_3_22),.I1(un4_v_low_s_3_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc996.INIT=32'hACACFF00;
  LUT5 desc997(.I0(un4_v_high_s_2_22),.I1(un4_v_low_s_2_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc997.INIT=32'hACACFF00;
  LUT5 desc998(.I0(un4_v_high_s_1_22),.I1(un4_v_low_s_1_22),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_46[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc998.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[46:46]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc999(.I0(acs_prob_tdata_28[0:0]),.I1(acs_prob_tdata_29[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc999.INIT=16'h9669;
  LUT2 desc1000(.I0(un4_v_high_s_1_22),.I1(un4_v_low_s_1_22),.O(v_diff_1_axb_1));
defparam desc1000.INIT=4'h9;
  LUT2 desc1001(.I0(un4_v_high_s_2_22),.I1(un4_v_low_s_2_22),.O(v_diff_1_axb_2));
defparam desc1001.INIT=4'h9;
  LUT2 desc1002(.I0(un4_v_high_s_3_22),.I1(un4_v_low_s_3_22),.O(v_diff_1_axb_3));
defparam desc1002.INIT=4'h9;
  LUT2 desc1003(.I0(un4_v_high_s_4_22),.I1(un4_v_low_s_4_22),.O(v_diff_1_axb_4));
defparam desc1003.INIT=4'h9;
  LUT2 desc1004(.I0(un4_v_high_s_5_22),.I1(un4_v_low_s_5_22),.O(v_diff_1_axb_5));
defparam desc1004.INIT=4'h9;
  LUT2 desc1005(.I0(un4_v_high_s_6_22),.I1(un4_v_low_s_6_22),.O(v_diff_1_axb_6));
defparam desc1005.INIT=4'h9;
  LUT2 desc1006(.I0(un4_v_high_s_7_22),.I1(un4_v_low_s_7_22),.O(v_diff_1_axb_7));
defparam desc1006.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_28[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_28[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_28[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_28[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_28[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_28[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_28[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_29[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_29[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_29[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_29[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_29[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_29[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_29[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_29[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1007(.I0(acs_prob_tdata_28[0:0]),.I1(acs_prob_tdata_29[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1908));
defparam desc1007.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_29[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_28[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1008(.I0(un4_v_high_s_8_22),.I1(un4_v_low_s_8_22),.O(v_diff_1_axb_8));
defparam desc1008.INIT=4'h9;
  LUT6 desc1009(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1009.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI6DHT(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI6DHT.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIOFM01_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIOFM01));
defparam s_axis_inbranch_tlast_d_RNIOFM01_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_28[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNINIBL_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_22));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_22));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_29[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_22));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_29[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_22));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_29[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_22));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_29[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_22));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_29[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_22));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_29[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_22));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_29[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_29[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_22));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_22));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_28[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_22));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_28[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_22));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_28[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_22));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_28[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_22));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_28[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_22));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_28[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_22));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_28[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_28[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1010(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1011(.DI(un4_v_low_s_7_22),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1012(.DI(un4_v_low_s_6_22),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1013(.DI(un4_v_low_s_5_22),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1014(.DI(un4_v_low_s_4_22),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1015(.DI(un4_v_low_s_3_22),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1016(.DI(un4_v_low_s_2_22),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1017(.DI(un4_v_low_s_1_22),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1018(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1019(.Q(acs_prob_tdata_46[0:0]),.D(N_1908),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOFM01),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1019_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1020(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNINIBL_O6));
defparam desc1020.INIT=16'hF4F0;
  LUT2 desc1021(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1021.INIT=4'h8;
endmodule
module acsZ0_23_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_19,acs_prob_tdata_18,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_9,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1028_p_O_FD,p_desc1029_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1058_p_O_FDRE);
input branch_tlast ;
output [9:9] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_19 ;
input [8:0] acs_prob_tdata_18 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_9 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI42D91_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIML781 ;
wire un4_v_high_s_7_23 ;
wire un4_v_low_s_7_23 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_23 ;
wire un4_v_low_s_8_23 ;
wire un4_v_high_s_6_23 ;
wire un4_v_low_s_6_23 ;
wire un4_v_high_s_5_23 ;
wire un4_v_low_s_5_23 ;
wire un4_v_high_s_4_23 ;
wire un4_v_low_s_4_23 ;
wire un4_v_high_s_3_23 ;
wire un4_v_low_s_3_23 ;
wire un4_v_high_s_2_23 ;
wire un4_v_low_s_2_23 ;
wire un4_v_high_s_1_23 ;
wire un4_v_low_s_1_23 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1888 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1028_p_O_FD ;
input p_desc1029_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1058_p_O_FDRE ;
// instances
  FDR desc1022(.Q(acs_prob_tdata_9[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  FDR desc1023(.Q(acs_prob_tdata_9[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  FDR desc1024(.Q(acs_prob_tdata_9[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  FDR desc1025(.Q(acs_prob_tdata_9[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  FDR desc1026(.Q(acs_prob_tdata_9[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  FDR desc1027(.Q(acs_prob_tdata_9[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781));
  p_O_FD desc1028(.Q(acs_prob_tdata_9[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1028_p_O_FD));
  p_O_FD desc1029(.Q(acs_prob_tdata_9[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1029_p_O_FD));
  LUT6 desc1030(.I0(un4_v_high_s_7_23),.I1(un4_v_low_s_7_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIML781),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1030.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1031(.I0(un4_v_high_s_8_23),.I1(un4_v_low_s_8_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIML781),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1031.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1032(.I0(un4_v_high_s_6_23),.I1(un4_v_low_s_6_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1032.INIT=32'hACACFF00;
  LUT5 desc1033(.I0(un4_v_high_s_5_23),.I1(un4_v_low_s_5_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1033.INIT=32'hACACFF00;
  LUT5 desc1034(.I0(un4_v_high_s_4_23),.I1(un4_v_low_s_4_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1034.INIT=32'hACACFF00;
  LUT5 desc1035(.I0(un4_v_high_s_3_23),.I1(un4_v_low_s_3_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1035.INIT=32'hACACFF00;
  LUT5 desc1036(.I0(un4_v_high_s_2_23),.I1(un4_v_low_s_2_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1036.INIT=32'hACACFF00;
  LUT5 desc1037(.I0(un4_v_high_s_1_23),.I1(un4_v_low_s_1_23),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_9[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1037.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[9:9]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1038(.I0(acs_prob_tdata_18[0:0]),.I1(acs_prob_tdata_19[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1038.INIT=16'h9669;
  LUT2 desc1039(.I0(un4_v_high_s_1_23),.I1(un4_v_low_s_1_23),.O(v_diff_1_axb_1));
defparam desc1039.INIT=4'h9;
  LUT2 desc1040(.I0(un4_v_high_s_2_23),.I1(un4_v_low_s_2_23),.O(v_diff_1_axb_2));
defparam desc1040.INIT=4'h9;
  LUT2 desc1041(.I0(un4_v_high_s_3_23),.I1(un4_v_low_s_3_23),.O(v_diff_1_axb_3));
defparam desc1041.INIT=4'h9;
  LUT2 desc1042(.I0(un4_v_high_s_4_23),.I1(un4_v_low_s_4_23),.O(v_diff_1_axb_4));
defparam desc1042.INIT=4'h9;
  LUT2 desc1043(.I0(un4_v_high_s_5_23),.I1(un4_v_low_s_5_23),.O(v_diff_1_axb_5));
defparam desc1043.INIT=4'h9;
  LUT2 desc1044(.I0(un4_v_high_s_6_23),.I1(un4_v_low_s_6_23),.O(v_diff_1_axb_6));
defparam desc1044.INIT=4'h9;
  LUT2 desc1045(.I0(un4_v_high_s_7_23),.I1(un4_v_low_s_7_23),.O(v_diff_1_axb_7));
defparam desc1045.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_18[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_18[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_18[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_18[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_18[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_18[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_18[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_19[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_19[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_19[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_19[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_19[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_19[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_19[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_19[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1046(.I0(acs_prob_tdata_18[0:0]),.I1(acs_prob_tdata_19[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1888));
defparam desc1046.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_19[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_18[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1047(.I0(un4_v_high_s_8_23),.I1(un4_v_low_s_8_23),.O(v_diff_1_axb_8));
defparam desc1047.INIT=4'h9;
  LUT6 desc1048(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1048.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI4J251(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI4J251.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIML781_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIML781));
defparam s_axis_inbranch_tlast_d_RNIML781_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_18[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI42D91_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_23));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_23));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_19[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_23));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_19[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_23));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_19[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_23));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_19[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_23));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_19[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_23));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_19[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_23));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_19[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_19[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_23));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_23));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_18[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_23));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_18[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_23));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_18[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_23));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_18[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_23));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_18[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_23));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_18[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_23));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_18[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_18[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1049(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1050(.DI(un4_v_low_s_7_23),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1051(.DI(un4_v_low_s_6_23),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1052(.DI(un4_v_low_s_5_23),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1053(.DI(un4_v_low_s_4_23),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1054(.DI(un4_v_low_s_3_23),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1055(.DI(un4_v_low_s_2_23),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1056(.DI(un4_v_low_s_1_23),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1057(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1058(.Q(acs_prob_tdata_9[0:0]),.D(N_1888),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIML781),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1058_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1059(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI42D91_O6));
defparam desc1059.INIT=16'hF4F0;
  LUT2 desc1060(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1060.INIT=4'h8;
endmodule
module acsZ0_24_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_5,acs_prob_tdata_4,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_2,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_4_rep1,N_1756_1,aresetn,p_desc1067_p_O_FD,p_desc1068_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1097_p_O_FDRE);
input branch_tlast ;
output [2:2] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_5 ;
input [8:0] acs_prob_tdata_4 ;
input [1:0] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_2 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_4_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_4_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIF7F41_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI80I91 ;
wire un4_v_high_s_7_24 ;
wire un4_v_low_s_7_24 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_24 ;
wire un4_v_low_s_8_24 ;
wire un4_v_high_s_6_24 ;
wire un4_v_low_s_6_24 ;
wire un4_v_high_s_5_24 ;
wire un4_v_low_s_5_24 ;
wire un4_v_high_s_4_24 ;
wire un4_v_low_s_4_24 ;
wire un4_v_high_s_3_24 ;
wire un4_v_low_s_3_24 ;
wire un4_v_high_s_2_24 ;
wire un4_v_low_s_2_24 ;
wire un4_v_high_s_1_24 ;
wire un4_v_low_s_1_24 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1868 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1067_p_O_FD ;
input p_desc1068_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1097_p_O_FDRE ;
// instances
  FDR desc1061(.Q(acs_prob_tdata_2[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  FDR desc1062(.Q(acs_prob_tdata_2[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  FDR desc1063(.Q(acs_prob_tdata_2[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  FDR desc1064(.Q(acs_prob_tdata_2[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  FDR desc1065(.Q(acs_prob_tdata_2[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  FDR desc1066(.Q(acs_prob_tdata_2[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91));
  p_O_FD desc1067(.Q(acs_prob_tdata_2[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1067_p_O_FD));
  p_O_FD desc1068(.Q(acs_prob_tdata_2[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1068_p_O_FD));
  LUT6 desc1069(.I0(un4_v_high_s_7_24),.I1(un4_v_low_s_7_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI80I91),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1069.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1070(.I0(un4_v_high_s_8_24),.I1(un4_v_low_s_8_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI80I91),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1070.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1071(.I0(un4_v_high_s_6_24),.I1(un4_v_low_s_6_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1071.INIT=32'hACACFF00;
  LUT5 desc1072(.I0(un4_v_high_s_5_24),.I1(un4_v_low_s_5_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1072.INIT=32'hACACFF00;
  LUT5 desc1073(.I0(un4_v_high_s_4_24),.I1(un4_v_low_s_4_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1073.INIT=32'hACACFF00;
  LUT5 desc1074(.I0(un4_v_high_s_3_24),.I1(un4_v_low_s_3_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1074.INIT=32'hACACFF00;
  LUT5 desc1075(.I0(un4_v_high_s_2_24),.I1(un4_v_low_s_2_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1075.INIT=32'hACACFF00;
  LUT5 desc1076(.I0(un4_v_high_s_1_24),.I1(un4_v_low_s_1_24),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_2[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1076.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[2:2]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1077(.I0(acs_prob_tdata_4[0:0]),.I1(acs_prob_tdata_5[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1077.INIT=16'h9669;
  LUT2 desc1078(.I0(un4_v_high_s_1_24),.I1(un4_v_low_s_1_24),.O(v_diff_1_axb_1));
defparam desc1078.INIT=4'h9;
  LUT2 desc1079(.I0(un4_v_high_s_2_24),.I1(un4_v_low_s_2_24),.O(v_diff_1_axb_2));
defparam desc1079.INIT=4'h9;
  LUT2 desc1080(.I0(un4_v_high_s_3_24),.I1(un4_v_low_s_3_24),.O(v_diff_1_axb_3));
defparam desc1080.INIT=4'h9;
  LUT2 desc1081(.I0(un4_v_high_s_4_24),.I1(un4_v_low_s_4_24),.O(v_diff_1_axb_4));
defparam desc1081.INIT=4'h9;
  LUT2 desc1082(.I0(un4_v_high_s_5_24),.I1(un4_v_low_s_5_24),.O(v_diff_1_axb_5));
defparam desc1082.INIT=4'h9;
  LUT2 desc1083(.I0(un4_v_high_s_6_24),.I1(un4_v_low_s_6_24),.O(v_diff_1_axb_6));
defparam desc1083.INIT=4'h9;
  LUT2 desc1084(.I0(un4_v_high_s_7_24),.I1(un4_v_low_s_7_24),.O(v_diff_1_axb_7));
defparam desc1084.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_4[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_4[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_4[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_4[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_4[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_4[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_4[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_5[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_5[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_5[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_5[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_5[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_5[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_5[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_5[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1085(.I0(acs_prob_tdata_4[0:0]),.I1(acs_prob_tdata_5[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1868));
defparam desc1085.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_5[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_4[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1086(.I0(un4_v_high_s_8_24),.I1(un4_v_low_s_8_24),.O(v_diff_1_axb_8));
defparam desc1086.INIT=4'h9;
  LUT6 desc1087(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4_rep1),.I2(write_ram_fsm[0:0]),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1087.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIMTC61(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIMTC61.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI80I91_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI80I91));
defparam s_axis_inbranch_tlast_d_RNI80I91_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_4[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIF7F41_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_24));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_24));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_5[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_24));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_5[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_24));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_5[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_24));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_5[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_24));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_5[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_24));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_5[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_24));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_5[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_5[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_24));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_24));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_4[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_24));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_4[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_24));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_4[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_24));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_4[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_24));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_4[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_24));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_4[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_24));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_4[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_4[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1088(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1089(.DI(un4_v_low_s_7_24),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1090(.DI(un4_v_low_s_6_24),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1091(.DI(un4_v_low_s_5_24),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1092(.DI(un4_v_low_s_4_24),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1093(.DI(un4_v_low_s_3_24),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1094(.DI(un4_v_low_s_2_24),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1095(.DI(un4_v_low_s_1_24),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1096(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1097(.Q(acs_prob_tdata_2[0:0]),.D(N_1868),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI80I91),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1097_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1098(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIF7F41_O6));
defparam desc1098.INIT=16'hF4F0;
  LUT2 desc1099(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1099.INIT=4'h8;
endmodule
module acsZ0_25_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_41,acs_prob_tdata_40,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_52,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,N_1756_1,aresetn,p_desc1106_p_O_FD,p_desc1107_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1136_p_O_FDRE);
input branch_tlast ;
output [52:52] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_41 ;
input [8:0] acs_prob_tdata_40 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_52 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIEJ2S_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNII8GT ;
wire un4_v_high_s_7_25 ;
wire un4_v_low_s_7_25 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_25 ;
wire un4_v_low_s_8_25 ;
wire un4_v_high_s_6_25 ;
wire un4_v_low_s_6_25 ;
wire un4_v_high_s_5_25 ;
wire un4_v_low_s_5_25 ;
wire un4_v_high_s_4_25 ;
wire un4_v_low_s_4_25 ;
wire un4_v_high_s_3_25 ;
wire un4_v_low_s_3_25 ;
wire un4_v_high_s_2_25 ;
wire un4_v_low_s_2_25 ;
wire un4_v_high_s_1_25 ;
wire un4_v_low_s_1_25 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1848 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1106_p_O_FD ;
input p_desc1107_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1136_p_O_FDRE ;
// instances
  FDR desc1100(.Q(acs_prob_tdata_52[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  FDR desc1101(.Q(acs_prob_tdata_52[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  FDR desc1102(.Q(acs_prob_tdata_52[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  FDR desc1103(.Q(acs_prob_tdata_52[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  FDR desc1104(.Q(acs_prob_tdata_52[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  FDR desc1105(.Q(acs_prob_tdata_52[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT));
  p_O_FD desc1106(.Q(acs_prob_tdata_52[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1106_p_O_FD));
  p_O_FD desc1107(.Q(acs_prob_tdata_52[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1107_p_O_FD));
  LUT6 desc1108(.I0(un4_v_high_s_7_25),.I1(un4_v_low_s_7_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII8GT),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1108.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1109(.I0(un4_v_high_s_8_25),.I1(un4_v_low_s_8_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII8GT),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1109.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1110(.I0(un4_v_high_s_6_25),.I1(un4_v_low_s_6_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1110.INIT=32'hACACFF00;
  LUT5 desc1111(.I0(un4_v_high_s_5_25),.I1(un4_v_low_s_5_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1111.INIT=32'hACACFF00;
  LUT5 desc1112(.I0(un4_v_high_s_4_25),.I1(un4_v_low_s_4_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1112.INIT=32'hACACFF00;
  LUT5 desc1113(.I0(un4_v_high_s_3_25),.I1(un4_v_low_s_3_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1113.INIT=32'hACACFF00;
  LUT5 desc1114(.I0(un4_v_high_s_2_25),.I1(un4_v_low_s_2_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1114.INIT=32'hACACFF00;
  LUT5 desc1115(.I0(un4_v_high_s_1_25),.I1(un4_v_low_s_1_25),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_52[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1115.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[52:52]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1116(.I0(acs_prob_tdata_40[0:0]),.I1(acs_prob_tdata_41[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1116.INIT=16'h9669;
  LUT2 desc1117(.I0(un4_v_high_s_1_25),.I1(un4_v_low_s_1_25),.O(v_diff_1_axb_1));
defparam desc1117.INIT=4'h9;
  LUT2 desc1118(.I0(un4_v_high_s_2_25),.I1(un4_v_low_s_2_25),.O(v_diff_1_axb_2));
defparam desc1118.INIT=4'h9;
  LUT2 desc1119(.I0(un4_v_high_s_3_25),.I1(un4_v_low_s_3_25),.O(v_diff_1_axb_3));
defparam desc1119.INIT=4'h9;
  LUT2 desc1120(.I0(un4_v_high_s_4_25),.I1(un4_v_low_s_4_25),.O(v_diff_1_axb_4));
defparam desc1120.INIT=4'h9;
  LUT2 desc1121(.I0(un4_v_high_s_5_25),.I1(un4_v_low_s_5_25),.O(v_diff_1_axb_5));
defparam desc1121.INIT=4'h9;
  LUT2 desc1122(.I0(un4_v_high_s_6_25),.I1(un4_v_low_s_6_25),.O(v_diff_1_axb_6));
defparam desc1122.INIT=4'h9;
  LUT2 desc1123(.I0(un4_v_high_s_7_25),.I1(un4_v_low_s_7_25),.O(v_diff_1_axb_7));
defparam desc1123.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_40[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_40[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_40[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_40[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_40[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_40[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_40[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_41[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_41[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_41[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_41[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_41[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_41[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_41[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_41[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1124(.I0(acs_prob_tdata_40[0:0]),.I1(acs_prob_tdata_41[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1848));
defparam desc1124.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_41[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_40[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1125(.I0(un4_v_high_s_8_25),.I1(un4_v_low_s_8_25),.O(v_diff_1_axb_8));
defparam desc1125.INIT=4'h9;
  LUT6 desc1126(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1126.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI06BQ(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI06BQ.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNII8GT_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNII8GT));
defparam s_axis_inbranch_tlast_d_RNII8GT_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_40[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIEJ2S_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_25));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_25));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_41[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_25));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_41[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_25));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_41[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_25));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_41[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_25));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_41[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_25));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_41[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_25));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_41[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_41[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_25));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_25));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_40[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_25));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_40[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_25));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_40[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_25));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_40[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_25));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_40[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_25));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_40[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_25));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_40[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_40[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1127(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1128(.DI(un4_v_low_s_7_25),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1129(.DI(un4_v_low_s_6_25),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1130(.DI(un4_v_low_s_5_25),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1131(.DI(un4_v_low_s_4_25),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1132(.DI(un4_v_low_s_3_25),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1133(.DI(un4_v_low_s_2_25),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1134(.DI(un4_v_low_s_1_25),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1135(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1136(.Q(acs_prob_tdata_52[0:0]),.D(N_1848),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII8GT),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1136_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1137(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIEJ2S_O6));
defparam desc1137.INIT=16'hF4F0;
  LUT2 desc1138(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1138.INIT=4'h8;
endmodule
module acsZ0_26_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_21,acs_prob_tdata_20,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_10,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1145_p_O_FD,p_desc1146_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1175_p_O_FDRE);
input branch_tlast ;
output [10:10] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_21 ;
input [8:0] acs_prob_tdata_20 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_10 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIS2CR_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI6EH41 ;
wire un4_v_high_s_7_26 ;
wire un4_v_low_s_7_26 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_26 ;
wire un4_v_low_s_8_26 ;
wire un4_v_high_s_6_26 ;
wire un4_v_low_s_6_26 ;
wire un4_v_high_s_5_26 ;
wire un4_v_low_s_5_26 ;
wire un4_v_high_s_4_26 ;
wire un4_v_low_s_4_26 ;
wire un4_v_high_s_3_26 ;
wire un4_v_low_s_3_26 ;
wire un4_v_high_s_2_26 ;
wire un4_v_low_s_2_26 ;
wire un4_v_high_s_1_26 ;
wire un4_v_low_s_1_26 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1828 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1145_p_O_FD ;
input p_desc1146_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1175_p_O_FDRE ;
// instances
  FDR desc1139(.Q(acs_prob_tdata_10[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  FDR desc1140(.Q(acs_prob_tdata_10[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  FDR desc1141(.Q(acs_prob_tdata_10[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  FDR desc1142(.Q(acs_prob_tdata_10[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  FDR desc1143(.Q(acs_prob_tdata_10[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  FDR desc1144(.Q(acs_prob_tdata_10[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41));
  p_O_FD desc1145(.Q(acs_prob_tdata_10[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1145_p_O_FD));
  p_O_FD desc1146(.Q(acs_prob_tdata_10[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1146_p_O_FD));
  LUT6 desc1147(.I0(un4_v_high_s_7_26),.I1(un4_v_low_s_7_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI6EH41),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1147.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1148(.I0(un4_v_high_s_8_26),.I1(un4_v_low_s_8_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI6EH41),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1148.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1149(.I0(un4_v_high_s_6_26),.I1(un4_v_low_s_6_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1149.INIT=32'hACACFF00;
  LUT5 desc1150(.I0(un4_v_high_s_5_26),.I1(un4_v_low_s_5_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1150.INIT=32'hACACFF00;
  LUT5 desc1151(.I0(un4_v_high_s_4_26),.I1(un4_v_low_s_4_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1151.INIT=32'hACACFF00;
  LUT5 desc1152(.I0(un4_v_high_s_3_26),.I1(un4_v_low_s_3_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1152.INIT=32'hACACFF00;
  LUT5 desc1153(.I0(un4_v_high_s_2_26),.I1(un4_v_low_s_2_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1153.INIT=32'hACACFF00;
  LUT5 desc1154(.I0(un4_v_high_s_1_26),.I1(un4_v_low_s_1_26),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_10[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1154.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[10:10]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1155(.I0(acs_prob_tdata_20[0:0]),.I1(acs_prob_tdata_21[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1155.INIT=16'h9669;
  LUT2 desc1156(.I0(un4_v_high_s_1_26),.I1(un4_v_low_s_1_26),.O(v_diff_1_axb_1));
defparam desc1156.INIT=4'h9;
  LUT2 desc1157(.I0(un4_v_high_s_2_26),.I1(un4_v_low_s_2_26),.O(v_diff_1_axb_2));
defparam desc1157.INIT=4'h9;
  LUT2 desc1158(.I0(un4_v_high_s_3_26),.I1(un4_v_low_s_3_26),.O(v_diff_1_axb_3));
defparam desc1158.INIT=4'h9;
  LUT2 desc1159(.I0(un4_v_high_s_4_26),.I1(un4_v_low_s_4_26),.O(v_diff_1_axb_4));
defparam desc1159.INIT=4'h9;
  LUT2 desc1160(.I0(un4_v_high_s_5_26),.I1(un4_v_low_s_5_26),.O(v_diff_1_axb_5));
defparam desc1160.INIT=4'h9;
  LUT2 desc1161(.I0(un4_v_high_s_6_26),.I1(un4_v_low_s_6_26),.O(v_diff_1_axb_6));
defparam desc1161.INIT=4'h9;
  LUT2 desc1162(.I0(un4_v_high_s_7_26),.I1(un4_v_low_s_7_26),.O(v_diff_1_axb_7));
defparam desc1162.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_20[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_20[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_20[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_20[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_20[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_20[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_20[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_21[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_21[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_21[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_21[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_21[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_21[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_21[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_21[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1163(.I0(acs_prob_tdata_20[0:0]),.I1(acs_prob_tdata_21[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1828));
defparam desc1163.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_21[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_20[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1164(.I0(un4_v_high_s_8_26),.I1(un4_v_low_s_8_26),.O(v_diff_1_axb_8));
defparam desc1164.INIT=4'h9;
  LUT6 desc1165(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1165.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIKBC11(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIKBC11.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI6EH41_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI6EH41));
defparam s_axis_inbranch_tlast_d_RNI6EH41_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_20[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIS2CR_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_26));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_26));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_21[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_26));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_21[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_26));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_21[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_26));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_21[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_26));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_21[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_26));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_21[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_26));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_21[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_21[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_26));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_26));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_20[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_26));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_20[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_26));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_20[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_26));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_20[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_26));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_20[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_26));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_20[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_26));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_20[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_20[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1166(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1167(.DI(un4_v_low_s_7_26),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1168(.DI(un4_v_low_s_6_26),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1169(.DI(un4_v_low_s_5_26),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1170(.DI(un4_v_low_s_4_26),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1171(.DI(un4_v_low_s_3_26),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1172(.DI(un4_v_low_s_2_26),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1173(.DI(un4_v_low_s_1_26),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1174(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1175(.Q(acs_prob_tdata_10[0:0]),.D(N_1828),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI6EH41),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1175_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1176(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIS2CR_O6));
defparam desc1176.INIT=16'hF4F0;
  LUT2 desc1177(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1177.INIT=4'h8;
endmodule
module acsZ0_27_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_45,acs_prob_tdata_44,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_22,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1184_p_O_FD,p_desc1185_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1214_p_O_FDRE);
input branch_tlast ;
output [22:22] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_45 ;
input [8:0] acs_prob_tdata_44 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_22 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI58141_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNICPTD1 ;
wire un4_v_high_s_7_27 ;
wire un4_v_low_s_7_27 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_27 ;
wire un4_v_low_s_8_27 ;
wire un4_v_high_s_6_27 ;
wire un4_v_low_s_6_27 ;
wire un4_v_high_s_5_27 ;
wire un4_v_low_s_5_27 ;
wire un4_v_high_s_4_27 ;
wire un4_v_low_s_4_27 ;
wire un4_v_high_s_3_27 ;
wire un4_v_low_s_3_27 ;
wire un4_v_high_s_2_27 ;
wire un4_v_low_s_2_27 ;
wire un4_v_high_s_1_27 ;
wire un4_v_low_s_1_27 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1808 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1184_p_O_FD ;
input p_desc1185_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1214_p_O_FDRE ;
// instances
  FDR desc1178(.Q(acs_prob_tdata_22[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  FDR desc1179(.Q(acs_prob_tdata_22[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  FDR desc1180(.Q(acs_prob_tdata_22[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  FDR desc1181(.Q(acs_prob_tdata_22[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  FDR desc1182(.Q(acs_prob_tdata_22[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  FDR desc1183(.Q(acs_prob_tdata_22[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1));
  p_O_FD desc1184(.Q(acs_prob_tdata_22[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1184_p_O_FD));
  p_O_FD desc1185(.Q(acs_prob_tdata_22[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1185_p_O_FD));
  LUT6 desc1186(.I0(un4_v_high_s_7_27),.I1(un4_v_low_s_7_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICPTD1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1186.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1187(.I0(un4_v_high_s_8_27),.I1(un4_v_low_s_8_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICPTD1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1187.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1188(.I0(un4_v_high_s_6_27),.I1(un4_v_low_s_6_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1188.INIT=32'hACACFF00;
  LUT5 desc1189(.I0(un4_v_high_s_5_27),.I1(un4_v_low_s_5_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1189.INIT=32'hACACFF00;
  LUT5 desc1190(.I0(un4_v_high_s_4_27),.I1(un4_v_low_s_4_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1190.INIT=32'hACACFF00;
  LUT5 desc1191(.I0(un4_v_high_s_3_27),.I1(un4_v_low_s_3_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1191.INIT=32'hACACFF00;
  LUT5 desc1192(.I0(un4_v_high_s_2_27),.I1(un4_v_low_s_2_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1192.INIT=32'hACACFF00;
  LUT5 desc1193(.I0(un4_v_high_s_1_27),.I1(un4_v_low_s_1_27),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_22[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1193.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[22:22]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_44[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_44[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_44[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_44[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_44[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_44[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_44[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_45[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_45[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_45[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_45[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_45[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_45[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_45[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_45[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1194(.I0(acs_prob_tdata_44[0:0]),.I1(acs_prob_tdata_45[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1194.INIT=16'h9669;
  LUT2 desc1195(.I0(un4_v_high_s_1_27),.I1(un4_v_low_s_1_27),.O(v_diff_1_axb_1));
defparam desc1195.INIT=4'h9;
  LUT2 desc1196(.I0(un4_v_high_s_2_27),.I1(un4_v_low_s_2_27),.O(v_diff_1_axb_2));
defparam desc1196.INIT=4'h9;
  LUT2 desc1197(.I0(un4_v_high_s_3_27),.I1(un4_v_low_s_3_27),.O(v_diff_1_axb_3));
defparam desc1197.INIT=4'h9;
  LUT2 desc1198(.I0(un4_v_high_s_4_27),.I1(un4_v_low_s_4_27),.O(v_diff_1_axb_4));
defparam desc1198.INIT=4'h9;
  LUT2 desc1199(.I0(un4_v_high_s_5_27),.I1(un4_v_low_s_5_27),.O(v_diff_1_axb_5));
defparam desc1199.INIT=4'h9;
  LUT2 desc1200(.I0(un4_v_high_s_6_27),.I1(un4_v_low_s_6_27),.O(v_diff_1_axb_6));
defparam desc1200.INIT=4'h9;
  LUT2 desc1201(.I0(un4_v_high_s_7_27),.I1(un4_v_low_s_7_27),.O(v_diff_1_axb_7));
defparam desc1201.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1202(.I0(acs_prob_tdata_44[0:0]),.I1(acs_prob_tdata_45[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1808));
defparam desc1202.INIT=32'h33CC5A5A;
  LUT2 desc1203(.I0(un4_v_high_s_8_27),.I1(un4_v_low_s_8_27),.O(v_diff_1_axb_8));
defparam desc1203.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_45[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_44[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1204(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1204.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIQMOA1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQMOA1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNICPTD1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNICPTD1));
defparam s_axis_inbranch_tlast_d_RNICPTD1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_44[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI58141_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1205(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1206(.DI(un4_v_low_s_7_27),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1207(.DI(un4_v_low_s_6_27),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1208(.DI(un4_v_low_s_5_27),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1209(.DI(un4_v_low_s_4_27),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1210(.DI(un4_v_low_s_3_27),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1211(.DI(un4_v_low_s_2_27),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1212(.DI(un4_v_low_s_1_27),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1213(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_27));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_27));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_45[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_27));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_45[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_27));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_45[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_27));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_45[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_27));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_45[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_27));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_45[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_27));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_45[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_45[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_27));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_27));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_44[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_27));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_44[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_27));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_44[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_27));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_44[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_27));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_44[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_27));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_44[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_27));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_44[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_44[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1214(.Q(acs_prob_tdata_22[0:0]),.D(N_1808),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICPTD1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1214_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1215(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI58141_O6));
defparam desc1215.INIT=16'hF4F0;
  LUT2 desc1216(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1216.INIT=4'h8;
endmodule
module acsZ0_28_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_15,acs_prob_tdata_14,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_7,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1223_p_O_FD,p_desc1224_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1253_p_O_FDRE);
input branch_tlast ;
output [7:7] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_15 ;
input [8:0] acs_prob_tdata_14 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_7 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIULD31_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIIF141 ;
wire un4_v_high_s_7_28 ;
wire un4_v_low_s_7_28 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_28 ;
wire un4_v_low_s_8_28 ;
wire un4_v_high_s_6_28 ;
wire un4_v_low_s_6_28 ;
wire un4_v_high_s_5_28 ;
wire un4_v_low_s_5_28 ;
wire un4_v_high_s_4_28 ;
wire un4_v_low_s_4_28 ;
wire un4_v_high_s_3_28 ;
wire un4_v_low_s_3_28 ;
wire un4_v_high_s_2_28 ;
wire un4_v_low_s_2_28 ;
wire un4_v_high_s_1_28 ;
wire un4_v_low_s_1_28 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1788 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1223_p_O_FD ;
input p_desc1224_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1253_p_O_FDRE ;
// instances
  FDR desc1217(.Q(acs_prob_tdata_7[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  FDR desc1218(.Q(acs_prob_tdata_7[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  FDR desc1219(.Q(acs_prob_tdata_7[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  FDR desc1220(.Q(acs_prob_tdata_7[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  FDR desc1221(.Q(acs_prob_tdata_7[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  FDR desc1222(.Q(acs_prob_tdata_7[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141));
  p_O_FD desc1223(.Q(acs_prob_tdata_7[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1223_p_O_FD));
  p_O_FD desc1224(.Q(acs_prob_tdata_7[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1224_p_O_FD));
  LUT6 desc1225(.I0(un4_v_high_s_7_28),.I1(un4_v_low_s_7_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIIF141),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1225.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1226(.I0(un4_v_high_s_8_28),.I1(un4_v_low_s_8_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIIF141),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1226.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1227(.I0(un4_v_high_s_6_28),.I1(un4_v_low_s_6_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1227.INIT=32'hACACFF00;
  LUT5 desc1228(.I0(un4_v_high_s_5_28),.I1(un4_v_low_s_5_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1228.INIT=32'hACACFF00;
  LUT5 desc1229(.I0(un4_v_high_s_4_28),.I1(un4_v_low_s_4_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1229.INIT=32'hACACFF00;
  LUT5 desc1230(.I0(un4_v_high_s_3_28),.I1(un4_v_low_s_3_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1230.INIT=32'hACACFF00;
  LUT5 desc1231(.I0(un4_v_high_s_2_28),.I1(un4_v_low_s_2_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1231.INIT=32'hACACFF00;
  LUT5 desc1232(.I0(un4_v_high_s_1_28),.I1(un4_v_low_s_1_28),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_7[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1232.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[7:7]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_14[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_14[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_14[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_14[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_14[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_14[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_14[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_15[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_15[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_15[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_15[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_15[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_15[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_15[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_15[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1233(.I0(acs_prob_tdata_14[0:0]),.I1(acs_prob_tdata_15[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1233.INIT=16'h9669;
  LUT2 desc1234(.I0(un4_v_high_s_1_28),.I1(un4_v_low_s_1_28),.O(v_diff_1_axb_1));
defparam desc1234.INIT=4'h9;
  LUT2 desc1235(.I0(un4_v_high_s_2_28),.I1(un4_v_low_s_2_28),.O(v_diff_1_axb_2));
defparam desc1235.INIT=4'h9;
  LUT2 desc1236(.I0(un4_v_high_s_3_28),.I1(un4_v_low_s_3_28),.O(v_diff_1_axb_3));
defparam desc1236.INIT=4'h9;
  LUT2 desc1237(.I0(un4_v_high_s_4_28),.I1(un4_v_low_s_4_28),.O(v_diff_1_axb_4));
defparam desc1237.INIT=4'h9;
  LUT2 desc1238(.I0(un4_v_high_s_5_28),.I1(un4_v_low_s_5_28),.O(v_diff_1_axb_5));
defparam desc1238.INIT=4'h9;
  LUT2 desc1239(.I0(un4_v_high_s_6_28),.I1(un4_v_low_s_6_28),.O(v_diff_1_axb_6));
defparam desc1239.INIT=4'h9;
  LUT2 desc1240(.I0(un4_v_high_s_7_28),.I1(un4_v_low_s_7_28),.O(v_diff_1_axb_7));
defparam desc1240.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1241(.I0(acs_prob_tdata_14[0:0]),.I1(acs_prob_tdata_15[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1788));
defparam desc1241.INIT=32'h3C3C55AA;
  LUT2 desc1242(.I0(un4_v_high_s_8_28),.I1(un4_v_low_s_8_28),.O(v_diff_1_axb_8));
defparam desc1242.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_15[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_14[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1243(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1243.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI0DS01(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI0DS01.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIIF141_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIIF141));
defparam s_axis_inbranch_tlast_d_RNIIF141_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_14[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIULD31_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1244(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1245(.DI(un4_v_low_s_7_28),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1246(.DI(un4_v_low_s_6_28),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1247(.DI(un4_v_low_s_5_28),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1248(.DI(un4_v_low_s_4_28),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1249(.DI(un4_v_low_s_3_28),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1250(.DI(un4_v_low_s_2_28),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1251(.DI(un4_v_low_s_1_28),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1252(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_28));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_28));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_15[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_28));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_15[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_28));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_15[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_28));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_15[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_28));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_15[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_28));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_15[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_28));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_15[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_15[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_28));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_28));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_14[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_28));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_14[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_28));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_14[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_28));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_14[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_28));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_14[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_28));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_14[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_28));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_14[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_14[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1253(.Q(acs_prob_tdata_7[0:0]),.D(N_1788),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIIF141),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1253_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1254(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIULD31_O6));
defparam desc1254.INIT=16'hF4F0;
  LUT2 desc1255(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1255.INIT=4'h8;
endmodule
module acsZ0_29_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_15,acs_prob_tdata_14,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_39,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc1262_p_O_FD,p_desc1263_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1292_p_O_FDRE);
input branch_tlast ;
output [39:39] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_15 ;
input [8:0] acs_prob_tdata_14 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_39 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNITRKR_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNISJP11 ;
wire un4_v_high_s_7_29 ;
wire un4_v_low_s_7_29 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_29 ;
wire un4_v_low_s_8_29 ;
wire un4_v_high_s_6_29 ;
wire un4_v_low_s_6_29 ;
wire un4_v_high_s_5_29 ;
wire un4_v_low_s_5_29 ;
wire un4_v_high_s_4_29 ;
wire un4_v_low_s_4_29 ;
wire un4_v_high_s_3_29 ;
wire un4_v_low_s_3_29 ;
wire un4_v_high_s_2_29 ;
wire un4_v_low_s_2_29 ;
wire un4_v_high_s_1_29 ;
wire un4_v_low_s_1_29 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1768 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1262_p_O_FD ;
input p_desc1263_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1292_p_O_FDRE ;
// instances
  FDR desc1256(.Q(acs_prob_tdata_39[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  FDR desc1257(.Q(acs_prob_tdata_39[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  FDR desc1258(.Q(acs_prob_tdata_39[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  FDR desc1259(.Q(acs_prob_tdata_39[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  FDR desc1260(.Q(acs_prob_tdata_39[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  FDR desc1261(.Q(acs_prob_tdata_39[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11));
  p_O_FD desc1262(.Q(acs_prob_tdata_39[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1262_p_O_FD));
  p_O_FD desc1263(.Q(acs_prob_tdata_39[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1263_p_O_FD));
  LUT6 desc1264(.I0(un4_v_high_s_7_29),.I1(un4_v_low_s_7_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISJP11),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1264.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1265(.I0(un4_v_high_s_8_29),.I1(un4_v_low_s_8_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISJP11),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1265.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1266(.I0(un4_v_high_s_6_29),.I1(un4_v_low_s_6_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1266.INIT=32'hACACFF00;
  LUT5 desc1267(.I0(un4_v_high_s_5_29),.I1(un4_v_low_s_5_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1267.INIT=32'hACACFF00;
  LUT5 desc1268(.I0(un4_v_high_s_4_29),.I1(un4_v_low_s_4_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1268.INIT=32'hACACFF00;
  LUT5 desc1269(.I0(un4_v_high_s_3_29),.I1(un4_v_low_s_3_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1269.INIT=32'hACACFF00;
  LUT5 desc1270(.I0(un4_v_high_s_2_29),.I1(un4_v_low_s_2_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1270.INIT=32'hACACFF00;
  LUT5 desc1271(.I0(un4_v_high_s_1_29),.I1(un4_v_low_s_1_29),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_39[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1271.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[39:39]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1272(.I0(acs_prob_tdata_14[0:0]),.I1(acs_prob_tdata_15[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1272.INIT=16'h9669;
  LUT2 desc1273(.I0(un4_v_high_s_1_29),.I1(un4_v_low_s_1_29),.O(v_diff_1_axb_1));
defparam desc1273.INIT=4'h9;
  LUT2 desc1274(.I0(un4_v_high_s_2_29),.I1(un4_v_low_s_2_29),.O(v_diff_1_axb_2));
defparam desc1274.INIT=4'h9;
  LUT2 desc1275(.I0(un4_v_high_s_3_29),.I1(un4_v_low_s_3_29),.O(v_diff_1_axb_3));
defparam desc1275.INIT=4'h9;
  LUT2 desc1276(.I0(un4_v_high_s_4_29),.I1(un4_v_low_s_4_29),.O(v_diff_1_axb_4));
defparam desc1276.INIT=4'h9;
  LUT2 desc1277(.I0(un4_v_high_s_5_29),.I1(un4_v_low_s_5_29),.O(v_diff_1_axb_5));
defparam desc1277.INIT=4'h9;
  LUT2 desc1278(.I0(un4_v_high_s_6_29),.I1(un4_v_low_s_6_29),.O(v_diff_1_axb_6));
defparam desc1278.INIT=4'h9;
  LUT2 desc1279(.I0(un4_v_high_s_7_29),.I1(un4_v_low_s_7_29),.O(v_diff_1_axb_7));
defparam desc1279.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_14[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_14[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_14[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_14[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_14[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_14[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_14[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_15[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_15[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_15[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_15[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_15[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_15[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_15[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_15[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1280(.I0(acs_prob_tdata_14[0:0]),.I1(acs_prob_tdata_15[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1768));
defparam desc1280.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_15[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_14[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1281(.I0(un4_v_high_s_8_29),.I1(un4_v_low_s_8_29),.O(v_diff_1_axb_8));
defparam desc1281.INIT=4'h9;
  LUT6 desc1282(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1282.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIAHKU(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIAHKU.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNISJP11_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNISJP11));
defparam s_axis_inbranch_tlast_d_RNISJP11_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_14[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNITRKR_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_29));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_29));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_15[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_29));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_15[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_29));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_15[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_29));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_15[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_29));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_15[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_29));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_15[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_29));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_15[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_15[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_29));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_29));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_14[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_29));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_14[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_29));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_14[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_29));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_14[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_29));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_14[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_29));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_14[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_29));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_14[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_14[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1283(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1284(.DI(un4_v_low_s_7_29),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1285(.DI(un4_v_low_s_6_29),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1286(.DI(un4_v_low_s_5_29),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1287(.DI(un4_v_low_s_4_29),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1288(.DI(un4_v_low_s_3_29),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1289(.DI(un4_v_low_s_2_29),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1290(.DI(un4_v_low_s_1_29),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1291(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1292(.Q(acs_prob_tdata_39[0:0]),.D(N_1768),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISJP11),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1292_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1293(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNITRKR_O6));
defparam desc1293.INIT=16'hF4F0;
  LUT2 desc1294(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1294.INIT=4'h8;
endmodule
module acsZ0_30_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_39,acs_prob_tdata_38,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_51,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,N_1756_1,aresetn,p_desc1301_p_O_FD,p_desc1302_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1331_p_O_FDRE);
input branch_tlast ;
output [51:51] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_39 ;
input [8:0] acs_prob_tdata_38 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_51 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIBT291_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIG5DB1 ;
wire un4_v_high_s_7_30 ;
wire un4_v_low_s_7_30 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_30 ;
wire un4_v_low_s_8_30 ;
wire un4_v_high_s_6_30 ;
wire un4_v_low_s_6_30 ;
wire un4_v_high_s_5_30 ;
wire un4_v_low_s_5_30 ;
wire un4_v_high_s_4_30 ;
wire un4_v_low_s_4_30 ;
wire un4_v_high_s_3_30 ;
wire un4_v_low_s_3_30 ;
wire un4_v_high_s_2_30 ;
wire un4_v_low_s_2_30 ;
wire un4_v_high_s_1_30 ;
wire un4_v_low_s_1_30 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1748 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1301_p_O_FD ;
input p_desc1302_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1331_p_O_FDRE ;
// instances
  FDR desc1295(.Q(acs_prob_tdata_51[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  FDR desc1296(.Q(acs_prob_tdata_51[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  FDR desc1297(.Q(acs_prob_tdata_51[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  FDR desc1298(.Q(acs_prob_tdata_51[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  FDR desc1299(.Q(acs_prob_tdata_51[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  FDR desc1300(.Q(acs_prob_tdata_51[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1));
  p_O_FD desc1301(.Q(acs_prob_tdata_51[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1301_p_O_FD));
  p_O_FD desc1302(.Q(acs_prob_tdata_51[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1302_p_O_FD));
  LUT6 desc1303(.I0(un4_v_high_s_7_30),.I1(un4_v_low_s_7_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG5DB1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1303.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1304(.I0(un4_v_high_s_8_30),.I1(un4_v_low_s_8_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG5DB1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1304.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1305(.I0(un4_v_high_s_6_30),.I1(un4_v_low_s_6_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1305.INIT=32'hACACFF00;
  LUT5 desc1306(.I0(un4_v_high_s_5_30),.I1(un4_v_low_s_5_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1306.INIT=32'hACACFF00;
  LUT5 desc1307(.I0(un4_v_high_s_4_30),.I1(un4_v_low_s_4_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1307.INIT=32'hACACFF00;
  LUT5 desc1308(.I0(un4_v_high_s_3_30),.I1(un4_v_low_s_3_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1308.INIT=32'hACACFF00;
  LUT5 desc1309(.I0(un4_v_high_s_2_30),.I1(un4_v_low_s_2_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1309.INIT=32'hACACFF00;
  LUT5 desc1310(.I0(un4_v_high_s_1_30),.I1(un4_v_low_s_1_30),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_51[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1310.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[51:51]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1311(.I0(acs_prob_tdata_38[0:0]),.I1(acs_prob_tdata_39[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1311.INIT=16'h9669;
  LUT2 desc1312(.I0(un4_v_high_s_1_30),.I1(un4_v_low_s_1_30),.O(v_diff_1_axb_1));
defparam desc1312.INIT=4'h9;
  LUT2 desc1313(.I0(un4_v_high_s_2_30),.I1(un4_v_low_s_2_30),.O(v_diff_1_axb_2));
defparam desc1313.INIT=4'h9;
  LUT2 desc1314(.I0(un4_v_high_s_3_30),.I1(un4_v_low_s_3_30),.O(v_diff_1_axb_3));
defparam desc1314.INIT=4'h9;
  LUT2 desc1315(.I0(un4_v_high_s_4_30),.I1(un4_v_low_s_4_30),.O(v_diff_1_axb_4));
defparam desc1315.INIT=4'h9;
  LUT2 desc1316(.I0(un4_v_high_s_5_30),.I1(un4_v_low_s_5_30),.O(v_diff_1_axb_5));
defparam desc1316.INIT=4'h9;
  LUT2 desc1317(.I0(un4_v_high_s_6_30),.I1(un4_v_low_s_6_30),.O(v_diff_1_axb_6));
defparam desc1317.INIT=4'h9;
  LUT2 desc1318(.I0(un4_v_high_s_7_30),.I1(un4_v_low_s_7_30),.O(v_diff_1_axb_7));
defparam desc1318.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_38[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_38[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_38[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_38[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_38[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_38[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_38[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_39[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_39[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_39[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_39[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_39[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_39[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_39[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_39[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1319(.I0(acs_prob_tdata_38[0:0]),.I1(acs_prob_tdata_39[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1748));
defparam desc1319.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_39[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_38[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1320(.I0(un4_v_high_s_8_30),.I1(un4_v_low_s_8_30),.O(v_diff_1_axb_8));
defparam desc1320.INIT=4'h9;
  LUT6 desc1321(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1321.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIU2881(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIU2881.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIG5DB1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIG5DB1));
defparam s_axis_inbranch_tlast_d_RNIG5DB1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_38[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIBT291_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_30));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_30));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_39[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_30));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_39[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_30));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_39[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_30));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_39[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_30));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_39[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_30));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_39[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_30));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_39[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_39[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_30));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_30));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_38[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_30));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_38[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_30));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_38[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_30));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_38[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_30));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_38[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_30));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_38[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_30));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_38[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_38[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1322(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1323(.DI(un4_v_low_s_7_30),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1324(.DI(un4_v_low_s_6_30),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1325(.DI(un4_v_low_s_5_30),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1326(.DI(un4_v_low_s_4_30),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1327(.DI(un4_v_low_s_3_30),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1328(.DI(un4_v_low_s_2_30),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1329(.DI(un4_v_low_s_1_30),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1330(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1331(.Q(acs_prob_tdata_51[0:0]),.D(N_1748),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG5DB1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1331_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1332(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIBT291_O6));
defparam desc1332.INIT=16'hF4F0;
  LUT2 desc1333(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1333.INIT=4'h8;
endmodule
module acsZ0_31_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_9,acs_prob_tdata_8,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_36,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc1340_p_O_FD,p_desc1341_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1370_p_O_FDRE);
input branch_tlast ;
output [36:36] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_9 ;
input [8:0] acs_prob_tdata_8 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_36 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIKPL21_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIMAGB1 ;
wire un4_v_high_s_7_31 ;
wire un4_v_low_s_7_31 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_31 ;
wire un4_v_low_s_8_31 ;
wire un4_v_high_s_6_31 ;
wire un4_v_low_s_6_31 ;
wire un4_v_high_s_5_31 ;
wire un4_v_low_s_5_31 ;
wire un4_v_high_s_4_31 ;
wire un4_v_low_s_4_31 ;
wire un4_v_high_s_3_31 ;
wire un4_v_low_s_3_31 ;
wire un4_v_high_s_2_31 ;
wire un4_v_low_s_2_31 ;
wire un4_v_high_s_1_31 ;
wire un4_v_low_s_1_31 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1728 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1340_p_O_FD ;
input p_desc1341_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1370_p_O_FDRE ;
// instances
  FDR desc1334(.Q(acs_prob_tdata_36[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  FDR desc1335(.Q(acs_prob_tdata_36[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  FDR desc1336(.Q(acs_prob_tdata_36[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  FDR desc1337(.Q(acs_prob_tdata_36[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  FDR desc1338(.Q(acs_prob_tdata_36[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  FDR desc1339(.Q(acs_prob_tdata_36[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1));
  p_O_FD desc1340(.Q(acs_prob_tdata_36[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1340_p_O_FD));
  p_O_FD desc1341(.Q(acs_prob_tdata_36[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1341_p_O_FD));
  LUT6 desc1342(.I0(un4_v_high_s_7_31),.I1(un4_v_low_s_7_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMAGB1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1342.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1343(.I0(un4_v_high_s_8_31),.I1(un4_v_low_s_8_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMAGB1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1343.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1344(.I0(un4_v_high_s_6_31),.I1(un4_v_low_s_6_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1344.INIT=32'hACACFF00;
  LUT5 desc1345(.I0(un4_v_high_s_5_31),.I1(un4_v_low_s_5_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1345.INIT=32'hACACFF00;
  LUT5 desc1346(.I0(un4_v_high_s_4_31),.I1(un4_v_low_s_4_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1346.INIT=32'hACACFF00;
  LUT5 desc1347(.I0(un4_v_high_s_3_31),.I1(un4_v_low_s_3_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1347.INIT=32'hACACFF00;
  LUT5 desc1348(.I0(un4_v_high_s_2_31),.I1(un4_v_low_s_2_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1348.INIT=32'hACACFF00;
  LUT5 desc1349(.I0(un4_v_high_s_1_31),.I1(un4_v_low_s_1_31),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_36[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1349.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[36:36]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1350(.I0(acs_prob_tdata_8[0:0]),.I1(acs_prob_tdata_9[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1350.INIT=16'h9669;
  LUT2 desc1351(.I0(un4_v_high_s_1_31),.I1(un4_v_low_s_1_31),.O(v_diff_1_axb_1));
defparam desc1351.INIT=4'h9;
  LUT2 desc1352(.I0(un4_v_high_s_2_31),.I1(un4_v_low_s_2_31),.O(v_diff_1_axb_2));
defparam desc1352.INIT=4'h9;
  LUT2 desc1353(.I0(un4_v_high_s_3_31),.I1(un4_v_low_s_3_31),.O(v_diff_1_axb_3));
defparam desc1353.INIT=4'h9;
  LUT2 desc1354(.I0(un4_v_high_s_4_31),.I1(un4_v_low_s_4_31),.O(v_diff_1_axb_4));
defparam desc1354.INIT=4'h9;
  LUT2 desc1355(.I0(un4_v_high_s_5_31),.I1(un4_v_low_s_5_31),.O(v_diff_1_axb_5));
defparam desc1355.INIT=4'h9;
  LUT2 desc1356(.I0(un4_v_high_s_6_31),.I1(un4_v_low_s_6_31),.O(v_diff_1_axb_6));
defparam desc1356.INIT=4'h9;
  LUT2 desc1357(.I0(un4_v_high_s_7_31),.I1(un4_v_low_s_7_31),.O(v_diff_1_axb_7));
defparam desc1357.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_8[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_8[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_8[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_8[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_8[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_8[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_8[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_9[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_9[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_9[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_9[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_9[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_9[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_9[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_9[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1358(.I0(acs_prob_tdata_8[0:0]),.I1(acs_prob_tdata_9[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1728));
defparam desc1358.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_9[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_8[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1359(.I0(un4_v_high_s_8_31),.I1(un4_v_low_s_8_31),.O(v_diff_1_axb_8));
defparam desc1359.INIT=4'h9;
  LUT6 desc1360(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1360.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI48B81(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI48B81.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIMAGB1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIMAGB1));
defparam s_axis_inbranch_tlast_d_RNIMAGB1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_8[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIKPL21_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_31));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_31));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_9[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_31));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_9[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_31));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_9[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_31));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_9[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_31));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_9[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_31));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_9[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_31));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_9[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_9[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_31));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_31));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_8[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_31));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_8[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_31));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_8[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_31));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_8[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_31));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_8[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_31));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_8[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_31));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_8[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_8[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1361(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1362(.DI(un4_v_low_s_7_31),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1363(.DI(un4_v_low_s_6_31),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1364(.DI(un4_v_low_s_5_31),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1365(.DI(un4_v_low_s_4_31),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1366(.DI(un4_v_low_s_3_31),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1367(.DI(un4_v_low_s_2_31),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1368(.DI(un4_v_low_s_1_31),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1369(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1370(.Q(acs_prob_tdata_36[0:0]),.D(N_1728),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMAGB1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1370_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1371(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIKPL21_O6));
defparam desc1371.INIT=16'hF4F0;
  LUT2 desc1372(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1372.INIT=4'h8;
endmodule
module acsZ0_32_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_43,acs_prob_tdata_42,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_21,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1379_p_O_FD,p_desc1380_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1409_p_O_FDRE);
input branch_tlast ;
output [21:21] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_43 ;
input [8:0] acs_prob_tdata_42 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_21 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI2I111_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIAMQB1 ;
wire un4_v_high_s_7_32 ;
wire un4_v_low_s_7_32 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_32 ;
wire un4_v_low_s_8_32 ;
wire un4_v_high_s_6_32 ;
wire un4_v_low_s_6_32 ;
wire un4_v_high_s_5_32 ;
wire un4_v_low_s_5_32 ;
wire un4_v_high_s_4_32 ;
wire un4_v_low_s_4_32 ;
wire un4_v_high_s_3_32 ;
wire un4_v_low_s_3_32 ;
wire un4_v_high_s_2_32 ;
wire un4_v_low_s_2_32 ;
wire un4_v_high_s_1_32 ;
wire un4_v_low_s_1_32 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1708 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1379_p_O_FD ;
input p_desc1380_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1409_p_O_FDRE ;
// instances
  FDR desc1373(.Q(acs_prob_tdata_21[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  FDR desc1374(.Q(acs_prob_tdata_21[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  FDR desc1375(.Q(acs_prob_tdata_21[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  FDR desc1376(.Q(acs_prob_tdata_21[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  FDR desc1377(.Q(acs_prob_tdata_21[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  FDR desc1378(.Q(acs_prob_tdata_21[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1));
  p_O_FD desc1379(.Q(acs_prob_tdata_21[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1379_p_O_FD));
  p_O_FD desc1380(.Q(acs_prob_tdata_21[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1380_p_O_FD));
  LUT6 desc1381(.I0(un4_v_high_s_7_32),.I1(un4_v_low_s_7_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAMQB1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1381.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1382(.I0(un4_v_high_s_8_32),.I1(un4_v_low_s_8_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAMQB1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1382.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1383(.I0(un4_v_high_s_6_32),.I1(un4_v_low_s_6_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1383.INIT=32'hACACFF00;
  LUT5 desc1384(.I0(un4_v_high_s_5_32),.I1(un4_v_low_s_5_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1384.INIT=32'hACACFF00;
  LUT5 desc1385(.I0(un4_v_high_s_4_32),.I1(un4_v_low_s_4_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1385.INIT=32'hACACFF00;
  LUT5 desc1386(.I0(un4_v_high_s_3_32),.I1(un4_v_low_s_3_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1386.INIT=32'hACACFF00;
  LUT5 desc1387(.I0(un4_v_high_s_2_32),.I1(un4_v_low_s_2_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1387.INIT=32'hACACFF00;
  LUT5 desc1388(.I0(un4_v_high_s_1_32),.I1(un4_v_low_s_1_32),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_21[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1388.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[21:21]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1389(.I0(acs_prob_tdata_42[0:0]),.I1(acs_prob_tdata_43[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1389.INIT=16'h9669;
  LUT2 desc1390(.I0(un4_v_high_s_1_32),.I1(un4_v_low_s_1_32),.O(v_diff_1_axb_1));
defparam desc1390.INIT=4'h9;
  LUT2 desc1391(.I0(un4_v_high_s_2_32),.I1(un4_v_low_s_2_32),.O(v_diff_1_axb_2));
defparam desc1391.INIT=4'h9;
  LUT2 desc1392(.I0(un4_v_high_s_3_32),.I1(un4_v_low_s_3_32),.O(v_diff_1_axb_3));
defparam desc1392.INIT=4'h9;
  LUT2 desc1393(.I0(un4_v_high_s_4_32),.I1(un4_v_low_s_4_32),.O(v_diff_1_axb_4));
defparam desc1393.INIT=4'h9;
  LUT2 desc1394(.I0(un4_v_high_s_5_32),.I1(un4_v_low_s_5_32),.O(v_diff_1_axb_5));
defparam desc1394.INIT=4'h9;
  LUT2 desc1395(.I0(un4_v_high_s_6_32),.I1(un4_v_low_s_6_32),.O(v_diff_1_axb_6));
defparam desc1395.INIT=4'h9;
  LUT2 desc1396(.I0(un4_v_high_s_7_32),.I1(un4_v_low_s_7_32),.O(v_diff_1_axb_7));
defparam desc1396.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_42[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_42[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_42[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_42[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_42[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_42[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_42[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_43[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_43[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_43[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_43[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_43[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_43[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_43[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_43[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1397(.I0(acs_prob_tdata_42[0:0]),.I1(acs_prob_tdata_43[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1708));
defparam desc1397.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_43[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_42[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1398(.I0(un4_v_high_s_8_32),.I1(un4_v_low_s_8_32),.O(v_diff_1_axb_8));
defparam desc1398.INIT=4'h9;
  LUT6 desc1399(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1399.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIOJL81(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIOJL81.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIAMQB1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIAMQB1));
defparam s_axis_inbranch_tlast_d_RNIAMQB1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_42[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI2I111_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_32));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_32));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_43[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_32));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_43[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_32));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_43[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_32));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_43[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_32));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_43[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_32));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_43[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_32));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_43[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_43[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_32));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_32));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_42[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_32));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_42[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_32));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_42[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_32));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_42[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_32));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_42[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_32));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_42[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_32));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_42[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_42[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1400(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1401(.DI(un4_v_low_s_7_32),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1402(.DI(un4_v_low_s_6_32),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1403(.DI(un4_v_low_s_5_32),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1404(.DI(un4_v_low_s_4_32),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1405(.DI(un4_v_low_s_3_32),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1406(.DI(un4_v_low_s_2_32),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1407(.DI(un4_v_low_s_1_32),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1408(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1409(.Q(acs_prob_tdata_21[0:0]),.D(N_1708),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAMQB1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1409_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1410(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI2I111_O6));
defparam desc1410.INIT=16'hF4F0;
  LUT2 desc1411(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1411.INIT=4'h8;
endmodule
module acsZ0_33_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_43,acs_prob_tdata_42,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_53,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,N_1756_1,aresetn,p_desc1418_p_O_FD,p_desc1419_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1448_p_O_FDRE);
input branch_tlast ;
output [53:53] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_43 ;
input [8:0] acs_prob_tdata_42 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_53 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIH92V_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIKBJV ;
wire un4_v_high_s_7_33 ;
wire un4_v_low_s_7_33 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_33 ;
wire un4_v_low_s_8_33 ;
wire un4_v_high_s_6_33 ;
wire un4_v_low_s_6_33 ;
wire un4_v_high_s_5_33 ;
wire un4_v_low_s_5_33 ;
wire un4_v_high_s_4_33 ;
wire un4_v_low_s_4_33 ;
wire un4_v_high_s_3_33 ;
wire un4_v_low_s_3_33 ;
wire un4_v_high_s_2_33 ;
wire un4_v_low_s_2_33 ;
wire un4_v_high_s_1_33 ;
wire un4_v_low_s_1_33 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1688 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1418_p_O_FD ;
input p_desc1419_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1448_p_O_FDRE ;
// instances
  FDR desc1412(.Q(acs_prob_tdata_53[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  FDR desc1413(.Q(acs_prob_tdata_53[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  FDR desc1414(.Q(acs_prob_tdata_53[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  FDR desc1415(.Q(acs_prob_tdata_53[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  FDR desc1416(.Q(acs_prob_tdata_53[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  FDR desc1417(.Q(acs_prob_tdata_53[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV));
  p_O_FD desc1418(.Q(acs_prob_tdata_53[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1418_p_O_FD));
  p_O_FD desc1419(.Q(acs_prob_tdata_53[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1419_p_O_FD));
  LUT6 desc1420(.I0(un4_v_high_s_7_33),.I1(un4_v_low_s_7_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKBJV),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1420.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1421(.I0(un4_v_high_s_8_33),.I1(un4_v_low_s_8_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKBJV),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1421.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1422(.I0(un4_v_high_s_6_33),.I1(un4_v_low_s_6_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1422.INIT=32'hACACFF00;
  LUT5 desc1423(.I0(un4_v_high_s_5_33),.I1(un4_v_low_s_5_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1423.INIT=32'hACACFF00;
  LUT5 desc1424(.I0(un4_v_high_s_4_33),.I1(un4_v_low_s_4_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1424.INIT=32'hACACFF00;
  LUT5 desc1425(.I0(un4_v_high_s_3_33),.I1(un4_v_low_s_3_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1425.INIT=32'hACACFF00;
  LUT5 desc1426(.I0(un4_v_high_s_2_33),.I1(un4_v_low_s_2_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1426.INIT=32'hACACFF00;
  LUT5 desc1427(.I0(un4_v_high_s_1_33),.I1(un4_v_low_s_1_33),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_53[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1427.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[53:53]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1428(.I0(acs_prob_tdata_42[0:0]),.I1(acs_prob_tdata_43[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1428.INIT=16'h9669;
  LUT2 desc1429(.I0(un4_v_high_s_1_33),.I1(un4_v_low_s_1_33),.O(v_diff_1_axb_1));
defparam desc1429.INIT=4'h9;
  LUT2 desc1430(.I0(un4_v_high_s_2_33),.I1(un4_v_low_s_2_33),.O(v_diff_1_axb_2));
defparam desc1430.INIT=4'h9;
  LUT2 desc1431(.I0(un4_v_high_s_3_33),.I1(un4_v_low_s_3_33),.O(v_diff_1_axb_3));
defparam desc1431.INIT=4'h9;
  LUT2 desc1432(.I0(un4_v_high_s_4_33),.I1(un4_v_low_s_4_33),.O(v_diff_1_axb_4));
defparam desc1432.INIT=4'h9;
  LUT2 desc1433(.I0(un4_v_high_s_5_33),.I1(un4_v_low_s_5_33),.O(v_diff_1_axb_5));
defparam desc1433.INIT=4'h9;
  LUT2 desc1434(.I0(un4_v_high_s_6_33),.I1(un4_v_low_s_6_33),.O(v_diff_1_axb_6));
defparam desc1434.INIT=4'h9;
  LUT2 desc1435(.I0(un4_v_high_s_7_33),.I1(un4_v_low_s_7_33),.O(v_diff_1_axb_7));
defparam desc1435.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_42[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_42[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_42[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_42[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_42[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_42[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_42[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_43[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_43[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_43[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_43[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_43[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_43[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_43[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_43[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1436(.I0(acs_prob_tdata_42[0:0]),.I1(acs_prob_tdata_43[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1688));
defparam desc1436.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_43[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_42[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1437(.I0(un4_v_high_s_8_33),.I1(un4_v_low_s_8_33),.O(v_diff_1_axb_8));
defparam desc1437.INIT=4'h9;
  LUT6 desc1438(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1438.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI29ES(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI29ES.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIKBJV_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIKBJV));
defparam s_axis_inbranch_tlast_d_RNIKBJV_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_42[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIH92V_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_33));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_33));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_43[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_33));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_43[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_33));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_43[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_33));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_43[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_33));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_43[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_33));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_43[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_33));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_43[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_43[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_33));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_33));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_42[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_33));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_42[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_33));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_42[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_33));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_42[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_33));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_42[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_33));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_42[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_33));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_42[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_42[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1439(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1440(.DI(un4_v_low_s_7_33),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1441(.DI(un4_v_low_s_6_33),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1442(.DI(un4_v_low_s_5_33),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1443(.DI(un4_v_low_s_4_33),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1444(.DI(un4_v_low_s_3_33),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1445(.DI(un4_v_low_s_2_33),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1446(.DI(un4_v_low_s_1_33),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1447(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1448(.Q(acs_prob_tdata_53[0:0]),.D(N_1688),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKBJV),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1448_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1449(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIH92V_O6));
defparam desc1449.INIT=16'hF4F0;
  LUT2 desc1450(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1450.INIT=4'h8;
endmodule
module acsZ0_34_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_23,acs_prob_tdata_22,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_11,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1457_p_O_FD,p_desc1458_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1487_p_O_FDRE);
input branch_tlast ;
output [11:11] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_23 ;
input [8:0] acs_prob_tdata_22 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_11 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIVOBU_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI8HK61 ;
wire un4_v_high_s_7_34 ;
wire un4_v_low_s_7_34 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_34 ;
wire un4_v_low_s_8_34 ;
wire un4_v_high_s_6_34 ;
wire un4_v_low_s_6_34 ;
wire un4_v_high_s_5_34 ;
wire un4_v_low_s_5_34 ;
wire un4_v_high_s_4_34 ;
wire un4_v_low_s_4_34 ;
wire un4_v_high_s_3_34 ;
wire un4_v_low_s_3_34 ;
wire un4_v_high_s_2_34 ;
wire un4_v_low_s_2_34 ;
wire un4_v_high_s_1_34 ;
wire un4_v_low_s_1_34 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1668 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1457_p_O_FD ;
input p_desc1458_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1487_p_O_FDRE ;
// instances
  FDR desc1451(.Q(acs_prob_tdata_11[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  FDR desc1452(.Q(acs_prob_tdata_11[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  FDR desc1453(.Q(acs_prob_tdata_11[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  FDR desc1454(.Q(acs_prob_tdata_11[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  FDR desc1455(.Q(acs_prob_tdata_11[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  FDR desc1456(.Q(acs_prob_tdata_11[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61));
  p_O_FD desc1457(.Q(acs_prob_tdata_11[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1457_p_O_FD));
  p_O_FD desc1458(.Q(acs_prob_tdata_11[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1458_p_O_FD));
  LUT6 desc1459(.I0(un4_v_high_s_7_34),.I1(un4_v_low_s_7_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI8HK61),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1459.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1460(.I0(un4_v_high_s_8_34),.I1(un4_v_low_s_8_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI8HK61),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1460.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1461(.I0(un4_v_high_s_6_34),.I1(un4_v_low_s_6_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1461.INIT=32'hACACFF00;
  LUT5 desc1462(.I0(un4_v_high_s_5_34),.I1(un4_v_low_s_5_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1462.INIT=32'hACACFF00;
  LUT5 desc1463(.I0(un4_v_high_s_4_34),.I1(un4_v_low_s_4_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1463.INIT=32'hACACFF00;
  LUT5 desc1464(.I0(un4_v_high_s_3_34),.I1(un4_v_low_s_3_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1464.INIT=32'hACACFF00;
  LUT5 desc1465(.I0(un4_v_high_s_2_34),.I1(un4_v_low_s_2_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1465.INIT=32'hACACFF00;
  LUT5 desc1466(.I0(un4_v_high_s_1_34),.I1(un4_v_low_s_1_34),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_11[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1466.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[11:11]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_22[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_22[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_22[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_22[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_22[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_22[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_22[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_23[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_23[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_23[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_23[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_23[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_23[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_23[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_23[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1467(.I0(acs_prob_tdata_22[0:0]),.I1(acs_prob_tdata_23[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1467.INIT=16'h9669;
  LUT2 desc1468(.I0(un4_v_high_s_1_34),.I1(un4_v_low_s_1_34),.O(v_diff_1_axb_1));
defparam desc1468.INIT=4'h9;
  LUT2 desc1469(.I0(un4_v_high_s_2_34),.I1(un4_v_low_s_2_34),.O(v_diff_1_axb_2));
defparam desc1469.INIT=4'h9;
  LUT2 desc1470(.I0(un4_v_high_s_3_34),.I1(un4_v_low_s_3_34),.O(v_diff_1_axb_3));
defparam desc1470.INIT=4'h9;
  LUT2 desc1471(.I0(un4_v_high_s_4_34),.I1(un4_v_low_s_4_34),.O(v_diff_1_axb_4));
defparam desc1471.INIT=4'h9;
  LUT2 desc1472(.I0(un4_v_high_s_5_34),.I1(un4_v_low_s_5_34),.O(v_diff_1_axb_5));
defparam desc1472.INIT=4'h9;
  LUT2 desc1473(.I0(un4_v_high_s_6_34),.I1(un4_v_low_s_6_34),.O(v_diff_1_axb_6));
defparam desc1473.INIT=4'h9;
  LUT2 desc1474(.I0(un4_v_high_s_7_34),.I1(un4_v_low_s_7_34),.O(v_diff_1_axb_7));
defparam desc1474.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1475(.I0(acs_prob_tdata_22[0:0]),.I1(acs_prob_tdata_23[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1668));
defparam desc1475.INIT=32'h3C3C55AA;
  LUT2 desc1476(.I0(un4_v_high_s_8_34),.I1(un4_v_low_s_8_34),.O(v_diff_1_axb_8));
defparam desc1476.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_23[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_22[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1477(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1477.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIMEF31(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIMEF31.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI8HK61_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI8HK61));
defparam s_axis_inbranch_tlast_d_RNI8HK61_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_22[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIVOBU_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1478(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1479(.DI(un4_v_low_s_7_34),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1480(.DI(un4_v_low_s_6_34),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1481(.DI(un4_v_low_s_5_34),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1482(.DI(un4_v_low_s_4_34),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1483(.DI(un4_v_low_s_3_34),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1484(.DI(un4_v_low_s_2_34),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1485(.DI(un4_v_low_s_1_34),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1486(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_34));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_34));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_23[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_34));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_23[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_34));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_23[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_34));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_23[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_34));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_23[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_34));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_23[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_34));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_23[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_23[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_34));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_34));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_22[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_34));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_22[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_34));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_22[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_34));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_22[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_34));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_22[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_34));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_22[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_34));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_22[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_22[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1487(.Q(acs_prob_tdata_11[0:0]),.D(N_1668),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8HK61),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1487_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1488(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIVOBU_O6));
defparam desc1488.INIT=16'hF4F0;
  LUT2 desc1489(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1489.INIT=4'h8;
endmodule
module acsZ0_35_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_47,acs_prob_tdata_46,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_23,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_3_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1496_p_O_FD,p_desc1497_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1526_p_O_FDRE);
input branch_tlast ;
output [23:23] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_47 ;
input [8:0] acs_prob_tdata_46 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_23 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_3_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_3_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI8U071_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIES0G1 ;
wire un4_v_high_s_7_35 ;
wire un4_v_low_s_7_35 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_35 ;
wire un4_v_low_s_8_35 ;
wire un4_v_high_s_6_35 ;
wire un4_v_low_s_6_35 ;
wire un4_v_high_s_5_35 ;
wire un4_v_low_s_5_35 ;
wire un4_v_high_s_4_35 ;
wire un4_v_low_s_4_35 ;
wire un4_v_high_s_3_35 ;
wire un4_v_low_s_3_35 ;
wire un4_v_high_s_2_35 ;
wire un4_v_low_s_2_35 ;
wire un4_v_high_s_1_35 ;
wire un4_v_low_s_1_35 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1648 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1496_p_O_FD ;
input p_desc1497_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1526_p_O_FDRE ;
// instances
  FDR desc1490(.Q(acs_prob_tdata_23[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  FDR desc1491(.Q(acs_prob_tdata_23[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  FDR desc1492(.Q(acs_prob_tdata_23[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  FDR desc1493(.Q(acs_prob_tdata_23[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  FDR desc1494(.Q(acs_prob_tdata_23[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  FDR desc1495(.Q(acs_prob_tdata_23[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1));
  p_O_FD desc1496(.Q(acs_prob_tdata_23[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1496_p_O_FD));
  p_O_FD desc1497(.Q(acs_prob_tdata_23[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1497_p_O_FD));
  LUT6 desc1498(.I0(un4_v_high_s_7_35),.I1(un4_v_low_s_7_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIES0G1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1498.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1499(.I0(un4_v_high_s_8_35),.I1(un4_v_low_s_8_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIES0G1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1499.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1500(.I0(un4_v_high_s_6_35),.I1(un4_v_low_s_6_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1500.INIT=32'hACACFF00;
  LUT5 desc1501(.I0(un4_v_high_s_5_35),.I1(un4_v_low_s_5_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1501.INIT=32'hACACFF00;
  LUT5 desc1502(.I0(un4_v_high_s_4_35),.I1(un4_v_low_s_4_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1502.INIT=32'hACACFF00;
  LUT5 desc1503(.I0(un4_v_high_s_3_35),.I1(un4_v_low_s_3_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1503.INIT=32'hACACFF00;
  LUT5 desc1504(.I0(un4_v_high_s_2_35),.I1(un4_v_low_s_2_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1504.INIT=32'hACACFF00;
  LUT5 desc1505(.I0(un4_v_high_s_1_35),.I1(un4_v_low_s_1_35),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_23[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1505.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[23:23]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_46[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_46[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_46[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_46[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_46[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_46[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_46[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_47[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_47[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_47[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_47[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_47[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_47[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_47[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_47[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1506(.I0(acs_prob_tdata_46[0:0]),.I1(acs_prob_tdata_47[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1506.INIT=16'h9669;
  LUT2 desc1507(.I0(un4_v_high_s_1_35),.I1(un4_v_low_s_1_35),.O(v_diff_1_axb_1));
defparam desc1507.INIT=4'h9;
  LUT2 desc1508(.I0(un4_v_high_s_2_35),.I1(un4_v_low_s_2_35),.O(v_diff_1_axb_2));
defparam desc1508.INIT=4'h9;
  LUT2 desc1509(.I0(un4_v_high_s_3_35),.I1(un4_v_low_s_3_35),.O(v_diff_1_axb_3));
defparam desc1509.INIT=4'h9;
  LUT2 desc1510(.I0(un4_v_high_s_4_35),.I1(un4_v_low_s_4_35),.O(v_diff_1_axb_4));
defparam desc1510.INIT=4'h9;
  LUT2 desc1511(.I0(un4_v_high_s_5_35),.I1(un4_v_low_s_5_35),.O(v_diff_1_axb_5));
defparam desc1511.INIT=4'h9;
  LUT2 desc1512(.I0(un4_v_high_s_6_35),.I1(un4_v_low_s_6_35),.O(v_diff_1_axb_6));
defparam desc1512.INIT=4'h9;
  LUT2 desc1513(.I0(un4_v_high_s_7_35),.I1(un4_v_low_s_7_35),.O(v_diff_1_axb_7));
defparam desc1513.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1514(.I0(acs_prob_tdata_46[0:0]),.I1(acs_prob_tdata_47[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1648));
defparam desc1514.INIT=32'h33CC5A5A;
  LUT2 desc1515(.I0(un4_v_high_s_8_35),.I1(un4_v_low_s_8_35),.O(v_diff_1_axb_8));
defparam desc1515.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_47[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_46[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1516(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1516.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNISPRC1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNISPRC1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIES0G1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIES0G1));
defparam s_axis_inbranch_tlast_d_RNIES0G1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_46[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI8U071_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1517(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1518(.DI(un4_v_low_s_7_35),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1519(.DI(un4_v_low_s_6_35),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1520(.DI(un4_v_low_s_5_35),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1521(.DI(un4_v_low_s_4_35),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1522(.DI(un4_v_low_s_3_35),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1523(.DI(un4_v_low_s_2_35),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1524(.DI(un4_v_low_s_1_35),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1525(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_35));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_35));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_47[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_35));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_47[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_35));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_47[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_35));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_47[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_35));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_47[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_35));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_47[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_35));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_47[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_47[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_35));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_35));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_46[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_35));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_46[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_35));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_46[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_35));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_46[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_35));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_46[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_35));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_46[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_35));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_46[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_46[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1526(.Q(acs_prob_tdata_23[0:0]),.D(N_1648),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIES0G1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1526_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1527(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI8U071_O6));
defparam desc1527.INIT=16'hF4F0;
  LUT2 desc1528(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1528.INIT=4'h8;
endmodule
module acsZ0_36_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_16,acs_prob_tdata_17,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_8,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1535_p_O_FD,p_desc1536_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1565_p_O_FDRE);
input branch_tlast ;
output [8:8] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_16 ;
input [8:0] acs_prob_tdata_17 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_8 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI1CD61_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIKI461 ;
wire un4_v_high_s_7_36 ;
wire un4_v_low_s_7_36 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_36 ;
wire un4_v_low_s_8_36 ;
wire un4_v_high_s_6_36 ;
wire un4_v_low_s_6_36 ;
wire un4_v_high_s_5_36 ;
wire un4_v_low_s_5_36 ;
wire un4_v_high_s_4_36 ;
wire un4_v_low_s_4_36 ;
wire un4_v_high_s_3_36 ;
wire un4_v_low_s_3_36 ;
wire un4_v_high_s_2_36 ;
wire un4_v_low_s_2_36 ;
wire un4_v_high_s_1_36 ;
wire un4_v_low_s_1_36 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire N_1628 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire GND ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire N_1 ;
input p_desc1535_p_O_FD ;
input p_desc1536_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1565_p_O_FDRE ;
// instances
  FDR desc1529(.Q(acs_prob_tdata_8[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  FDR desc1530(.Q(acs_prob_tdata_8[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  FDR desc1531(.Q(acs_prob_tdata_8[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  FDR desc1532(.Q(acs_prob_tdata_8[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  FDR desc1533(.Q(acs_prob_tdata_8[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  FDR desc1534(.Q(acs_prob_tdata_8[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461));
  p_O_FD desc1535(.Q(acs_prob_tdata_8[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1535_p_O_FD));
  p_O_FD desc1536(.Q(acs_prob_tdata_8[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1536_p_O_FD));
  LUT6 desc1537(.I0(un4_v_high_s_7_36),.I1(un4_v_low_s_7_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKI461),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1537.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1538(.I0(un4_v_high_s_8_36),.I1(un4_v_low_s_8_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIKI461),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1538.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1539(.I0(un4_v_high_s_6_36),.I1(un4_v_low_s_6_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1539.INIT=32'hACACFF00;
  LUT5 desc1540(.I0(un4_v_high_s_5_36),.I1(un4_v_low_s_5_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1540.INIT=32'hACACFF00;
  LUT5 desc1541(.I0(un4_v_high_s_4_36),.I1(un4_v_low_s_4_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1541.INIT=32'hACACFF00;
  LUT5 desc1542(.I0(un4_v_high_s_3_36),.I1(un4_v_low_s_3_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1542.INIT=32'hACACFF00;
  LUT5 desc1543(.I0(un4_v_high_s_2_36),.I1(un4_v_low_s_2_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1543.INIT=32'hACACFF00;
  LUT5 desc1544(.I0(un4_v_high_s_1_36),.I1(un4_v_low_s_1_36),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_8[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1544.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[8:8]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_17[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_17[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_17[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_17[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_17[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_17[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_17[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_17[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1545(.I0(acs_prob_tdata_16[0:0]),.I1(acs_prob_tdata_17[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1545.INIT=16'h9669;
  LUT2 desc1546(.I0(un4_v_high_s_1_36),.I1(un4_v_low_s_1_36),.O(v_diff_1_axb_1));
defparam desc1546.INIT=4'h9;
  LUT2 desc1547(.I0(un4_v_high_s_2_36),.I1(un4_v_low_s_2_36),.O(v_diff_1_axb_2));
defparam desc1547.INIT=4'h9;
  LUT2 desc1548(.I0(un4_v_high_s_3_36),.I1(un4_v_low_s_3_36),.O(v_diff_1_axb_3));
defparam desc1548.INIT=4'h9;
  LUT2 desc1549(.I0(un4_v_high_s_4_36),.I1(un4_v_low_s_4_36),.O(v_diff_1_axb_4));
defparam desc1549.INIT=4'h9;
  LUT2 desc1550(.I0(un4_v_high_s_5_36),.I1(un4_v_low_s_5_36),.O(v_diff_1_axb_5));
defparam desc1550.INIT=4'h9;
  LUT2 desc1551(.I0(un4_v_high_s_6_36),.I1(un4_v_low_s_6_36),.O(v_diff_1_axb_6));
defparam desc1551.INIT=4'h9;
  LUT2 desc1552(.I0(un4_v_high_s_7_36),.I1(un4_v_low_s_7_36),.O(v_diff_1_axb_7));
defparam desc1552.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_16[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_16[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_16[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_16[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_16[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_16[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_16[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1553(.I0(acs_prob_tdata_16[0:0]),.I1(acs_prob_tdata_17[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1628));
defparam desc1553.INIT=32'h3C3C55AA;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_16[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1554(.I0(un4_v_high_s_8_36),.I1(un4_v_low_s_8_36),.O(v_diff_1_axb_8));
defparam desc1554.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_17[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT6 desc1555(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1555.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI2GV21(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI2GV21.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIKI461_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIKI461));
defparam s_axis_inbranch_tlast_d_RNIKI461_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_16[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI1CD61_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_36));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_36));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_16[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_36));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_16[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_36));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_16[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_36));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_16[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_36));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_16[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_36));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_16[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_36));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_16[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_16[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1556(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1557(.DI(un4_v_low_s_7_36),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1558(.DI(un4_v_low_s_6_36),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1559(.DI(un4_v_low_s_5_36),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1560(.DI(un4_v_low_s_4_36),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1561(.DI(un4_v_low_s_3_36),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1562(.DI(un4_v_low_s_2_36),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1563(.DI(un4_v_low_s_1_36),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1564(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_36));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_36));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_17[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_36));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_17[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_36));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_17[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_36));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_17[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_36));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_17[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_36));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_17[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_36));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_17[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_17[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  p_O_FDRE desc1565(.Q(acs_prob_tdata_8[0:0]),.D(N_1628),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIKI461),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1565_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1566(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI1CD61_O6));
defparam desc1566.INIT=16'hF4F0;
  LUT2 desc1567(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1567.INIT=4'h8;
endmodule
module acsZ0_37_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_17,acs_prob_tdata_16,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_40,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc1574_p_O_FD,p_desc1575_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1604_p_O_FDRE);
input branch_tlast ;
output [40:40] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_17 ;
input [8:0] acs_prob_tdata_16 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_40 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI5ED31_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNICT341 ;
wire un4_v_high_s_7_37 ;
wire un4_v_low_s_7_37 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_37 ;
wire un4_v_low_s_8_37 ;
wire un4_v_high_s_6_37 ;
wire un4_v_low_s_6_37 ;
wire un4_v_high_s_5_37 ;
wire un4_v_low_s_5_37 ;
wire un4_v_high_s_4_37 ;
wire un4_v_low_s_4_37 ;
wire un4_v_high_s_3_37 ;
wire un4_v_low_s_3_37 ;
wire un4_v_high_s_2_37 ;
wire un4_v_low_s_2_37 ;
wire un4_v_high_s_1_37 ;
wire un4_v_low_s_1_37 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1608 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1574_p_O_FD ;
input p_desc1575_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1604_p_O_FDRE ;
// instances
  FDR desc1568(.Q(acs_prob_tdata_40[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  FDR desc1569(.Q(acs_prob_tdata_40[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  FDR desc1570(.Q(acs_prob_tdata_40[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  FDR desc1571(.Q(acs_prob_tdata_40[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  FDR desc1572(.Q(acs_prob_tdata_40[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  FDR desc1573(.Q(acs_prob_tdata_40[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341));
  p_O_FD desc1574(.Q(acs_prob_tdata_40[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1574_p_O_FD));
  p_O_FD desc1575(.Q(acs_prob_tdata_40[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1575_p_O_FD));
  LUT6 desc1576(.I0(un4_v_high_s_7_37),.I1(un4_v_low_s_7_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICT341),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1576.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1577(.I0(un4_v_high_s_8_37),.I1(un4_v_low_s_8_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICT341),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1577.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1578(.I0(un4_v_high_s_6_37),.I1(un4_v_low_s_6_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1578.INIT=32'hACACFF00;
  LUT5 desc1579(.I0(un4_v_high_s_5_37),.I1(un4_v_low_s_5_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1579.INIT=32'hACACFF00;
  LUT5 desc1580(.I0(un4_v_high_s_4_37),.I1(un4_v_low_s_4_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1580.INIT=32'hACACFF00;
  LUT5 desc1581(.I0(un4_v_high_s_3_37),.I1(un4_v_low_s_3_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1581.INIT=32'hACACFF00;
  LUT5 desc1582(.I0(un4_v_high_s_2_37),.I1(un4_v_low_s_2_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1582.INIT=32'hACACFF00;
  LUT5 desc1583(.I0(un4_v_high_s_1_37),.I1(un4_v_low_s_1_37),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_40[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1583.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[40:40]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1584(.I0(acs_prob_tdata_16[0:0]),.I1(acs_prob_tdata_17[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1584.INIT=16'h9669;
  LUT2 desc1585(.I0(un4_v_high_s_1_37),.I1(un4_v_low_s_1_37),.O(v_diff_1_axb_1));
defparam desc1585.INIT=4'h9;
  LUT2 desc1586(.I0(un4_v_high_s_2_37),.I1(un4_v_low_s_2_37),.O(v_diff_1_axb_2));
defparam desc1586.INIT=4'h9;
  LUT2 desc1587(.I0(un4_v_high_s_3_37),.I1(un4_v_low_s_3_37),.O(v_diff_1_axb_3));
defparam desc1587.INIT=4'h9;
  LUT2 desc1588(.I0(un4_v_high_s_4_37),.I1(un4_v_low_s_4_37),.O(v_diff_1_axb_4));
defparam desc1588.INIT=4'h9;
  LUT2 desc1589(.I0(un4_v_high_s_5_37),.I1(un4_v_low_s_5_37),.O(v_diff_1_axb_5));
defparam desc1589.INIT=4'h9;
  LUT2 desc1590(.I0(un4_v_high_s_6_37),.I1(un4_v_low_s_6_37),.O(v_diff_1_axb_6));
defparam desc1590.INIT=4'h9;
  LUT2 desc1591(.I0(un4_v_high_s_7_37),.I1(un4_v_low_s_7_37),.O(v_diff_1_axb_7));
defparam desc1591.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_16[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_16[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_16[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_16[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_16[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_16[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_16[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_17[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_17[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_17[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_17[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_17[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_17[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_17[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_17[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1592(.I0(acs_prob_tdata_16[0:0]),.I1(acs_prob_tdata_17[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1608));
defparam desc1592.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_17[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_16[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1593(.I0(un4_v_high_s_8_37),.I1(un4_v_low_s_8_37),.O(v_diff_1_axb_8));
defparam desc1593.INIT=4'h9;
  LUT6 desc1594(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1594.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIQQU01(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQQU01.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNICT341_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNICT341));
defparam s_axis_inbranch_tlast_d_RNICT341_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_16[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI5ED31_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_37));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_37));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_17[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_37));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_17[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_37));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_17[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_37));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_17[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_37));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_17[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_37));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_17[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_37));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_17[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_17[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_37));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_37));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_16[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_37));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_16[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_37));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_16[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_37));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_16[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_37));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_16[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_37));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_16[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_37));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_16[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_16[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1595(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1596(.DI(un4_v_low_s_7_37),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1597(.DI(un4_v_low_s_6_37),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1598(.DI(un4_v_low_s_5_37),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1599(.DI(un4_v_low_s_4_37),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1600(.DI(un4_v_low_s_3_37),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1601(.DI(un4_v_low_s_2_37),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1602(.DI(un4_v_low_s_1_37),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1603(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1604(.Q(acs_prob_tdata_40[0:0]),.D(N_1608),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICT341),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1604_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1605(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI5ED31_O6));
defparam desc1605.INIT=16'hF4F0;
  LUT2 desc1606(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1606.INIT=4'h8;
endmodule
module acsZ0_38_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_35,acs_prob_tdata_34,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_17,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1613_p_O_FD,p_desc1614_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1643_p_O_FDRE);
input branch_tlast ;
output [17:17] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_35 ;
input [8:0] acs_prob_tdata_34 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_17 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIHT901_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIK3731 ;
wire un4_v_high_s_7_38 ;
wire un4_v_low_s_7_38 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_38 ;
wire un4_v_low_s_8_38 ;
wire un4_v_high_s_6_38 ;
wire un4_v_low_s_6_38 ;
wire un4_v_high_s_5_38 ;
wire un4_v_low_s_5_38 ;
wire un4_v_high_s_4_38 ;
wire un4_v_low_s_4_38 ;
wire un4_v_high_s_3_38 ;
wire un4_v_low_s_3_38 ;
wire un4_v_high_s_2_38 ;
wire un4_v_low_s_2_38 ;
wire un4_v_high_s_1_38 ;
wire un4_v_low_s_1_38 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1588 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1613_p_O_FD ;
input p_desc1614_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1643_p_O_FDRE ;
// instances
  FDR desc1607(.Q(acs_prob_tdata_17[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  FDR desc1608(.Q(acs_prob_tdata_17[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  FDR desc1609(.Q(acs_prob_tdata_17[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  FDR desc1610(.Q(acs_prob_tdata_17[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  FDR desc1611(.Q(acs_prob_tdata_17[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  FDR desc1612(.Q(acs_prob_tdata_17[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731));
  p_O_FD desc1613(.Q(acs_prob_tdata_17[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1613_p_O_FD));
  p_O_FD desc1614(.Q(acs_prob_tdata_17[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1614_p_O_FD));
  LUT6 desc1615(.I0(un4_v_high_s_7_38),.I1(un4_v_low_s_7_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK3731),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1615.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1616(.I0(un4_v_high_s_8_38),.I1(un4_v_low_s_8_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK3731),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1616.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1617(.I0(un4_v_high_s_6_38),.I1(un4_v_low_s_6_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1617.INIT=32'hACACFF00;
  LUT5 desc1618(.I0(un4_v_high_s_5_38),.I1(un4_v_low_s_5_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1618.INIT=32'hACACFF00;
  LUT5 desc1619(.I0(un4_v_high_s_4_38),.I1(un4_v_low_s_4_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1619.INIT=32'hACACFF00;
  LUT5 desc1620(.I0(un4_v_high_s_3_38),.I1(un4_v_low_s_3_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1620.INIT=32'hACACFF00;
  LUT5 desc1621(.I0(un4_v_high_s_2_38),.I1(un4_v_low_s_2_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1621.INIT=32'hACACFF00;
  LUT5 desc1622(.I0(un4_v_high_s_1_38),.I1(un4_v_low_s_1_38),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_17[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1622.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[17:17]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1623(.I0(acs_prob_tdata_34[0:0]),.I1(acs_prob_tdata_35[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1623.INIT=16'h9669;
  LUT2 desc1624(.I0(un4_v_high_s_1_38),.I1(un4_v_low_s_1_38),.O(v_diff_1_axb_1));
defparam desc1624.INIT=4'h9;
  LUT2 desc1625(.I0(un4_v_high_s_2_38),.I1(un4_v_low_s_2_38),.O(v_diff_1_axb_2));
defparam desc1625.INIT=4'h9;
  LUT2 desc1626(.I0(un4_v_high_s_3_38),.I1(un4_v_low_s_3_38),.O(v_diff_1_axb_3));
defparam desc1626.INIT=4'h9;
  LUT2 desc1627(.I0(un4_v_high_s_4_38),.I1(un4_v_low_s_4_38),.O(v_diff_1_axb_4));
defparam desc1627.INIT=4'h9;
  LUT2 desc1628(.I0(un4_v_high_s_5_38),.I1(un4_v_low_s_5_38),.O(v_diff_1_axb_5));
defparam desc1628.INIT=4'h9;
  LUT2 desc1629(.I0(un4_v_high_s_6_38),.I1(un4_v_low_s_6_38),.O(v_diff_1_axb_6));
defparam desc1629.INIT=4'h9;
  LUT2 desc1630(.I0(un4_v_high_s_7_38),.I1(un4_v_low_s_7_38),.O(v_diff_1_axb_7));
defparam desc1630.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_34[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_34[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_34[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_34[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_34[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_34[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_34[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_35[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_35[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_35[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_35[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_35[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_35[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_35[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_35[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1631(.I0(acs_prob_tdata_34[0:0]),.I1(acs_prob_tdata_35[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1588));
defparam desc1631.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_35[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_34[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1632(.I0(un4_v_high_s_8_38),.I1(un4_v_low_s_8_38),.O(v_diff_1_axb_8));
defparam desc1632.INIT=4'h9;
  LUT6 desc1633(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1633.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI21201(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI21201.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIK3731_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIK3731));
defparam s_axis_inbranch_tlast_d_RNIK3731_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_34[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIHT901_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_38));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_38));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_35[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_38));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_35[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_38));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_35[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_38));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_35[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_38));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_35[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_38));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_35[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_38));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_35[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_35[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_38));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_38));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_34[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_38));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_34[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_38));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_34[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_38));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_34[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_38));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_34[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_38));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_34[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_38));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_34[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_34[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1634(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1635(.DI(un4_v_low_s_7_38),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1636(.DI(un4_v_low_s_6_38),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1637(.DI(un4_v_low_s_5_38),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1638(.DI(un4_v_low_s_4_38),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1639(.DI(un4_v_low_s_3_38),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1640(.DI(un4_v_low_s_2_38),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1641(.DI(un4_v_low_s_1_38),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1642(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1643(.Q(acs_prob_tdata_17[0:0]),.D(N_1588),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK3731),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1643_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1644(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIHT901_O6));
defparam desc1644.INIT=16'hF4F0;
  LUT2 desc1645(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1645.INIT=4'h8;
endmodule
module acsZ0_39_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_37,acs_prob_tdata_36,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_50,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,N_1756_1,aresetn,p_desc1652_p_O_FD,p_desc1653_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1682_p_O_FDRE);
input branch_tlast ;
output [50:50] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_37 ;
input [8:0] acs_prob_tdata_36 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_50 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI87361_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIE2A91 ;
wire un4_v_high_s_7_39 ;
wire un4_v_low_s_7_39 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_39 ;
wire un4_v_low_s_8_39 ;
wire un4_v_high_s_6_39 ;
wire un4_v_low_s_6_39 ;
wire un4_v_high_s_5_39 ;
wire un4_v_low_s_5_39 ;
wire un4_v_high_s_4_39 ;
wire un4_v_low_s_4_39 ;
wire un4_v_high_s_3_39 ;
wire un4_v_low_s_3_39 ;
wire un4_v_high_s_2_39 ;
wire un4_v_low_s_2_39 ;
wire un4_v_high_s_1_39 ;
wire un4_v_low_s_1_39 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1568 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1652_p_O_FD ;
input p_desc1653_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1682_p_O_FDRE ;
// instances
  FDR desc1646(.Q(acs_prob_tdata_50[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  FDR desc1647(.Q(acs_prob_tdata_50[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  FDR desc1648(.Q(acs_prob_tdata_50[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  FDR desc1649(.Q(acs_prob_tdata_50[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  FDR desc1650(.Q(acs_prob_tdata_50[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  FDR desc1651(.Q(acs_prob_tdata_50[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91));
  p_O_FD desc1652(.Q(acs_prob_tdata_50[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1652_p_O_FD));
  p_O_FD desc1653(.Q(acs_prob_tdata_50[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1653_p_O_FD));
  LUT6 desc1654(.I0(un4_v_high_s_7_39),.I1(un4_v_low_s_7_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE2A91),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1654.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1655(.I0(un4_v_high_s_8_39),.I1(un4_v_low_s_8_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE2A91),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1655.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1656(.I0(un4_v_high_s_6_39),.I1(un4_v_low_s_6_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1656.INIT=32'hACACFF00;
  LUT5 desc1657(.I0(un4_v_high_s_5_39),.I1(un4_v_low_s_5_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1657.INIT=32'hACACFF00;
  LUT5 desc1658(.I0(un4_v_high_s_4_39),.I1(un4_v_low_s_4_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1658.INIT=32'hACACFF00;
  LUT5 desc1659(.I0(un4_v_high_s_3_39),.I1(un4_v_low_s_3_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1659.INIT=32'hACACFF00;
  LUT5 desc1660(.I0(un4_v_high_s_2_39),.I1(un4_v_low_s_2_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1660.INIT=32'hACACFF00;
  LUT5 desc1661(.I0(un4_v_high_s_1_39),.I1(un4_v_low_s_1_39),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_50[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1661.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[50:50]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1662(.I0(acs_prob_tdata_36[0:0]),.I1(acs_prob_tdata_37[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1662.INIT=16'h9669;
  LUT2 desc1663(.I0(un4_v_high_s_1_39),.I1(un4_v_low_s_1_39),.O(v_diff_1_axb_1));
defparam desc1663.INIT=4'h9;
  LUT2 desc1664(.I0(un4_v_high_s_2_39),.I1(un4_v_low_s_2_39),.O(v_diff_1_axb_2));
defparam desc1664.INIT=4'h9;
  LUT2 desc1665(.I0(un4_v_high_s_3_39),.I1(un4_v_low_s_3_39),.O(v_diff_1_axb_3));
defparam desc1665.INIT=4'h9;
  LUT2 desc1666(.I0(un4_v_high_s_4_39),.I1(un4_v_low_s_4_39),.O(v_diff_1_axb_4));
defparam desc1666.INIT=4'h9;
  LUT2 desc1667(.I0(un4_v_high_s_5_39),.I1(un4_v_low_s_5_39),.O(v_diff_1_axb_5));
defparam desc1667.INIT=4'h9;
  LUT2 desc1668(.I0(un4_v_high_s_6_39),.I1(un4_v_low_s_6_39),.O(v_diff_1_axb_6));
defparam desc1668.INIT=4'h9;
  LUT2 desc1669(.I0(un4_v_high_s_7_39),.I1(un4_v_low_s_7_39),.O(v_diff_1_axb_7));
defparam desc1669.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_36[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_36[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_36[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_36[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_36[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_36[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_36[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_37[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_37[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_37[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_37[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_37[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_37[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_37[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_37[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1670(.I0(acs_prob_tdata_36[0:0]),.I1(acs_prob_tdata_37[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1568));
defparam desc1670.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_37[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_36[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1671(.I0(un4_v_high_s_8_39),.I1(un4_v_low_s_8_39),.O(v_diff_1_axb_8));
defparam desc1671.INIT=4'h9;
  LUT6 desc1672(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1672.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNISV461(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNISV461.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIE2A91_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIE2A91));
defparam s_axis_inbranch_tlast_d_RNIE2A91_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_36[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI87361_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_39));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_39));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_37[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_39));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_37[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_39));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_37[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_39));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_37[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_39));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_37[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_39));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_37[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_39));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_37[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_37[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_39));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_39));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_36[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_39));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_36[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_39));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_36[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_39));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_36[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_39));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_36[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_39));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_36[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_39));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_36[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_36[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1673(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1674(.DI(un4_v_low_s_7_39),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1675(.DI(un4_v_low_s_6_39),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1676(.DI(un4_v_low_s_5_39),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1677(.DI(un4_v_low_s_4_39),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1678(.DI(un4_v_low_s_3_39),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1679(.DI(un4_v_low_s_2_39),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1680(.DI(un4_v_low_s_1_39),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1681(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1682(.Q(acs_prob_tdata_50[0:0]),.D(N_1568),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE2A91),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1682_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1683(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI87361_O6));
defparam desc1683.INIT=16'hF4F0;
  LUT2 desc1684(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1684.INIT=4'h8;
endmodule
module acsZ0_40_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_7,acs_prob_tdata_6,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_35,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1691_p_O_FD,p_desc1692_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1721_p_O_FDRE);
input branch_tlast ;
output [35:35] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_7 ;
input [8:0] acs_prob_tdata_6 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_35 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIH3MV_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIK7D91 ;
wire un4_v_high_s_7_40 ;
wire un4_v_low_s_7_40 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_40 ;
wire un4_v_low_s_8_40 ;
wire un4_v_high_s_6_40 ;
wire un4_v_low_s_6_40 ;
wire un4_v_high_s_5_40 ;
wire un4_v_low_s_5_40 ;
wire un4_v_high_s_4_40 ;
wire un4_v_low_s_4_40 ;
wire un4_v_high_s_3_40 ;
wire un4_v_low_s_3_40 ;
wire un4_v_high_s_2_40 ;
wire un4_v_low_s_2_40 ;
wire un4_v_high_s_1_40 ;
wire un4_v_low_s_1_40 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1548 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1691_p_O_FD ;
input p_desc1692_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1721_p_O_FDRE ;
// instances
  FDR desc1685(.Q(acs_prob_tdata_35[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  FDR desc1686(.Q(acs_prob_tdata_35[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  FDR desc1687(.Q(acs_prob_tdata_35[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  FDR desc1688(.Q(acs_prob_tdata_35[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  FDR desc1689(.Q(acs_prob_tdata_35[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  FDR desc1690(.Q(acs_prob_tdata_35[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91));
  p_O_FD desc1691(.Q(acs_prob_tdata_35[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1691_p_O_FD));
  p_O_FD desc1692(.Q(acs_prob_tdata_35[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1692_p_O_FD));
  LUT6 desc1693(.I0(un4_v_high_s_7_40),.I1(un4_v_low_s_7_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK7D91),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1693.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1694(.I0(un4_v_high_s_8_40),.I1(un4_v_low_s_8_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK7D91),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1694.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1695(.I0(un4_v_high_s_6_40),.I1(un4_v_low_s_6_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1695.INIT=32'hACACFF00;
  LUT5 desc1696(.I0(un4_v_high_s_5_40),.I1(un4_v_low_s_5_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1696.INIT=32'hACACFF00;
  LUT5 desc1697(.I0(un4_v_high_s_4_40),.I1(un4_v_low_s_4_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1697.INIT=32'hACACFF00;
  LUT5 desc1698(.I0(un4_v_high_s_3_40),.I1(un4_v_low_s_3_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1698.INIT=32'hACACFF00;
  LUT5 desc1699(.I0(un4_v_high_s_2_40),.I1(un4_v_low_s_2_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1699.INIT=32'hACACFF00;
  LUT5 desc1700(.I0(un4_v_high_s_1_40),.I1(un4_v_low_s_1_40),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_35[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1700.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[35:35]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1701(.I0(acs_prob_tdata_6[0:0]),.I1(acs_prob_tdata_7[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1701.INIT=16'h9669;
  LUT2 desc1702(.I0(un4_v_high_s_1_40),.I1(un4_v_low_s_1_40),.O(v_diff_1_axb_1));
defparam desc1702.INIT=4'h9;
  LUT2 desc1703(.I0(un4_v_high_s_2_40),.I1(un4_v_low_s_2_40),.O(v_diff_1_axb_2));
defparam desc1703.INIT=4'h9;
  LUT2 desc1704(.I0(un4_v_high_s_3_40),.I1(un4_v_low_s_3_40),.O(v_diff_1_axb_3));
defparam desc1704.INIT=4'h9;
  LUT2 desc1705(.I0(un4_v_high_s_4_40),.I1(un4_v_low_s_4_40),.O(v_diff_1_axb_4));
defparam desc1705.INIT=4'h9;
  LUT2 desc1706(.I0(un4_v_high_s_5_40),.I1(un4_v_low_s_5_40),.O(v_diff_1_axb_5));
defparam desc1706.INIT=4'h9;
  LUT2 desc1707(.I0(un4_v_high_s_6_40),.I1(un4_v_low_s_6_40),.O(v_diff_1_axb_6));
defparam desc1707.INIT=4'h9;
  LUT2 desc1708(.I0(un4_v_high_s_7_40),.I1(un4_v_low_s_7_40),.O(v_diff_1_axb_7));
defparam desc1708.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_6[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_6[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_6[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_6[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_6[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_6[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_6[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_7[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_7[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_7[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_7[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_7[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_7[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_7[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_7[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1709(.I0(acs_prob_tdata_6[0:0]),.I1(acs_prob_tdata_7[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1548));
defparam desc1709.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_7[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_6[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1710(.I0(un4_v_high_s_8_40),.I1(un4_v_low_s_8_40),.O(v_diff_1_axb_8));
defparam desc1710.INIT=4'h9;
  LUT6 desc1711(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1711.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI25861(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI25861.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIK7D91_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIK7D91));
defparam s_axis_inbranch_tlast_d_RNIK7D91_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_6[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIH3MV_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_40));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_40));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_7[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_40));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_7[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_40));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_7[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_40));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_7[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_40));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_7[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_40));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_7[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_40));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_7[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_7[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_40));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_40));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_6[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_40));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_6[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_40));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_6[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_40));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_6[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_40));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_6[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_40));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_6[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_40));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_6[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_6[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1712(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1713(.DI(un4_v_low_s_7_40),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1714(.DI(un4_v_low_s_6_40),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1715(.DI(un4_v_low_s_5_40),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1716(.DI(un4_v_low_s_4_40),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1717(.DI(un4_v_low_s_3_40),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1718(.DI(un4_v_low_s_2_40),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1719(.DI(un4_v_low_s_1_40),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1720(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1721(.Q(acs_prob_tdata_35[0:0]),.D(N_1548),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK7D91),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1721_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1722(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIH3MV_O6));
defparam desc1722.INIT=16'hF4F0;
  LUT2 desc1723(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1723.INIT=4'h8;
endmodule
module acsZ0_41_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_13,acs_prob_tdata_12,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_6,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1730_p_O_FD,p_desc1731_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1760_p_O_FDRE);
input branch_tlast ;
output [6:6] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_13 ;
input [8:0] acs_prob_tdata_12 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_6 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIRVDG1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIGCUH1 ;
wire un4_v_high_s_7_41 ;
wire un4_v_low_s_7_41 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_41 ;
wire un4_v_low_s_8_41 ;
wire un4_v_high_s_6_41 ;
wire un4_v_low_s_6_41 ;
wire un4_v_high_s_5_41 ;
wire un4_v_low_s_5_41 ;
wire un4_v_high_s_4_41 ;
wire un4_v_low_s_4_41 ;
wire un4_v_high_s_3_41 ;
wire un4_v_low_s_3_41 ;
wire un4_v_high_s_2_41 ;
wire un4_v_low_s_2_41 ;
wire un4_v_high_s_1_41 ;
wire un4_v_low_s_1_41 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1528 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1730_p_O_FD ;
input p_desc1731_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1760_p_O_FDRE ;
// instances
  FDR desc1724(.Q(acs_prob_tdata_6[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  FDR desc1725(.Q(acs_prob_tdata_6[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  FDR desc1726(.Q(acs_prob_tdata_6[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  FDR desc1727(.Q(acs_prob_tdata_6[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  FDR desc1728(.Q(acs_prob_tdata_6[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  FDR desc1729(.Q(acs_prob_tdata_6[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1));
  p_O_FD desc1730(.Q(acs_prob_tdata_6[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1730_p_O_FD));
  p_O_FD desc1731(.Q(acs_prob_tdata_6[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1731_p_O_FD));
  LUT6 desc1732(.I0(un4_v_high_s_7_41),.I1(un4_v_low_s_7_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGCUH1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1732.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1733(.I0(un4_v_high_s_8_41),.I1(un4_v_low_s_8_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGCUH1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1733.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1734(.I0(un4_v_high_s_6_41),.I1(un4_v_low_s_6_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1734.INIT=32'hACACFF00;
  LUT5 desc1735(.I0(un4_v_high_s_5_41),.I1(un4_v_low_s_5_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1735.INIT=32'hACACFF00;
  LUT5 desc1736(.I0(un4_v_high_s_4_41),.I1(un4_v_low_s_4_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1736.INIT=32'hACACFF00;
  LUT5 desc1737(.I0(un4_v_high_s_3_41),.I1(un4_v_low_s_3_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1737.INIT=32'hACACFF00;
  LUT5 desc1738(.I0(un4_v_high_s_2_41),.I1(un4_v_low_s_2_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1738.INIT=32'hACACFF00;
  LUT5 desc1739(.I0(un4_v_high_s_1_41),.I1(un4_v_low_s_1_41),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_6[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1739.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[6:6]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1740(.I0(acs_prob_tdata_12[0:0]),.I1(acs_prob_tdata_13[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1740.INIT=16'h9669;
  LUT2 desc1741(.I0(un4_v_high_s_1_41),.I1(un4_v_low_s_1_41),.O(v_diff_1_axb_1));
defparam desc1741.INIT=4'h9;
  LUT2 desc1742(.I0(un4_v_high_s_2_41),.I1(un4_v_low_s_2_41),.O(v_diff_1_axb_2));
defparam desc1742.INIT=4'h9;
  LUT2 desc1743(.I0(un4_v_high_s_3_41),.I1(un4_v_low_s_3_41),.O(v_diff_1_axb_3));
defparam desc1743.INIT=4'h9;
  LUT2 desc1744(.I0(un4_v_high_s_4_41),.I1(un4_v_low_s_4_41),.O(v_diff_1_axb_4));
defparam desc1744.INIT=4'h9;
  LUT2 desc1745(.I0(un4_v_high_s_5_41),.I1(un4_v_low_s_5_41),.O(v_diff_1_axb_5));
defparam desc1745.INIT=4'h9;
  LUT2 desc1746(.I0(un4_v_high_s_6_41),.I1(un4_v_low_s_6_41),.O(v_diff_1_axb_6));
defparam desc1746.INIT=4'h9;
  LUT2 desc1747(.I0(un4_v_high_s_7_41),.I1(un4_v_low_s_7_41),.O(v_diff_1_axb_7));
defparam desc1747.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_12[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_12[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_12[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_12[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_12[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_12[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_12[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_13[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_13[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_13[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_13[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_13[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_13[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_13[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_13[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1748(.I0(acs_prob_tdata_12[0:0]),.I1(acs_prob_tdata_13[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1528));
defparam desc1748.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_13[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_12[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1749(.I0(un4_v_high_s_8_41),.I1(un4_v_low_s_8_41),.O(v_diff_1_axb_8));
defparam desc1749.INIT=4'h9;
  LUT6 desc1750(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1750.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIU9PE1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIU9PE1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIGCUH1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIGCUH1));
defparam s_axis_inbranch_tlast_d_RNIGCUH1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_12[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIRVDG1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_41));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_41));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_13[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_41));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_13[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_41));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_13[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_41));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_13[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_41));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_13[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_41));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_13[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_41));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_13[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_13[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_41));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_41));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_12[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_41));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_12[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_41));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_12[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_41));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_12[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_41));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_12[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_41));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_12[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_41));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_12[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_12[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1751(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1752(.DI(un4_v_low_s_7_41),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1753(.DI(un4_v_low_s_6_41),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1754(.DI(un4_v_low_s_5_41),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1755(.DI(un4_v_low_s_4_41),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1756(.DI(un4_v_low_s_3_41),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1757(.DI(un4_v_low_s_2_41),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1758(.DI(un4_v_low_s_1_41),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1759(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1760(.Q(acs_prob_tdata_6[0:0]),.D(N_1528),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGCUH1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1760_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1761(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIRVDG1_O6));
defparam desc1761.INIT=16'hF4F0;
  LUT2 desc1762(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1762.INIT=4'h8;
endmodule
module acsZ0_42_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_33,acs_prob_tdata_32,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_48,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,N_1756_1,aresetn,p_desc1769_p_O_FD,p_desc1770_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1799_p_O_FDRE);
input branch_tlast ;
output [48:48] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_33 ;
input [8:0] acs_prob_tdata_32 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_48 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNITUAR_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNISLS41 ;
wire un4_v_high_s_7_42 ;
wire un4_v_low_s_7_42 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_42 ;
wire un4_v_low_s_8_42 ;
wire un4_v_high_s_6_42 ;
wire un4_v_low_s_6_42 ;
wire un4_v_high_s_5_42 ;
wire un4_v_low_s_5_42 ;
wire un4_v_high_s_4_42 ;
wire un4_v_low_s_4_42 ;
wire un4_v_high_s_3_42 ;
wire un4_v_low_s_3_42 ;
wire un4_v_high_s_2_42 ;
wire un4_v_low_s_2_42 ;
wire un4_v_high_s_1_42 ;
wire un4_v_low_s_1_42 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1508 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1769_p_O_FD ;
input p_desc1770_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1799_p_O_FDRE ;
// instances
  FDR desc1763(.Q(acs_prob_tdata_48[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  FDR desc1764(.Q(acs_prob_tdata_48[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  FDR desc1765(.Q(acs_prob_tdata_48[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  FDR desc1766(.Q(acs_prob_tdata_48[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  FDR desc1767(.Q(acs_prob_tdata_48[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  FDR desc1768(.Q(acs_prob_tdata_48[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41));
  p_O_FD desc1769(.Q(acs_prob_tdata_48[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1769_p_O_FD));
  p_O_FD desc1770(.Q(acs_prob_tdata_48[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1770_p_O_FD));
  LUT6 desc1771(.I0(un4_v_high_s_7_42),.I1(un4_v_low_s_7_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISLS41),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1771.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1772(.I0(un4_v_high_s_8_42),.I1(un4_v_low_s_8_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNISLS41),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1772.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1773(.I0(un4_v_high_s_6_42),.I1(un4_v_low_s_6_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1773.INIT=32'hACACFF00;
  LUT5 desc1774(.I0(un4_v_high_s_5_42),.I1(un4_v_low_s_5_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1774.INIT=32'hACACFF00;
  LUT5 desc1775(.I0(un4_v_high_s_4_42),.I1(un4_v_low_s_4_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1775.INIT=32'hACACFF00;
  LUT5 desc1776(.I0(un4_v_high_s_3_42),.I1(un4_v_low_s_3_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1776.INIT=32'hACACFF00;
  LUT5 desc1777(.I0(un4_v_high_s_2_42),.I1(un4_v_low_s_2_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1777.INIT=32'hACACFF00;
  LUT5 desc1778(.I0(un4_v_high_s_1_42),.I1(un4_v_low_s_1_42),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_48[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1778.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[48:48]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_32[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_32[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_32[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_32[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_32[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_32[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_32[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_33[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_33[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_33[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_33[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_33[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_33[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_33[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_33[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1779(.I0(acs_prob_tdata_32[0:0]),.I1(acs_prob_tdata_33[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1779.INIT=16'h9669;
  LUT2 desc1780(.I0(un4_v_high_s_1_42),.I1(un4_v_low_s_1_42),.O(v_diff_1_axb_1));
defparam desc1780.INIT=4'h9;
  LUT2 desc1781(.I0(un4_v_high_s_2_42),.I1(un4_v_low_s_2_42),.O(v_diff_1_axb_2));
defparam desc1781.INIT=4'h9;
  LUT2 desc1782(.I0(un4_v_high_s_3_42),.I1(un4_v_low_s_3_42),.O(v_diff_1_axb_3));
defparam desc1782.INIT=4'h9;
  LUT2 desc1783(.I0(un4_v_high_s_4_42),.I1(un4_v_low_s_4_42),.O(v_diff_1_axb_4));
defparam desc1783.INIT=4'h9;
  LUT2 desc1784(.I0(un4_v_high_s_5_42),.I1(un4_v_low_s_5_42),.O(v_diff_1_axb_5));
defparam desc1784.INIT=4'h9;
  LUT2 desc1785(.I0(un4_v_high_s_6_42),.I1(un4_v_low_s_6_42),.O(v_diff_1_axb_6));
defparam desc1785.INIT=4'h9;
  LUT2 desc1786(.I0(un4_v_high_s_7_42),.I1(un4_v_low_s_7_42),.O(v_diff_1_axb_7));
defparam desc1786.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1787(.I0(acs_prob_tdata_32[0:0]),.I1(acs_prob_tdata_33[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1508));
defparam desc1787.INIT=32'h33CC5A5A;
  LUT2 desc1788(.I0(un4_v_high_s_8_42),.I1(un4_v_low_s_8_42),.O(v_diff_1_axb_8));
defparam desc1788.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_33[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_32[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1789(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1789.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIAJN11(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIAJN11.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNISLS41_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNISLS41));
defparam s_axis_inbranch_tlast_d_RNISLS41_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_32[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNITUAR_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1790(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1791(.DI(un4_v_low_s_7_42),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1792(.DI(un4_v_low_s_6_42),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1793(.DI(un4_v_low_s_5_42),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1794(.DI(un4_v_low_s_4_42),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1795(.DI(un4_v_low_s_3_42),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1796(.DI(un4_v_low_s_2_42),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1797(.DI(un4_v_low_s_1_42),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1798(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_42));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_42));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_33[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_42));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_33[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_42));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_33[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_42));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_33[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_42));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_33[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_42));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_33[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_42));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_33[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_33[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_42));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_42));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_32[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_42));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_32[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_42));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_32[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_42));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_32[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_42));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_32[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_42));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_32[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_42));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_32[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_32[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1799(.Q(acs_prob_tdata_48[0:0]),.D(N_1508),.C(aclk),.R(s_axis_inbranch_tlast_d_RNISLS41),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1799_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1800(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNITUAR_O6));
defparam desc1800.INIT=16'hF4F0;
  LUT2 desc1801(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1801.INIT=4'h8;
endmodule
module acsZ0_43_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_41,acs_prob_tdata_40,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_20,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1808_p_O_FD,p_desc1809_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1838_p_O_FDRE);
input branch_tlast ;
output [20:20] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_41 ;
input [8:0] acs_prob_tdata_40 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_20 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIVR1U_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI8JN91 ;
wire un4_v_high_s_7_43 ;
wire un4_v_low_s_7_43 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_43 ;
wire un4_v_low_s_8_43 ;
wire un4_v_high_s_6_43 ;
wire un4_v_low_s_6_43 ;
wire un4_v_high_s_5_43 ;
wire un4_v_low_s_5_43 ;
wire un4_v_high_s_4_43 ;
wire un4_v_low_s_4_43 ;
wire un4_v_high_s_3_43 ;
wire un4_v_low_s_3_43 ;
wire un4_v_high_s_2_43 ;
wire un4_v_low_s_2_43 ;
wire un4_v_high_s_1_43 ;
wire un4_v_low_s_1_43 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1488 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc1808_p_O_FD ;
input p_desc1809_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1838_p_O_FDRE ;
// instances
  FDR desc1802(.Q(acs_prob_tdata_20[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  FDR desc1803(.Q(acs_prob_tdata_20[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  FDR desc1804(.Q(acs_prob_tdata_20[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  FDR desc1805(.Q(acs_prob_tdata_20[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  FDR desc1806(.Q(acs_prob_tdata_20[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  FDR desc1807(.Q(acs_prob_tdata_20[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91));
  p_O_FD desc1808(.Q(acs_prob_tdata_20[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1808_p_O_FD));
  p_O_FD desc1809(.Q(acs_prob_tdata_20[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1809_p_O_FD));
  LUT6 desc1810(.I0(un4_v_high_s_7_43),.I1(un4_v_low_s_7_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI8JN91),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1810.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1811(.I0(un4_v_high_s_8_43),.I1(un4_v_low_s_8_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI8JN91),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1811.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1812(.I0(un4_v_high_s_6_43),.I1(un4_v_low_s_6_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1812.INIT=32'hACACFF00;
  LUT5 desc1813(.I0(un4_v_high_s_5_43),.I1(un4_v_low_s_5_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1813.INIT=32'hACACFF00;
  LUT5 desc1814(.I0(un4_v_high_s_4_43),.I1(un4_v_low_s_4_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1814.INIT=32'hACACFF00;
  LUT5 desc1815(.I0(un4_v_high_s_3_43),.I1(un4_v_low_s_3_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1815.INIT=32'hACACFF00;
  LUT5 desc1816(.I0(un4_v_high_s_2_43),.I1(un4_v_low_s_2_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1816.INIT=32'hACACFF00;
  LUT5 desc1817(.I0(un4_v_high_s_1_43),.I1(un4_v_low_s_1_43),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_20[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1817.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[20:20]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_40[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_40[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_40[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_40[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_40[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_40[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_40[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_41[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_41[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_41[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_41[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_41[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_41[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_41[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_41[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc1818(.I0(acs_prob_tdata_40[0:0]),.I1(acs_prob_tdata_41[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1818.INIT=16'h9669;
  LUT2 desc1819(.I0(un4_v_high_s_1_43),.I1(un4_v_low_s_1_43),.O(v_diff_1_axb_1));
defparam desc1819.INIT=4'h9;
  LUT2 desc1820(.I0(un4_v_high_s_2_43),.I1(un4_v_low_s_2_43),.O(v_diff_1_axb_2));
defparam desc1820.INIT=4'h9;
  LUT2 desc1821(.I0(un4_v_high_s_3_43),.I1(un4_v_low_s_3_43),.O(v_diff_1_axb_3));
defparam desc1821.INIT=4'h9;
  LUT2 desc1822(.I0(un4_v_high_s_4_43),.I1(un4_v_low_s_4_43),.O(v_diff_1_axb_4));
defparam desc1822.INIT=4'h9;
  LUT2 desc1823(.I0(un4_v_high_s_5_43),.I1(un4_v_low_s_5_43),.O(v_diff_1_axb_5));
defparam desc1823.INIT=4'h9;
  LUT2 desc1824(.I0(un4_v_high_s_6_43),.I1(un4_v_low_s_6_43),.O(v_diff_1_axb_6));
defparam desc1824.INIT=4'h9;
  LUT2 desc1825(.I0(un4_v_high_s_7_43),.I1(un4_v_low_s_7_43),.O(v_diff_1_axb_7));
defparam desc1825.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1826(.I0(acs_prob_tdata_40[0:0]),.I1(acs_prob_tdata_41[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1488));
defparam desc1826.INIT=32'h33CC5A5A;
  LUT2 desc1827(.I0(un4_v_high_s_8_43),.I1(un4_v_low_s_8_43),.O(v_diff_1_axb_8));
defparam desc1827.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_41[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_40[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc1828(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1828.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIMGI61(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIMGI61.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI8JN91_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI8JN91));
defparam s_axis_inbranch_tlast_d_RNI8JN91_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_40[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIVR1U_O6),.C(aclk),.R(aresetn_i));
  XORCY desc1829(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1830(.DI(un4_v_low_s_7_43),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1831(.DI(un4_v_low_s_6_43),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1832(.DI(un4_v_low_s_5_43),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1833(.DI(un4_v_low_s_4_43),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1834(.DI(un4_v_low_s_3_43),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1835(.DI(un4_v_low_s_2_43),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1836(.DI(un4_v_low_s_1_43),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1837(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_43));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_43));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_41[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_43));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_41[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_43));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_41[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_43));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_41[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_43));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_41[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_43));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_41[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_43));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_41[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_41[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_43));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_43));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_40[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_43));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_40[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_43));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_40[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_43));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_40[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_43));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_40[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_43));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_40[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_43));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_40[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_40[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc1838(.Q(acs_prob_tdata_20[0:0]),.D(N_1488),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI8JN91),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1838_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1839(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIVR1U_O6));
defparam desc1839.INIT=16'hF4F0;
  LUT2 desc1840(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1840.INIT=4'h8;
endmodule
module acsZ0_44_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_13,acs_prob_tdata_12,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_38,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc1847_p_O_FD,p_desc1848_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1877_p_O_FDRE);
input branch_tlast ;
output [38:38] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_13 ;
input [8:0] acs_prob_tdata_12 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_38 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIQ5LO_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIQGMV ;
wire un4_v_high_s_7_44 ;
wire un4_v_low_s_7_44 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_44 ;
wire un4_v_low_s_8_44 ;
wire un4_v_high_s_6_44 ;
wire un4_v_low_s_6_44 ;
wire un4_v_high_s_5_44 ;
wire un4_v_low_s_5_44 ;
wire un4_v_high_s_4_44 ;
wire un4_v_low_s_4_44 ;
wire un4_v_high_s_3_44 ;
wire un4_v_low_s_3_44 ;
wire un4_v_high_s_2_44 ;
wire un4_v_low_s_2_44 ;
wire un4_v_high_s_1_44 ;
wire un4_v_low_s_1_44 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1468 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1847_p_O_FD ;
input p_desc1848_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1877_p_O_FDRE ;
// instances
  FDR desc1841(.Q(acs_prob_tdata_38[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  FDR desc1842(.Q(acs_prob_tdata_38[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  FDR desc1843(.Q(acs_prob_tdata_38[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  FDR desc1844(.Q(acs_prob_tdata_38[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  FDR desc1845(.Q(acs_prob_tdata_38[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  FDR desc1846(.Q(acs_prob_tdata_38[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV));
  p_O_FD desc1847(.Q(acs_prob_tdata_38[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1847_p_O_FD));
  p_O_FD desc1848(.Q(acs_prob_tdata_38[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1848_p_O_FD));
  LUT6 desc1849(.I0(un4_v_high_s_7_44),.I1(un4_v_low_s_7_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQGMV),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1849.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1850(.I0(un4_v_high_s_8_44),.I1(un4_v_low_s_8_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQGMV),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1850.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1851(.I0(un4_v_high_s_6_44),.I1(un4_v_low_s_6_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1851.INIT=32'hACACFF00;
  LUT5 desc1852(.I0(un4_v_high_s_5_44),.I1(un4_v_low_s_5_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1852.INIT=32'hACACFF00;
  LUT5 desc1853(.I0(un4_v_high_s_4_44),.I1(un4_v_low_s_4_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1853.INIT=32'hACACFF00;
  LUT5 desc1854(.I0(un4_v_high_s_3_44),.I1(un4_v_low_s_3_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1854.INIT=32'hACACFF00;
  LUT5 desc1855(.I0(un4_v_high_s_2_44),.I1(un4_v_low_s_2_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1855.INIT=32'hACACFF00;
  LUT5 desc1856(.I0(un4_v_high_s_1_44),.I1(un4_v_low_s_1_44),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_38[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1856.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[38:38]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1857(.I0(acs_prob_tdata_12[0:0]),.I1(acs_prob_tdata_13[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc1857.INIT=16'h9669;
  LUT2 desc1858(.I0(un4_v_high_s_1_44),.I1(un4_v_low_s_1_44),.O(v_diff_1_axb_1));
defparam desc1858.INIT=4'h9;
  LUT2 desc1859(.I0(un4_v_high_s_2_44),.I1(un4_v_low_s_2_44),.O(v_diff_1_axb_2));
defparam desc1859.INIT=4'h9;
  LUT2 desc1860(.I0(un4_v_high_s_3_44),.I1(un4_v_low_s_3_44),.O(v_diff_1_axb_3));
defparam desc1860.INIT=4'h9;
  LUT2 desc1861(.I0(un4_v_high_s_4_44),.I1(un4_v_low_s_4_44),.O(v_diff_1_axb_4));
defparam desc1861.INIT=4'h9;
  LUT2 desc1862(.I0(un4_v_high_s_5_44),.I1(un4_v_low_s_5_44),.O(v_diff_1_axb_5));
defparam desc1862.INIT=4'h9;
  LUT2 desc1863(.I0(un4_v_high_s_6_44),.I1(un4_v_low_s_6_44),.O(v_diff_1_axb_6));
defparam desc1863.INIT=4'h9;
  LUT2 desc1864(.I0(un4_v_high_s_7_44),.I1(un4_v_low_s_7_44),.O(v_diff_1_axb_7));
defparam desc1864.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_12[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_12[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_12[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_12[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_12[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_12[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_12[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_13[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_13[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_13[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_13[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_13[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_13[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_13[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_13[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1865(.I0(acs_prob_tdata_12[0:0]),.I1(acs_prob_tdata_13[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1468));
defparam desc1865.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_13[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_12[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1866(.I0(un4_v_high_s_8_44),.I1(un4_v_low_s_8_44),.O(v_diff_1_axb_8));
defparam desc1866.INIT=4'h9;
  LUT6 desc1867(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1867.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI8EHS(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI8EHS.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIQGMV_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIQGMV));
defparam s_axis_inbranch_tlast_d_RNIQGMV_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_12[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIQ5LO_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_44));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_44));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_13[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_44));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_13[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_44));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_13[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_44));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_13[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_44));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_13[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_44));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_13[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_44));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_13[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_13[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_44));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_44));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_12[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_44));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_12[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_44));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_12[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_44));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_12[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_44));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_12[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_44));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_12[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_44));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_12[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_12[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1868(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1869(.DI(un4_v_low_s_7_44),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1870(.DI(un4_v_low_s_6_44),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1871(.DI(un4_v_low_s_5_44),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1872(.DI(un4_v_low_s_4_44),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1873(.DI(un4_v_low_s_3_44),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1874(.DI(un4_v_low_s_2_44),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1875(.DI(un4_v_low_s_1_44),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1876(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1877(.Q(acs_prob_tdata_38[0:0]),.D(N_1468),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQGMV),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1877_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1878(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIQ5LO_O6));
defparam desc1878.INIT=16'hF4F0;
  LUT2 desc1879(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1879.INIT=4'h8;
endmodule
module acsZ0_45_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_19,acs_prob_tdata_18,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_41,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc1886_p_O_FD,p_desc1887_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1916_p_O_FDRE);
input branch_tlast ;
output [41:41] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_19 ;
input [8:0] acs_prob_tdata_18 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_41 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI84D61_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIE0761 ;
wire un4_v_high_s_7_45 ;
wire un4_v_low_s_7_45 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_45 ;
wire un4_v_low_s_8_45 ;
wire un4_v_high_s_6_45 ;
wire un4_v_low_s_6_45 ;
wire un4_v_high_s_5_45 ;
wire un4_v_low_s_5_45 ;
wire un4_v_high_s_4_45 ;
wire un4_v_low_s_4_45 ;
wire un4_v_high_s_3_45 ;
wire un4_v_low_s_3_45 ;
wire un4_v_high_s_2_45 ;
wire un4_v_low_s_2_45 ;
wire un4_v_high_s_1_45 ;
wire un4_v_low_s_1_45 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1448 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1886_p_O_FD ;
input p_desc1887_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1916_p_O_FDRE ;
// instances
  FDR desc1880(.Q(acs_prob_tdata_41[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  FDR desc1881(.Q(acs_prob_tdata_41[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  FDR desc1882(.Q(acs_prob_tdata_41[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  FDR desc1883(.Q(acs_prob_tdata_41[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  FDR desc1884(.Q(acs_prob_tdata_41[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  FDR desc1885(.Q(acs_prob_tdata_41[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761));
  p_O_FD desc1886(.Q(acs_prob_tdata_41[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1886_p_O_FD));
  p_O_FD desc1887(.Q(acs_prob_tdata_41[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1887_p_O_FD));
  LUT6 desc1888(.I0(un4_v_high_s_7_45),.I1(un4_v_low_s_7_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE0761),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1888.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1889(.I0(un4_v_high_s_8_45),.I1(un4_v_low_s_8_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIE0761),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1889.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1890(.I0(un4_v_high_s_6_45),.I1(un4_v_low_s_6_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1890.INIT=32'hACACFF00;
  LUT5 desc1891(.I0(un4_v_high_s_5_45),.I1(un4_v_low_s_5_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1891.INIT=32'hACACFF00;
  LUT5 desc1892(.I0(un4_v_high_s_4_45),.I1(un4_v_low_s_4_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1892.INIT=32'hACACFF00;
  LUT5 desc1893(.I0(un4_v_high_s_3_45),.I1(un4_v_low_s_3_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1893.INIT=32'hACACFF00;
  LUT5 desc1894(.I0(un4_v_high_s_2_45),.I1(un4_v_low_s_2_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1894.INIT=32'hACACFF00;
  LUT5 desc1895(.I0(un4_v_high_s_1_45),.I1(un4_v_low_s_1_45),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_41[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1895.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[41:41]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1896(.I0(acs_prob_tdata_18[0:0]),.I1(acs_prob_tdata_19[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1896.INIT=16'h9669;
  LUT2 desc1897(.I0(un4_v_high_s_1_45),.I1(un4_v_low_s_1_45),.O(v_diff_1_axb_1));
defparam desc1897.INIT=4'h9;
  LUT2 desc1898(.I0(un4_v_high_s_2_45),.I1(un4_v_low_s_2_45),.O(v_diff_1_axb_2));
defparam desc1898.INIT=4'h9;
  LUT2 desc1899(.I0(un4_v_high_s_3_45),.I1(un4_v_low_s_3_45),.O(v_diff_1_axb_3));
defparam desc1899.INIT=4'h9;
  LUT2 desc1900(.I0(un4_v_high_s_4_45),.I1(un4_v_low_s_4_45),.O(v_diff_1_axb_4));
defparam desc1900.INIT=4'h9;
  LUT2 desc1901(.I0(un4_v_high_s_5_45),.I1(un4_v_low_s_5_45),.O(v_diff_1_axb_5));
defparam desc1901.INIT=4'h9;
  LUT2 desc1902(.I0(un4_v_high_s_6_45),.I1(un4_v_low_s_6_45),.O(v_diff_1_axb_6));
defparam desc1902.INIT=4'h9;
  LUT2 desc1903(.I0(un4_v_high_s_7_45),.I1(un4_v_low_s_7_45),.O(v_diff_1_axb_7));
defparam desc1903.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_18[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_18[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_18[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_18[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_18[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_18[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_18[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_19[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_19[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_19[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_19[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_19[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_19[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_19[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_19[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1904(.I0(acs_prob_tdata_18[0:0]),.I1(acs_prob_tdata_19[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1448));
defparam desc1904.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_19[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_18[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1905(.I0(un4_v_high_s_8_45),.I1(un4_v_low_s_8_45),.O(v_diff_1_axb_8));
defparam desc1905.INIT=4'h9;
  LUT6 desc1906(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1906.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIST131(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIST131.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIE0761_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIE0761));
defparam s_axis_inbranch_tlast_d_RNIE0761_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_18[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI84D61_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_45));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_45));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_19[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_45));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_19[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_45));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_19[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_45));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_19[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_45));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_19[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_45));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_19[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_45));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_19[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_19[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_45));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_45));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_18[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_45));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_18[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_45));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_18[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_45));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_18[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_45));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_18[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_45));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_18[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_45));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_18[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_18[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1907(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1908(.DI(un4_v_low_s_7_45),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1909(.DI(un4_v_low_s_6_45),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1910(.DI(un4_v_low_s_5_45),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1911(.DI(un4_v_low_s_4_45),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1912(.DI(un4_v_low_s_3_45),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1913(.DI(un4_v_low_s_2_45),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1914(.DI(un4_v_low_s_1_45),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1915(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1916(.Q(acs_prob_tdata_41[0:0]),.D(N_1448),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIE0761),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1916_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1917(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI84D61_O6));
defparam desc1917.INIT=16'hF4F0;
  LUT2 desc1918(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1918.INIT=4'h8;
endmodule
module acsZ0_46_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_53,acs_prob_tdata_52,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_26,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc1925_p_O_FD,p_desc1926_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1955_p_O_FDRE);
input branch_tlast ;
output [26:26] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_53 ;
input [8:0] acs_prob_tdata_52 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_26 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIH0001_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIK5A61 ;
wire un4_v_high_s_7_46 ;
wire un4_v_low_s_7_46 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_46 ;
wire un4_v_low_s_8_46 ;
wire un4_v_high_s_6_46 ;
wire un4_v_low_s_6_46 ;
wire un4_v_high_s_5_46 ;
wire un4_v_low_s_5_46 ;
wire un4_v_high_s_4_46 ;
wire un4_v_low_s_4_46 ;
wire un4_v_high_s_3_46 ;
wire un4_v_low_s_3_46 ;
wire un4_v_high_s_2_46 ;
wire un4_v_low_s_2_46 ;
wire un4_v_high_s_1_46 ;
wire un4_v_low_s_1_46 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1428 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1925_p_O_FD ;
input p_desc1926_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1955_p_O_FDRE ;
// instances
  FDR desc1919(.Q(acs_prob_tdata_26[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  FDR desc1920(.Q(acs_prob_tdata_26[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  FDR desc1921(.Q(acs_prob_tdata_26[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  FDR desc1922(.Q(acs_prob_tdata_26[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  FDR desc1923(.Q(acs_prob_tdata_26[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  FDR desc1924(.Q(acs_prob_tdata_26[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61));
  p_O_FD desc1925(.Q(acs_prob_tdata_26[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1925_p_O_FD));
  p_O_FD desc1926(.Q(acs_prob_tdata_26[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1926_p_O_FD));
  LUT6 desc1927(.I0(un4_v_high_s_7_46),.I1(un4_v_low_s_7_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK5A61),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1927.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1928(.I0(un4_v_high_s_8_46),.I1(un4_v_low_s_8_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK5A61),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1928.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1929(.I0(un4_v_high_s_6_46),.I1(un4_v_low_s_6_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1929.INIT=32'hACACFF00;
  LUT5 desc1930(.I0(un4_v_high_s_5_46),.I1(un4_v_low_s_5_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1930.INIT=32'hACACFF00;
  LUT5 desc1931(.I0(un4_v_high_s_4_46),.I1(un4_v_low_s_4_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1931.INIT=32'hACACFF00;
  LUT5 desc1932(.I0(un4_v_high_s_3_46),.I1(un4_v_low_s_3_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1932.INIT=32'hACACFF00;
  LUT5 desc1933(.I0(un4_v_high_s_2_46),.I1(un4_v_low_s_2_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1933.INIT=32'hACACFF00;
  LUT5 desc1934(.I0(un4_v_high_s_1_46),.I1(un4_v_low_s_1_46),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_26[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1934.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[26:26]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1935(.I0(acs_prob_tdata_52[0:0]),.I1(acs_prob_tdata_53[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1935.INIT=16'h9669;
  LUT2 desc1936(.I0(un4_v_high_s_1_46),.I1(un4_v_low_s_1_46),.O(v_diff_1_axb_1));
defparam desc1936.INIT=4'h9;
  LUT2 desc1937(.I0(un4_v_high_s_2_46),.I1(un4_v_low_s_2_46),.O(v_diff_1_axb_2));
defparam desc1937.INIT=4'h9;
  LUT2 desc1938(.I0(un4_v_high_s_3_46),.I1(un4_v_low_s_3_46),.O(v_diff_1_axb_3));
defparam desc1938.INIT=4'h9;
  LUT2 desc1939(.I0(un4_v_high_s_4_46),.I1(un4_v_low_s_4_46),.O(v_diff_1_axb_4));
defparam desc1939.INIT=4'h9;
  LUT2 desc1940(.I0(un4_v_high_s_5_46),.I1(un4_v_low_s_5_46),.O(v_diff_1_axb_5));
defparam desc1940.INIT=4'h9;
  LUT2 desc1941(.I0(un4_v_high_s_6_46),.I1(un4_v_low_s_6_46),.O(v_diff_1_axb_6));
defparam desc1941.INIT=4'h9;
  LUT2 desc1942(.I0(un4_v_high_s_7_46),.I1(un4_v_low_s_7_46),.O(v_diff_1_axb_7));
defparam desc1942.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_52[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_52[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_52[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_52[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_52[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_52[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_52[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_53[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_53[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_53[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_53[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_53[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_53[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_53[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_53[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1943(.I0(acs_prob_tdata_52[0:0]),.I1(acs_prob_tdata_53[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1428));
defparam desc1943.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_53[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_52[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1944(.I0(un4_v_high_s_8_46),.I1(un4_v_low_s_8_46),.O(v_diff_1_axb_8));
defparam desc1944.INIT=4'h9;
  LUT6 desc1945(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1945.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI23531(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI23531.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIK5A61_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIK5A61));
defparam s_axis_inbranch_tlast_d_RNIK5A61_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_52[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIH0001_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_46));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_46));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_53[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_46));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_53[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_46));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_53[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_46));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_53[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_46));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_53[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_46));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_53[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_46));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_53[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_53[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_46));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_46));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_52[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_46));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_52[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_46));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_52[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_46));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_52[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_46));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_52[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_46));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_52[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_46));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_52[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_52[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1946(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1947(.DI(un4_v_low_s_7_46),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1948(.DI(un4_v_low_s_6_46),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1949(.DI(un4_v_low_s_5_46),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1950(.DI(un4_v_low_s_4_46),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1951(.DI(un4_v_low_s_3_46),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1952(.DI(un4_v_low_s_2_46),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1953(.DI(un4_v_low_s_1_46),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1954(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1955(.Q(acs_prob_tdata_26[0:0]),.D(N_1428),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK5A61),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1955_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1956(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIH0001_O6));
defparam desc1956.INIT=16'hF4F0;
  LUT2 desc1957(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1957.INIT=4'h8;
endmodule
module acsZ0_47_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_53,acs_prob_tdata_52,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_58,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,N_1756_1,aresetn,p_desc1964_p_O_FD,p_desc1965_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc1994_p_O_FDRE);
input branch_tlast ;
output [58:58] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_53 ;
input [8:0] acs_prob_tdata_52 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_58 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI0O0E_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIUQ2Q ;
wire un4_v_high_s_7_47 ;
wire un4_v_low_s_7_47 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_47 ;
wire un4_v_low_s_8_47 ;
wire un4_v_high_s_6_47 ;
wire un4_v_low_s_6_47 ;
wire un4_v_high_s_5_47 ;
wire un4_v_low_s_5_47 ;
wire un4_v_high_s_4_47 ;
wire un4_v_low_s_4_47 ;
wire un4_v_high_s_3_47 ;
wire un4_v_low_s_3_47 ;
wire un4_v_high_s_2_47 ;
wire un4_v_low_s_2_47 ;
wire un4_v_high_s_1_47 ;
wire un4_v_low_s_1_47 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1408 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc1964_p_O_FD ;
input p_desc1965_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc1994_p_O_FDRE ;
// instances
  FDR desc1958(.Q(acs_prob_tdata_58[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  FDR desc1959(.Q(acs_prob_tdata_58[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  FDR desc1960(.Q(acs_prob_tdata_58[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  FDR desc1961(.Q(acs_prob_tdata_58[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  FDR desc1962(.Q(acs_prob_tdata_58[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  FDR desc1963(.Q(acs_prob_tdata_58[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q));
  p_O_FD desc1964(.Q(acs_prob_tdata_58[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc1964_p_O_FD));
  p_O_FD desc1965(.Q(acs_prob_tdata_58[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc1965_p_O_FD));
  LUT6 desc1966(.I0(un4_v_high_s_7_47),.I1(un4_v_low_s_7_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIUQ2Q),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc1966.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc1967(.I0(un4_v_high_s_8_47),.I1(un4_v_low_s_8_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIUQ2Q),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc1967.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc1968(.I0(un4_v_high_s_6_47),.I1(un4_v_low_s_6_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc1968.INIT=32'hACACFF00;
  LUT5 desc1969(.I0(un4_v_high_s_5_47),.I1(un4_v_low_s_5_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc1969.INIT=32'hACACFF00;
  LUT5 desc1970(.I0(un4_v_high_s_4_47),.I1(un4_v_low_s_4_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc1970.INIT=32'hACACFF00;
  LUT5 desc1971(.I0(un4_v_high_s_3_47),.I1(un4_v_low_s_3_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc1971.INIT=32'hACACFF00;
  LUT5 desc1972(.I0(un4_v_high_s_2_47),.I1(un4_v_low_s_2_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc1972.INIT=32'hACACFF00;
  LUT5 desc1973(.I0(un4_v_high_s_1_47),.I1(un4_v_low_s_1_47),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_58[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc1973.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[58:58]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc1974(.I0(acs_prob_tdata_52[0:0]),.I1(acs_prob_tdata_53[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc1974.INIT=16'h9669;
  LUT2 desc1975(.I0(un4_v_high_s_1_47),.I1(un4_v_low_s_1_47),.O(v_diff_1_axb_1));
defparam desc1975.INIT=4'h9;
  LUT2 desc1976(.I0(un4_v_high_s_2_47),.I1(un4_v_low_s_2_47),.O(v_diff_1_axb_2));
defparam desc1976.INIT=4'h9;
  LUT2 desc1977(.I0(un4_v_high_s_3_47),.I1(un4_v_low_s_3_47),.O(v_diff_1_axb_3));
defparam desc1977.INIT=4'h9;
  LUT2 desc1978(.I0(un4_v_high_s_4_47),.I1(un4_v_low_s_4_47),.O(v_diff_1_axb_4));
defparam desc1978.INIT=4'h9;
  LUT2 desc1979(.I0(un4_v_high_s_5_47),.I1(un4_v_low_s_5_47),.O(v_diff_1_axb_5));
defparam desc1979.INIT=4'h9;
  LUT2 desc1980(.I0(un4_v_high_s_6_47),.I1(un4_v_low_s_6_47),.O(v_diff_1_axb_6));
defparam desc1980.INIT=4'h9;
  LUT2 desc1981(.I0(un4_v_high_s_7_47),.I1(un4_v_low_s_7_47),.O(v_diff_1_axb_7));
defparam desc1981.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_52[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_52[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_52[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_52[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_52[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_52[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_52[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_53[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_53[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_53[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_53[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_53[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_53[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_53[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_53[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc1982(.I0(acs_prob_tdata_52[0:0]),.I1(acs_prob_tdata_53[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1408));
defparam desc1982.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_53[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_52[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc1983(.I0(un4_v_high_s_8_47),.I1(un4_v_low_s_8_47),.O(v_diff_1_axb_8));
defparam desc1983.INIT=4'h9;
  LUT6 desc1984(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc1984.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNICOTM(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNICOTM.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIUQ2Q_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIUQ2Q));
defparam s_axis_inbranch_tlast_d_RNIUQ2Q_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_52[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI0O0E_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_47));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_47));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_53[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_47));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_53[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_47));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_53[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_47));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_53[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_47));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_53[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_47));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_53[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_47));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_53[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_53[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_47));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_47));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_52[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_47));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_52[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_47));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_52[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_47));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_52[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_47));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_52[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_47));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_52[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_47));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_52[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_52[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc1985(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc1986(.DI(un4_v_low_s_7_47),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc1987(.DI(un4_v_low_s_6_47),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc1988(.DI(un4_v_low_s_5_47),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc1989(.DI(un4_v_low_s_4_47),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc1990(.DI(un4_v_low_s_3_47),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc1991(.DI(un4_v_low_s_2_47),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc1992(.DI(un4_v_low_s_1_47),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc1993(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc1994(.Q(acs_prob_tdata_58[0:0]),.D(N_1408),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIUQ2Q),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc1994_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1995(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI0O0E_O6));
defparam desc1995.INIT=16'hF4F0;
  LUT2 desc1996(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc1996.INIT=4'h8;
endmodule
module acsZ0_48_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_23,acs_prob_tdata_22,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_43,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc2003_p_O_FD,p_desc2004_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2033_p_O_FDRE);
input branch_tlast ;
output [43:43] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_23 ;
input [8:0] acs_prob_tdata_22 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_43 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIEGCC1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNII6DA1 ;
wire un4_v_high_s_7_48 ;
wire un4_v_low_s_7_48 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_48 ;
wire un4_v_low_s_8_48 ;
wire un4_v_high_s_6_48 ;
wire un4_v_low_s_6_48 ;
wire un4_v_high_s_5_48 ;
wire un4_v_low_s_5_48 ;
wire un4_v_high_s_4_48 ;
wire un4_v_low_s_4_48 ;
wire un4_v_high_s_3_48 ;
wire un4_v_low_s_3_48 ;
wire un4_v_high_s_2_48 ;
wire un4_v_low_s_2_48 ;
wire un4_v_high_s_1_48 ;
wire un4_v_low_s_1_48 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1388 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2003_p_O_FD ;
input p_desc2004_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2033_p_O_FDRE ;
// instances
  FDR desc1997(.Q(acs_prob_tdata_43[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  FDR desc1998(.Q(acs_prob_tdata_43[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  FDR desc1999(.Q(acs_prob_tdata_43[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  FDR desc2000(.Q(acs_prob_tdata_43[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  FDR desc2001(.Q(acs_prob_tdata_43[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  FDR desc2002(.Q(acs_prob_tdata_43[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1));
  p_O_FD desc2003(.Q(acs_prob_tdata_43[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2003_p_O_FD));
  p_O_FD desc2004(.Q(acs_prob_tdata_43[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2004_p_O_FD));
  LUT6 desc2005(.I0(un4_v_high_s_7_48),.I1(un4_v_low_s_7_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII6DA1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2005.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2006(.I0(un4_v_high_s_8_48),.I1(un4_v_low_s_8_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNII6DA1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2006.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2007(.I0(un4_v_high_s_6_48),.I1(un4_v_low_s_6_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2007.INIT=32'hACACFF00;
  LUT5 desc2008(.I0(un4_v_high_s_5_48),.I1(un4_v_low_s_5_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2008.INIT=32'hACACFF00;
  LUT5 desc2009(.I0(un4_v_high_s_4_48),.I1(un4_v_low_s_4_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2009.INIT=32'hACACFF00;
  LUT5 desc2010(.I0(un4_v_high_s_3_48),.I1(un4_v_low_s_3_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2010.INIT=32'hACACFF00;
  LUT5 desc2011(.I0(un4_v_high_s_2_48),.I1(un4_v_low_s_2_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2011.INIT=32'hACACFF00;
  LUT5 desc2012(.I0(un4_v_high_s_1_48),.I1(un4_v_low_s_1_48),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_43[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2012.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[43:43]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2013(.I0(acs_prob_tdata_22[0:0]),.I1(acs_prob_tdata_23[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2013.INIT=16'h9669;
  LUT2 desc2014(.I0(un4_v_high_s_1_48),.I1(un4_v_low_s_1_48),.O(v_diff_1_axb_1));
defparam desc2014.INIT=4'h9;
  LUT2 desc2015(.I0(un4_v_high_s_2_48),.I1(un4_v_low_s_2_48),.O(v_diff_1_axb_2));
defparam desc2015.INIT=4'h9;
  LUT2 desc2016(.I0(un4_v_high_s_3_48),.I1(un4_v_low_s_3_48),.O(v_diff_1_axb_3));
defparam desc2016.INIT=4'h9;
  LUT2 desc2017(.I0(un4_v_high_s_4_48),.I1(un4_v_low_s_4_48),.O(v_diff_1_axb_4));
defparam desc2017.INIT=4'h9;
  LUT2 desc2018(.I0(un4_v_high_s_5_48),.I1(un4_v_low_s_5_48),.O(v_diff_1_axb_5));
defparam desc2018.INIT=4'h9;
  LUT2 desc2019(.I0(un4_v_high_s_6_48),.I1(un4_v_low_s_6_48),.O(v_diff_1_axb_6));
defparam desc2019.INIT=4'h9;
  LUT2 desc2020(.I0(un4_v_high_s_7_48),.I1(un4_v_low_s_7_48),.O(v_diff_1_axb_7));
defparam desc2020.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_22[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_22[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_22[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_22[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_22[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_22[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_22[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_23[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_23[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_23[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_23[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_23[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_23[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_23[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_23[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2021(.I0(acs_prob_tdata_22[0:0]),.I1(acs_prob_tdata_23[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1388));
defparam desc2021.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_23[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_22[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2022(.I0(un4_v_high_s_8_48),.I1(un4_v_low_s_8_48),.O(v_diff_1_axb_8));
defparam desc2022.INIT=4'h9;
  LUT6 desc2023(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2023.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI04871(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI04871.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNII6DA1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNII6DA1));
defparam s_axis_inbranch_tlast_d_RNII6DA1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_22[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIEGCC1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_48));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_48));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_23[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_48));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_23[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_48));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_23[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_48));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_23[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_48));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_23[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_48));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_23[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_48));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_23[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_23[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_48));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_48));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_22[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_48));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_22[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_48));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_22[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_48));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_22[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_48));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_22[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_48));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_22[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_48));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_22[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_22[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2024(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2025(.DI(un4_v_low_s_7_48),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2026(.DI(un4_v_low_s_6_48),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2027(.DI(un4_v_low_s_5_48),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2028(.DI(un4_v_low_s_4_48),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2029(.DI(un4_v_low_s_3_48),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2030(.DI(un4_v_low_s_2_48),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2031(.DI(un4_v_low_s_1_48),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2032(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2033(.Q(acs_prob_tdata_43[0:0]),.D(N_1388),.C(aclk),.R(s_axis_inbranch_tlast_d_RNII6DA1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2033_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2034(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIEGCC1_O6));
defparam desc2034.INIT=16'hF4F0;
  LUT2 desc2035(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2035.INIT=4'h8;
endmodule
module acsZ0_49_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_47,acs_prob_tdata_46,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_55,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,N_1756_1,aresetn,p_desc2042_p_O_FD,p_desc2043_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2072_p_O_FDRE);
input branch_tlast ;
output [55:55] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_47 ;
input [8:0] acs_prob_tdata_46 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_55 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNINL151_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIOHP31 ;
wire un4_v_high_s_7_49 ;
wire un4_v_low_s_7_49 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_49 ;
wire un4_v_low_s_8_49 ;
wire un4_v_high_s_6_49 ;
wire un4_v_low_s_6_49 ;
wire un4_v_high_s_5_49 ;
wire un4_v_low_s_5_49 ;
wire un4_v_high_s_4_49 ;
wire un4_v_low_s_4_49 ;
wire un4_v_high_s_3_49 ;
wire un4_v_low_s_3_49 ;
wire un4_v_high_s_2_49 ;
wire un4_v_low_s_2_49 ;
wire un4_v_high_s_1_49 ;
wire un4_v_low_s_1_49 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1368 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc2042_p_O_FD ;
input p_desc2043_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2072_p_O_FDRE ;
// instances
  FDR desc2036(.Q(acs_prob_tdata_55[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  FDR desc2037(.Q(acs_prob_tdata_55[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  FDR desc2038(.Q(acs_prob_tdata_55[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  FDR desc2039(.Q(acs_prob_tdata_55[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  FDR desc2040(.Q(acs_prob_tdata_55[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  FDR desc2041(.Q(acs_prob_tdata_55[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31));
  p_O_FD desc2042(.Q(acs_prob_tdata_55[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2042_p_O_FD));
  p_O_FD desc2043(.Q(acs_prob_tdata_55[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2043_p_O_FD));
  LUT6 desc2044(.I0(un4_v_high_s_7_49),.I1(un4_v_low_s_7_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOHP31),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2044.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2045(.I0(un4_v_high_s_8_49),.I1(un4_v_low_s_8_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOHP31),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2045.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2046(.I0(un4_v_high_s_6_49),.I1(un4_v_low_s_6_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2046.INIT=32'hACACFF00;
  LUT5 desc2047(.I0(un4_v_high_s_5_49),.I1(un4_v_low_s_5_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2047.INIT=32'hACACFF00;
  LUT5 desc2048(.I0(un4_v_high_s_4_49),.I1(un4_v_low_s_4_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2048.INIT=32'hACACFF00;
  LUT5 desc2049(.I0(un4_v_high_s_3_49),.I1(un4_v_low_s_3_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2049.INIT=32'hACACFF00;
  LUT5 desc2050(.I0(un4_v_high_s_2_49),.I1(un4_v_low_s_2_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2050.INIT=32'hACACFF00;
  LUT5 desc2051(.I0(un4_v_high_s_1_49),.I1(un4_v_low_s_1_49),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_55[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2051.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[55:55]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_46[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_46[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_46[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_46[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_46[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_46[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_46[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_47[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_47[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_47[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_47[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_47[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_47[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_47[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_47[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc2052(.I0(acs_prob_tdata_46[0:0]),.I1(acs_prob_tdata_47[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2052.INIT=16'h9669;
  LUT2 desc2053(.I0(un4_v_high_s_1_49),.I1(un4_v_low_s_1_49),.O(v_diff_1_axb_1));
defparam desc2053.INIT=4'h9;
  LUT2 desc2054(.I0(un4_v_high_s_2_49),.I1(un4_v_low_s_2_49),.O(v_diff_1_axb_2));
defparam desc2054.INIT=4'h9;
  LUT2 desc2055(.I0(un4_v_high_s_3_49),.I1(un4_v_low_s_3_49),.O(v_diff_1_axb_3));
defparam desc2055.INIT=4'h9;
  LUT2 desc2056(.I0(un4_v_high_s_4_49),.I1(un4_v_low_s_4_49),.O(v_diff_1_axb_4));
defparam desc2056.INIT=4'h9;
  LUT2 desc2057(.I0(un4_v_high_s_5_49),.I1(un4_v_low_s_5_49),.O(v_diff_1_axb_5));
defparam desc2057.INIT=4'h9;
  LUT2 desc2058(.I0(un4_v_high_s_6_49),.I1(un4_v_low_s_6_49),.O(v_diff_1_axb_6));
defparam desc2058.INIT=4'h9;
  LUT2 desc2059(.I0(un4_v_high_s_7_49),.I1(un4_v_low_s_7_49),.O(v_diff_1_axb_7));
defparam desc2059.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2060(.I0(acs_prob_tdata_46[0:0]),.I1(acs_prob_tdata_47[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1368));
defparam desc2060.INIT=32'h3C3C55AA;
  LUT2 desc2061(.I0(un4_v_high_s_8_49),.I1(un4_v_low_s_8_49),.O(v_diff_1_axb_8));
defparam desc2061.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_47[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_46[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc2062(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2062.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI6FK01(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI6FK01.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIOHP31_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIOHP31));
defparam s_axis_inbranch_tlast_d_RNIOHP31_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_46[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNINL151_O6),.C(aclk),.R(aresetn_i));
  XORCY desc2063(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2064(.DI(un4_v_low_s_7_49),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2065(.DI(un4_v_low_s_6_49),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2066(.DI(un4_v_low_s_5_49),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2067(.DI(un4_v_low_s_4_49),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2068(.DI(un4_v_low_s_3_49),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2069(.DI(un4_v_low_s_2_49),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2070(.DI(un4_v_low_s_1_49),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2071(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_49));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_49));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_47[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_49));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_47[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_49));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_47[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_49));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_47[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_49));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_47[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_49));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_47[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_49));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_47[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_47[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_49));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_49));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_46[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_49));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_46[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_49));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_46[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_49));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_46[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_49));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_46[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_49));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_46[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_49));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_46[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_46[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc2072(.Q(acs_prob_tdata_55[0:0]),.D(N_1368),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOHP31),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2072_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2073(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNINL151_O6));
defparam desc2073.INIT=16'hF4F0;
  LUT2 desc2074(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2074.INIT=4'h8;
endmodule
module acsZ0_50_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_27,acs_prob_tdata_26,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_13,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_2_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,write_ram_fsm_0_rep1,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2081_p_O_FD,p_desc2082_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2111_p_O_FDRE);
input branch_tlast ;
output [13:13] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_27 ;
input [8:0] acs_prob_tdata_26 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_13 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_2_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input write_ram_fsm_0_rep1 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI55B41_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNICNQA1 ;
wire un4_v_high_s_7_50 ;
wire un4_v_low_s_7_50 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_50 ;
wire un4_v_low_s_8_50 ;
wire un4_v_high_s_6_50 ;
wire un4_v_low_s_6_50 ;
wire un4_v_high_s_5_50 ;
wire un4_v_low_s_5_50 ;
wire un4_v_high_s_4_50 ;
wire un4_v_low_s_4_50 ;
wire un4_v_high_s_3_50 ;
wire un4_v_low_s_3_50 ;
wire un4_v_high_s_2_50 ;
wire un4_v_low_s_2_50 ;
wire un4_v_high_s_1_50 ;
wire un4_v_low_s_1_50 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1348 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc2081_p_O_FD ;
input p_desc2082_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2111_p_O_FDRE ;
// instances
  FDR desc2075(.Q(acs_prob_tdata_13[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  FDR desc2076(.Q(acs_prob_tdata_13[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  FDR desc2077(.Q(acs_prob_tdata_13[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  FDR desc2078(.Q(acs_prob_tdata_13[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  FDR desc2079(.Q(acs_prob_tdata_13[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  FDR desc2080(.Q(acs_prob_tdata_13[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1));
  p_O_FD desc2081(.Q(acs_prob_tdata_13[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2081_p_O_FD));
  p_O_FD desc2082(.Q(acs_prob_tdata_13[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2082_p_O_FD));
  LUT6 desc2083(.I0(un4_v_high_s_7_50),.I1(un4_v_low_s_7_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICNQA1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2083.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2084(.I0(un4_v_high_s_8_50),.I1(un4_v_low_s_8_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICNQA1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2084.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2085(.I0(un4_v_high_s_6_50),.I1(un4_v_low_s_6_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2085.INIT=32'hACACFF00;
  LUT5 desc2086(.I0(un4_v_high_s_5_50),.I1(un4_v_low_s_5_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2086.INIT=32'hACACFF00;
  LUT5 desc2087(.I0(un4_v_high_s_4_50),.I1(un4_v_low_s_4_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2087.INIT=32'hACACFF00;
  LUT5 desc2088(.I0(un4_v_high_s_3_50),.I1(un4_v_low_s_3_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2088.INIT=32'hACACFF00;
  LUT5 desc2089(.I0(un4_v_high_s_2_50),.I1(un4_v_low_s_2_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2089.INIT=32'hACACFF00;
  LUT5 desc2090(.I0(un4_v_high_s_1_50),.I1(un4_v_low_s_1_50),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_13[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2090.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[13:13]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_26[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_26[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_26[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_26[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_26[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_26[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_26[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_27[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_27[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_27[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_27[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_27[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_27[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_27[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_27[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc2091(.I0(acs_prob_tdata_26[0:0]),.I1(acs_prob_tdata_27[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2091.INIT=16'h9669;
  LUT2 desc2092(.I0(un4_v_high_s_1_50),.I1(un4_v_low_s_1_50),.O(v_diff_1_axb_1));
defparam desc2092.INIT=4'h9;
  LUT2 desc2093(.I0(un4_v_high_s_2_50),.I1(un4_v_low_s_2_50),.O(v_diff_1_axb_2));
defparam desc2093.INIT=4'h9;
  LUT2 desc2094(.I0(un4_v_high_s_3_50),.I1(un4_v_low_s_3_50),.O(v_diff_1_axb_3));
defparam desc2094.INIT=4'h9;
  LUT2 desc2095(.I0(un4_v_high_s_4_50),.I1(un4_v_low_s_4_50),.O(v_diff_1_axb_4));
defparam desc2095.INIT=4'h9;
  LUT2 desc2096(.I0(un4_v_high_s_5_50),.I1(un4_v_low_s_5_50),.O(v_diff_1_axb_5));
defparam desc2096.INIT=4'h9;
  LUT2 desc2097(.I0(un4_v_high_s_6_50),.I1(un4_v_low_s_6_50),.O(v_diff_1_axb_6));
defparam desc2097.INIT=4'h9;
  LUT2 desc2098(.I0(un4_v_high_s_7_50),.I1(un4_v_low_s_7_50),.O(v_diff_1_axb_7));
defparam desc2098.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2099(.I0(acs_prob_tdata_26[0:0]),.I1(acs_prob_tdata_27[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1348));
defparam desc2099.INIT=32'h33CC5A5A;
  LUT2 desc2100(.I0(un4_v_high_s_8_50),.I1(un4_v_low_s_8_50),.O(v_diff_1_axb_8));
defparam desc2100.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_27[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_26[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc2101(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep1),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2101.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIQKL71(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQKL71.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNICNQA1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNICNQA1));
defparam s_axis_inbranch_tlast_d_RNICNQA1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_26[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI55B41_O6),.C(aclk),.R(aresetn_i));
  XORCY desc2102(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2103(.DI(un4_v_low_s_7_50),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2104(.DI(un4_v_low_s_6_50),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2105(.DI(un4_v_low_s_5_50),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2106(.DI(un4_v_low_s_4_50),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2107(.DI(un4_v_low_s_3_50),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2108(.DI(un4_v_low_s_2_50),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2109(.DI(un4_v_low_s_1_50),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2110(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_50));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_50));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_27[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_50));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_27[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_50));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_27[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_50));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_27[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_50));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_27[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_50));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_27[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_50));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_27[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_27[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_50));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_50));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_26[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_50));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_26[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_50));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_26[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_50));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_26[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_50));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_26[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_50));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_26[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_50));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_26[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_26[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc2111(.Q(acs_prob_tdata_13[0:0]),.D(N_1348),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICNQA1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2111_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2112(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI55B41_O6));
defparam desc2112.INIT=16'hF4F0;
  LUT2 desc2113(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2113.INIT=4'h8;
endmodule
module acsZ0_51_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_26,acs_prob_tdata_27,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_45,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,N_1756_1,aresetn,p_desc2120_p_O_FD,p_desc2121_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2150_p_O_FDRE);
input branch_tlast ;
output [45:45] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_26 ;
input [8:0] acs_prob_tdata_27 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_45 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIKSBI_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIMCJU ;
wire un4_v_high_s_7_51 ;
wire un4_v_low_s_7_51 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_51 ;
wire un4_v_low_s_8_51 ;
wire un4_v_high_s_6_51 ;
wire un4_v_low_s_6_51 ;
wire un4_v_high_s_5_51 ;
wire un4_v_low_s_5_51 ;
wire un4_v_high_s_4_51 ;
wire un4_v_low_s_4_51 ;
wire un4_v_high_s_3_51 ;
wire un4_v_low_s_3_51 ;
wire un4_v_high_s_2_51 ;
wire un4_v_low_s_2_51 ;
wire un4_v_high_s_1_51 ;
wire un4_v_low_s_1_51 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire N_1328 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire GND ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire N_1 ;
input p_desc2120_p_O_FD ;
input p_desc2121_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2150_p_O_FDRE ;
// instances
  FDR desc2114(.Q(acs_prob_tdata_45[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  FDR desc2115(.Q(acs_prob_tdata_45[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  FDR desc2116(.Q(acs_prob_tdata_45[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  FDR desc2117(.Q(acs_prob_tdata_45[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  FDR desc2118(.Q(acs_prob_tdata_45[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  FDR desc2119(.Q(acs_prob_tdata_45[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU));
  p_O_FD desc2120(.Q(acs_prob_tdata_45[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2120_p_O_FD));
  p_O_FD desc2121(.Q(acs_prob_tdata_45[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2121_p_O_FD));
  LUT6 desc2122(.I0(un4_v_high_s_7_51),.I1(un4_v_low_s_7_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMCJU),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2122.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2123(.I0(un4_v_high_s_8_51),.I1(un4_v_low_s_8_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIMCJU),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2123.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2124(.I0(un4_v_high_s_6_51),.I1(un4_v_low_s_6_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2124.INIT=32'hACACFF00;
  LUT5 desc2125(.I0(un4_v_high_s_5_51),.I1(un4_v_low_s_5_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2125.INIT=32'hACACFF00;
  LUT5 desc2126(.I0(un4_v_high_s_4_51),.I1(un4_v_low_s_4_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2126.INIT=32'hACACFF00;
  LUT5 desc2127(.I0(un4_v_high_s_3_51),.I1(un4_v_low_s_3_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2127.INIT=32'hACACFF00;
  LUT5 desc2128(.I0(un4_v_high_s_2_51),.I1(un4_v_low_s_2_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2128.INIT=32'hACACFF00;
  LUT5 desc2129(.I0(un4_v_high_s_1_51),.I1(un4_v_low_s_1_51),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_45[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2129.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[45:45]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_27[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_27[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_27[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_27[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_27[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_27[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_27[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_27[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc2130(.I0(acs_prob_tdata_26[0:0]),.I1(acs_prob_tdata_27[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2130.INIT=16'h9669;
  LUT2 desc2131(.I0(un4_v_high_s_1_51),.I1(un4_v_low_s_1_51),.O(v_diff_1_axb_1));
defparam desc2131.INIT=4'h9;
  LUT2 desc2132(.I0(un4_v_high_s_2_51),.I1(un4_v_low_s_2_51),.O(v_diff_1_axb_2));
defparam desc2132.INIT=4'h9;
  LUT2 desc2133(.I0(un4_v_high_s_3_51),.I1(un4_v_low_s_3_51),.O(v_diff_1_axb_3));
defparam desc2133.INIT=4'h9;
  LUT2 desc2134(.I0(un4_v_high_s_4_51),.I1(un4_v_low_s_4_51),.O(v_diff_1_axb_4));
defparam desc2134.INIT=4'h9;
  LUT2 desc2135(.I0(un4_v_high_s_5_51),.I1(un4_v_low_s_5_51),.O(v_diff_1_axb_5));
defparam desc2135.INIT=4'h9;
  LUT2 desc2136(.I0(un4_v_high_s_6_51),.I1(un4_v_low_s_6_51),.O(v_diff_1_axb_6));
defparam desc2136.INIT=4'h9;
  LUT2 desc2137(.I0(un4_v_high_s_7_51),.I1(un4_v_low_s_7_51),.O(v_diff_1_axb_7));
defparam desc2137.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_26[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_26[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_26[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_26[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_26[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_26[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_26[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2138(.I0(acs_prob_tdata_26[0:0]),.I1(acs_prob_tdata_27[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1328));
defparam desc2138.INIT=32'h3C3C55AA;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_26[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2139(.I0(un4_v_high_s_8_51),.I1(un4_v_low_s_8_51),.O(v_diff_1_axb_8));
defparam desc2139.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_27[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT6 desc2140(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2140.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI4AER(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI4AER.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIMCJU_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIMCJU));
defparam s_axis_inbranch_tlast_d_RNIMCJU_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_26[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIKSBI_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_51));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_51));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_26[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_51));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_26[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_51));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_26[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_51));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_26[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_51));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_26[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_51));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_26[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_51));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_26[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_26[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2141(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2142(.DI(un4_v_low_s_7_51),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2143(.DI(un4_v_low_s_6_51),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2144(.DI(un4_v_low_s_5_51),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2145(.DI(un4_v_low_s_4_51),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2146(.DI(un4_v_low_s_3_51),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2147(.DI(un4_v_low_s_2_51),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2148(.DI(un4_v_low_s_1_51),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2149(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_51));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_51));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_27[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_51));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_27[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_51));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_27[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_51));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_27[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_51));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_27[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_51));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_27[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_51));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_27[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_27[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  p_O_FDRE desc2150(.Q(acs_prob_tdata_45[0:0]),.D(N_1328),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIMCJU),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2150_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2151(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIKSBI_O6));
defparam desc2151.INIT=16'hF4F0;
  LUT2 desc2152(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2152.INIT=4'h8;
endmodule
module acsZ0_52_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_61,acs_prob_tdata_60,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_30,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2159_p_O_FD,p_desc2160_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2189_p_O_FDRE);
input branch_tlast ;
output [30:30] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_61 ;
input [8:0] acs_prob_tdata_60 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_30 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI2LNG1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIAOTE1 ;
wire un4_v_high_s_7_52 ;
wire un4_v_low_s_7_52 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_52 ;
wire un4_v_low_s_8_52 ;
wire un4_v_high_s_6_52 ;
wire un4_v_low_s_6_52 ;
wire un4_v_high_s_5_52 ;
wire un4_v_low_s_5_52 ;
wire un4_v_high_s_4_52 ;
wire un4_v_low_s_4_52 ;
wire un4_v_high_s_3_52 ;
wire un4_v_low_s_3_52 ;
wire un4_v_high_s_2_52 ;
wire un4_v_low_s_2_52 ;
wire un4_v_high_s_1_52 ;
wire un4_v_low_s_1_52 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1308 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2159_p_O_FD ;
input p_desc2160_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2189_p_O_FDRE ;
// instances
  FDR desc2153(.Q(acs_prob_tdata_30[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  FDR desc2154(.Q(acs_prob_tdata_30[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  FDR desc2155(.Q(acs_prob_tdata_30[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  FDR desc2156(.Q(acs_prob_tdata_30[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  FDR desc2157(.Q(acs_prob_tdata_30[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  FDR desc2158(.Q(acs_prob_tdata_30[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1));
  p_O_FD desc2159(.Q(acs_prob_tdata_30[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2159_p_O_FD));
  p_O_FD desc2160(.Q(acs_prob_tdata_30[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2160_p_O_FD));
  LUT6 desc2161(.I0(un4_v_high_s_7_52),.I1(un4_v_low_s_7_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAOTE1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2161.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2162(.I0(un4_v_high_s_8_52),.I1(un4_v_low_s_8_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIAOTE1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2162.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2163(.I0(un4_v_high_s_6_52),.I1(un4_v_low_s_6_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2163.INIT=32'hACACFF00;
  LUT5 desc2164(.I0(un4_v_high_s_5_52),.I1(un4_v_low_s_5_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2164.INIT=32'hACACFF00;
  LUT5 desc2165(.I0(un4_v_high_s_4_52),.I1(un4_v_low_s_4_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2165.INIT=32'hACACFF00;
  LUT5 desc2166(.I0(un4_v_high_s_3_52),.I1(un4_v_low_s_3_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2166.INIT=32'hACACFF00;
  LUT5 desc2167(.I0(un4_v_high_s_2_52),.I1(un4_v_low_s_2_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2167.INIT=32'hACACFF00;
  LUT5 desc2168(.I0(un4_v_high_s_1_52),.I1(un4_v_low_s_1_52),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_30[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2168.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[30:30]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2169(.I0(acs_prob_tdata_60[0:0]),.I1(acs_prob_tdata_61[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2169.INIT=16'h9669;
  LUT2 desc2170(.I0(un4_v_high_s_1_52),.I1(un4_v_low_s_1_52),.O(v_diff_1_axb_1));
defparam desc2170.INIT=4'h9;
  LUT2 desc2171(.I0(un4_v_high_s_2_52),.I1(un4_v_low_s_2_52),.O(v_diff_1_axb_2));
defparam desc2171.INIT=4'h9;
  LUT2 desc2172(.I0(un4_v_high_s_3_52),.I1(un4_v_low_s_3_52),.O(v_diff_1_axb_3));
defparam desc2172.INIT=4'h9;
  LUT2 desc2173(.I0(un4_v_high_s_4_52),.I1(un4_v_low_s_4_52),.O(v_diff_1_axb_4));
defparam desc2173.INIT=4'h9;
  LUT2 desc2174(.I0(un4_v_high_s_5_52),.I1(un4_v_low_s_5_52),.O(v_diff_1_axb_5));
defparam desc2174.INIT=4'h9;
  LUT2 desc2175(.I0(un4_v_high_s_6_52),.I1(un4_v_low_s_6_52),.O(v_diff_1_axb_6));
defparam desc2175.INIT=4'h9;
  LUT2 desc2176(.I0(un4_v_high_s_7_52),.I1(un4_v_low_s_7_52),.O(v_diff_1_axb_7));
defparam desc2176.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_60[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_60[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_60[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_60[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_60[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_60[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_60[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_61[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_61[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_61[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_61[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_61[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_61[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_61[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_61[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2177(.I0(acs_prob_tdata_60[0:0]),.I1(acs_prob_tdata_61[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1308));
defparam desc2177.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_61[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_60[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2178(.I0(un4_v_high_s_8_52),.I1(un4_v_low_s_8_52),.O(v_diff_1_axb_8));
defparam desc2178.INIT=4'h9;
  LUT6 desc2179(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2179.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIOLOB1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIOLOB1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIAOTE1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIAOTE1));
defparam s_axis_inbranch_tlast_d_RNIAOTE1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_60[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI2LNG1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_52));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_52));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_61[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_52));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_61[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_52));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_61[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_52));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_61[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_52));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_61[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_52));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_61[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_52));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_61[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_61[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_52));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_52));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_60[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_52));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_60[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_52));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_60[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_52));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_60[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_52));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_60[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_52));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_60[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_52));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_60[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_60[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2180(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2181(.DI(un4_v_low_s_7_52),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2182(.DI(un4_v_low_s_6_52),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2183(.DI(un4_v_low_s_5_52),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2184(.DI(un4_v_low_s_4_52),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2185(.DI(un4_v_low_s_3_52),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2186(.DI(un4_v_low_s_2_52),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2187(.DI(un4_v_low_s_1_52),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2188(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2189(.Q(acs_prob_tdata_30[0:0]),.D(N_1308),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIAOTE1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2189_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2190(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI2LNG1_O6));
defparam desc2190.INIT=16'hF4F0;
  LUT2 desc2191(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2191.INIT=4'h8;
endmodule
module acsZ0_53_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_31,acs_prob_tdata_30,write_ram_fsm,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_15,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2198_p_O_FD,p_desc2199_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2228_p_O_FDRE);
input branch_tlast ;
output [15:15] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_31 ;
input [8:0] acs_prob_tdata_30 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_15 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIBHAA1_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIGT0F1 ;
wire un4_v_high_s_7_53 ;
wire un4_v_low_s_7_53 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_53 ;
wire un4_v_low_s_8_53 ;
wire un4_v_high_s_6_53 ;
wire un4_v_low_s_6_53 ;
wire un4_v_high_s_5_53 ;
wire un4_v_low_s_5_53 ;
wire un4_v_high_s_4_53 ;
wire un4_v_low_s_4_53 ;
wire un4_v_high_s_3_53 ;
wire un4_v_low_s_3_53 ;
wire un4_v_high_s_2_53 ;
wire un4_v_low_s_2_53 ;
wire un4_v_high_s_1_53 ;
wire un4_v_low_s_1_53 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1288 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2198_p_O_FD ;
input p_desc2199_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2228_p_O_FDRE ;
// instances
  FDR desc2192(.Q(acs_prob_tdata_15[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  FDR desc2193(.Q(acs_prob_tdata_15[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  FDR desc2194(.Q(acs_prob_tdata_15[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  FDR desc2195(.Q(acs_prob_tdata_15[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  FDR desc2196(.Q(acs_prob_tdata_15[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  FDR desc2197(.Q(acs_prob_tdata_15[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1));
  p_O_FD desc2198(.Q(acs_prob_tdata_15[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2198_p_O_FD));
  p_O_FD desc2199(.Q(acs_prob_tdata_15[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2199_p_O_FD));
  LUT6 desc2200(.I0(un4_v_high_s_7_53),.I1(un4_v_low_s_7_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGT0F1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2200.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2201(.I0(un4_v_high_s_8_53),.I1(un4_v_low_s_8_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIGT0F1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2201.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2202(.I0(un4_v_high_s_6_53),.I1(un4_v_low_s_6_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2202.INIT=32'hACACFF00;
  LUT5 desc2203(.I0(un4_v_high_s_5_53),.I1(un4_v_low_s_5_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2203.INIT=32'hACACFF00;
  LUT5 desc2204(.I0(un4_v_high_s_4_53),.I1(un4_v_low_s_4_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2204.INIT=32'hACACFF00;
  LUT5 desc2205(.I0(un4_v_high_s_3_53),.I1(un4_v_low_s_3_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2205.INIT=32'hACACFF00;
  LUT5 desc2206(.I0(un4_v_high_s_2_53),.I1(un4_v_low_s_2_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2206.INIT=32'hACACFF00;
  LUT5 desc2207(.I0(un4_v_high_s_1_53),.I1(un4_v_low_s_1_53),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_15[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2207.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[15:15]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2208(.I0(acs_prob_tdata_30[0:0]),.I1(acs_prob_tdata_31[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2208.INIT=16'h9669;
  LUT2 desc2209(.I0(un4_v_high_s_1_53),.I1(un4_v_low_s_1_53),.O(v_diff_1_axb_1));
defparam desc2209.INIT=4'h9;
  LUT2 desc2210(.I0(un4_v_high_s_2_53),.I1(un4_v_low_s_2_53),.O(v_diff_1_axb_2));
defparam desc2210.INIT=4'h9;
  LUT2 desc2211(.I0(un4_v_high_s_3_53),.I1(un4_v_low_s_3_53),.O(v_diff_1_axb_3));
defparam desc2211.INIT=4'h9;
  LUT2 desc2212(.I0(un4_v_high_s_4_53),.I1(un4_v_low_s_4_53),.O(v_diff_1_axb_4));
defparam desc2212.INIT=4'h9;
  LUT2 desc2213(.I0(un4_v_high_s_5_53),.I1(un4_v_low_s_5_53),.O(v_diff_1_axb_5));
defparam desc2213.INIT=4'h9;
  LUT2 desc2214(.I0(un4_v_high_s_6_53),.I1(un4_v_low_s_6_53),.O(v_diff_1_axb_6));
defparam desc2214.INIT=4'h9;
  LUT2 desc2215(.I0(un4_v_high_s_7_53),.I1(un4_v_low_s_7_53),.O(v_diff_1_axb_7));
defparam desc2215.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_30[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_30[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_30[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_30[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_30[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_30[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_30[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_31[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_31[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_31[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_31[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_31[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_31[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_31[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_31[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2216(.I0(acs_prob_tdata_30[0:0]),.I1(acs_prob_tdata_31[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1288));
defparam desc2216.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_31[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_30[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2217(.I0(un4_v_high_s_8_53),.I1(un4_v_low_s_8_53),.O(v_diff_1_axb_8));
defparam desc2217.INIT=4'h9;
  LUT6 desc2218(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2218.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIUQRB1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIUQRB1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIGT0F1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIGT0F1));
defparam s_axis_inbranch_tlast_d_RNIGT0F1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_30[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIBHAA1_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_53));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_53));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_31[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_53));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_31[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_53));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_31[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_53));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_31[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_53));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_31[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_53));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_31[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_53));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_31[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_31[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_53));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_53));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_30[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_53));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_30[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_53));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_30[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_53));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_30[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_53));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_30[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_53));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_30[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_53));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_30[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_30[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2219(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2220(.DI(un4_v_low_s_7_53),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2221(.DI(un4_v_low_s_6_53),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2222(.DI(un4_v_low_s_5_53),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2223(.DI(un4_v_low_s_4_53),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2224(.DI(un4_v_low_s_3_53),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2225(.DI(un4_v_low_s_2_53),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2226(.DI(un4_v_low_s_1_53),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2227(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2228(.Q(acs_prob_tdata_15[0:0]),.D(N_1288),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIGT0F1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2228_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2229(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIBHAA1_O6));
defparam desc2229.INIT=16'hF4F0;
  LUT2 desc2230(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2230.INIT=4'h8;
endmodule
module acsZ0_54_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_55,acs_prob_tdata_54,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_27,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_3_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2237_p_O_FD,p_desc2238_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2267_p_O_FDRE);
input branch_tlast ;
output [27:27] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_55 ;
input [8:0] acs_prob_tdata_54 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_27 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_3_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIKMV21_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIM8D81 ;
wire un4_v_high_s_7_54 ;
wire un4_v_low_s_7_54 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_54 ;
wire un4_v_low_s_8_54 ;
wire un4_v_high_s_6_54 ;
wire un4_v_low_s_6_54 ;
wire un4_v_high_s_5_54 ;
wire un4_v_low_s_5_54 ;
wire un4_v_high_s_4_54 ;
wire un4_v_low_s_4_54 ;
wire un4_v_high_s_3_54 ;
wire un4_v_low_s_3_54 ;
wire un4_v_high_s_2_54 ;
wire un4_v_low_s_2_54 ;
wire un4_v_high_s_1_54 ;
wire un4_v_low_s_1_54 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1268 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2237_p_O_FD ;
input p_desc2238_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2267_p_O_FDRE ;
// instances
  FDR desc2231(.Q(acs_prob_tdata_27[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  FDR desc2232(.Q(acs_prob_tdata_27[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  FDR desc2233(.Q(acs_prob_tdata_27[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  FDR desc2234(.Q(acs_prob_tdata_27[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  FDR desc2235(.Q(acs_prob_tdata_27[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  FDR desc2236(.Q(acs_prob_tdata_27[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81));
  p_O_FD desc2237(.Q(acs_prob_tdata_27[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2237_p_O_FD));
  p_O_FD desc2238(.Q(acs_prob_tdata_27[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2238_p_O_FD));
  LUT6 desc2239(.I0(un4_v_high_s_7_54),.I1(un4_v_low_s_7_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIM8D81),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2239.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2240(.I0(un4_v_high_s_8_54),.I1(un4_v_low_s_8_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIM8D81),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2240.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2241(.I0(un4_v_high_s_6_54),.I1(un4_v_low_s_6_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2241.INIT=32'hACACFF00;
  LUT5 desc2242(.I0(un4_v_high_s_5_54),.I1(un4_v_low_s_5_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2242.INIT=32'hACACFF00;
  LUT5 desc2243(.I0(un4_v_high_s_4_54),.I1(un4_v_low_s_4_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2243.INIT=32'hACACFF00;
  LUT5 desc2244(.I0(un4_v_high_s_3_54),.I1(un4_v_low_s_3_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2244.INIT=32'hACACFF00;
  LUT5 desc2245(.I0(un4_v_high_s_2_54),.I1(un4_v_low_s_2_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2245.INIT=32'hACACFF00;
  LUT5 desc2246(.I0(un4_v_high_s_1_54),.I1(un4_v_low_s_1_54),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_27[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2246.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[27:27]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2247(.I0(acs_prob_tdata_54[0:0]),.I1(acs_prob_tdata_55[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2247.INIT=16'h9669;
  LUT2 desc2248(.I0(un4_v_high_s_1_54),.I1(un4_v_low_s_1_54),.O(v_diff_1_axb_1));
defparam desc2248.INIT=4'h9;
  LUT2 desc2249(.I0(un4_v_high_s_2_54),.I1(un4_v_low_s_2_54),.O(v_diff_1_axb_2));
defparam desc2249.INIT=4'h9;
  LUT2 desc2250(.I0(un4_v_high_s_3_54),.I1(un4_v_low_s_3_54),.O(v_diff_1_axb_3));
defparam desc2250.INIT=4'h9;
  LUT2 desc2251(.I0(un4_v_high_s_4_54),.I1(un4_v_low_s_4_54),.O(v_diff_1_axb_4));
defparam desc2251.INIT=4'h9;
  LUT2 desc2252(.I0(un4_v_high_s_5_54),.I1(un4_v_low_s_5_54),.O(v_diff_1_axb_5));
defparam desc2252.INIT=4'h9;
  LUT2 desc2253(.I0(un4_v_high_s_6_54),.I1(un4_v_low_s_6_54),.O(v_diff_1_axb_6));
defparam desc2253.INIT=4'h9;
  LUT2 desc2254(.I0(un4_v_high_s_7_54),.I1(un4_v_low_s_7_54),.O(v_diff_1_axb_7));
defparam desc2254.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_54[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_54[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_54[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_54[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_54[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_54[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_54[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_55[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_55[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_55[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_55[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_55[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_55[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_55[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_55[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2255(.I0(acs_prob_tdata_54[0:0]),.I1(acs_prob_tdata_55[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1268));
defparam desc2255.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_55[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_54[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2256(.I0(un4_v_high_s_8_54),.I1(un4_v_low_s_8_54),.O(v_diff_1_axb_8));
defparam desc2256.INIT=4'h9;
  LUT6 desc2257(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2257.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI46851(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI46851.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIM8D81_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIM8D81));
defparam s_axis_inbranch_tlast_d_RNIM8D81_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_54[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIKMV21_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_54));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_54));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_55[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_54));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_55[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_54));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_55[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_54));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_55[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_54));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_55[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_54));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_55[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_54));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_55[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_55[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_54));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_54));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_54[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_54));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_54[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_54));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_54[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_54));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_54[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_54));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_54[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_54));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_54[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_54));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_54[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_54[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2258(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2259(.DI(un4_v_low_s_7_54),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2260(.DI(un4_v_low_s_6_54),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2261(.DI(un4_v_low_s_5_54),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2262(.DI(un4_v_low_s_4_54),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2263(.DI(un4_v_low_s_3_54),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2264(.DI(un4_v_low_s_2_54),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2265(.DI(un4_v_low_s_1_54),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2266(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2267(.Q(acs_prob_tdata_27[0:0]),.D(N_1268),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIM8D81),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2267_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2268(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIKMV21_O6));
defparam desc2268.INIT=16'hF4F0;
  LUT2 desc2269(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2269.INIT=4'h8;
endmodule
module acsZ0_55_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_55,acs_prob_tdata_54,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_59,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,N_1756_1,aresetn,p_desc2276_p_O_FD,p_desc2277_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2306_p_O_FDRE);
input branch_tlast ;
output [59:59] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_55 ;
input [8:0] acs_prob_tdata_54 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_59 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI3E0H_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNI0U5S ;
wire un4_v_high_s_7_55 ;
wire un4_v_low_s_7_55 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_55 ;
wire un4_v_low_s_8_55 ;
wire un4_v_high_s_6_55 ;
wire un4_v_low_s_6_55 ;
wire un4_v_high_s_5_55 ;
wire un4_v_low_s_5_55 ;
wire un4_v_high_s_4_55 ;
wire un4_v_low_s_4_55 ;
wire un4_v_high_s_3_55 ;
wire un4_v_low_s_3_55 ;
wire un4_v_high_s_2_55 ;
wire un4_v_low_s_2_55 ;
wire un4_v_high_s_1_55 ;
wire un4_v_low_s_1_55 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1248 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2276_p_O_FD ;
input p_desc2277_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2306_p_O_FDRE ;
// instances
  FDR desc2270(.Q(acs_prob_tdata_59[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  FDR desc2271(.Q(acs_prob_tdata_59[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  FDR desc2272(.Q(acs_prob_tdata_59[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  FDR desc2273(.Q(acs_prob_tdata_59[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  FDR desc2274(.Q(acs_prob_tdata_59[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  FDR desc2275(.Q(acs_prob_tdata_59[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S));
  p_O_FD desc2276(.Q(acs_prob_tdata_59[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2276_p_O_FD));
  p_O_FD desc2277(.Q(acs_prob_tdata_59[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2277_p_O_FD));
  LUT6 desc2278(.I0(un4_v_high_s_7_55),.I1(un4_v_low_s_7_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI0U5S),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2278.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2279(.I0(un4_v_high_s_8_55),.I1(un4_v_low_s_8_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNI0U5S),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2279.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2280(.I0(un4_v_high_s_6_55),.I1(un4_v_low_s_6_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2280.INIT=32'hACACFF00;
  LUT5 desc2281(.I0(un4_v_high_s_5_55),.I1(un4_v_low_s_5_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2281.INIT=32'hACACFF00;
  LUT5 desc2282(.I0(un4_v_high_s_4_55),.I1(un4_v_low_s_4_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2282.INIT=32'hACACFF00;
  LUT5 desc2283(.I0(un4_v_high_s_3_55),.I1(un4_v_low_s_3_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2283.INIT=32'hACACFF00;
  LUT5 desc2284(.I0(un4_v_high_s_2_55),.I1(un4_v_low_s_2_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2284.INIT=32'hACACFF00;
  LUT5 desc2285(.I0(un4_v_high_s_1_55),.I1(un4_v_low_s_1_55),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_59[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2285.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[59:59]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2286(.I0(acs_prob_tdata_54[0:0]),.I1(acs_prob_tdata_55[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2286.INIT=16'h9669;
  LUT2 desc2287(.I0(un4_v_high_s_1_55),.I1(un4_v_low_s_1_55),.O(v_diff_1_axb_1));
defparam desc2287.INIT=4'h9;
  LUT2 desc2288(.I0(un4_v_high_s_2_55),.I1(un4_v_low_s_2_55),.O(v_diff_1_axb_2));
defparam desc2288.INIT=4'h9;
  LUT2 desc2289(.I0(un4_v_high_s_3_55),.I1(un4_v_low_s_3_55),.O(v_diff_1_axb_3));
defparam desc2289.INIT=4'h9;
  LUT2 desc2290(.I0(un4_v_high_s_4_55),.I1(un4_v_low_s_4_55),.O(v_diff_1_axb_4));
defparam desc2290.INIT=4'h9;
  LUT2 desc2291(.I0(un4_v_high_s_5_55),.I1(un4_v_low_s_5_55),.O(v_diff_1_axb_5));
defparam desc2291.INIT=4'h9;
  LUT2 desc2292(.I0(un4_v_high_s_6_55),.I1(un4_v_low_s_6_55),.O(v_diff_1_axb_6));
defparam desc2292.INIT=4'h9;
  LUT2 desc2293(.I0(un4_v_high_s_7_55),.I1(un4_v_low_s_7_55),.O(v_diff_1_axb_7));
defparam desc2293.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_54[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_54[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_54[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_54[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_54[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_54[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_54[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_55[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_55[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_55[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_55[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_55[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_55[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_55[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_55[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2294(.I0(acs_prob_tdata_54[0:0]),.I1(acs_prob_tdata_55[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1248));
defparam desc2294.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_55[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_54[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2295(.I0(un4_v_high_s_8_55),.I1(un4_v_low_s_8_55),.O(v_diff_1_axb_8));
defparam desc2295.INIT=4'h9;
  LUT6 desc2296(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2296.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIER0P(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIER0P.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNI0U5S_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNI0U5S));
defparam s_axis_inbranch_tlast_d_RNI0U5S_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_54[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI3E0H_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_55));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_55));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_55[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_55));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_55[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_55));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_55[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_55));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_55[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_55));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_55[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_55));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_55[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_55));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_55[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_55[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_55));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_55));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_54[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_55));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_54[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_55));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_54[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_55));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_54[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_55));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_54[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_55));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_54[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_55));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_54[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_54[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2297(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2298(.DI(un4_v_low_s_7_55),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2299(.DI(un4_v_low_s_6_55),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2300(.DI(un4_v_low_s_5_55),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2301(.DI(un4_v_low_s_4_55),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2302(.DI(un4_v_low_s_3_55),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2303(.DI(un4_v_low_s_2_55),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2304(.DI(un4_v_low_s_1_55),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2305(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2306(.Q(acs_prob_tdata_59[0:0]),.D(N_1248),.C(aclk),.R(s_axis_inbranch_tlast_d_RNI0U5S),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2306_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2307(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI3E0H_O6));
defparam desc2307.INIT=16'hF4F0;
  LUT2 desc2308(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2308.INIT=4'h8;
endmodule
module acsZ0_56_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_25,acs_prob_tdata_24,write_ram_fsm_3,write_ram_fsm_0,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_44,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,N_1756_1,aresetn,p_desc2315_p_O_FD,p_desc2316_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2345_p_O_FDRE);
input branch_tlast ;
output [44:44] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_25 ;
input [8:0] acs_prob_tdata_24 ;
input write_ram_fsm_3 ;
input write_ram_fsm_0 ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_44 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire write_ram_fsm_3 ;
wire write_ram_fsm_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIH6CV_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIK9GC1 ;
wire un4_v_high_s_7_56 ;
wire un4_v_low_s_7_56 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_56 ;
wire un4_v_low_s_8_56 ;
wire un4_v_high_s_6_56 ;
wire un4_v_low_s_6_56 ;
wire un4_v_high_s_5_56 ;
wire un4_v_low_s_5_56 ;
wire un4_v_high_s_4_56 ;
wire un4_v_low_s_4_56 ;
wire un4_v_high_s_3_56 ;
wire un4_v_low_s_3_56 ;
wire un4_v_high_s_2_56 ;
wire un4_v_low_s_2_56 ;
wire un4_v_high_s_1_56 ;
wire un4_v_low_s_1_56 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1228 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2315_p_O_FD ;
input p_desc2316_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2345_p_O_FDRE ;
// instances
  FDR desc2309(.Q(acs_prob_tdata_44[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  FDR desc2310(.Q(acs_prob_tdata_44[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  FDR desc2311(.Q(acs_prob_tdata_44[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  FDR desc2312(.Q(acs_prob_tdata_44[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  FDR desc2313(.Q(acs_prob_tdata_44[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  FDR desc2314(.Q(acs_prob_tdata_44[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1));
  p_O_FD desc2315(.Q(acs_prob_tdata_44[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2315_p_O_FD));
  p_O_FD desc2316(.Q(acs_prob_tdata_44[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2316_p_O_FD));
  LUT6 desc2317(.I0(un4_v_high_s_7_56),.I1(un4_v_low_s_7_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK9GC1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2317.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2318(.I0(un4_v_high_s_8_56),.I1(un4_v_low_s_8_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIK9GC1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2318.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2319(.I0(un4_v_high_s_6_56),.I1(un4_v_low_s_6_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2319.INIT=32'hACACFF00;
  LUT5 desc2320(.I0(un4_v_high_s_5_56),.I1(un4_v_low_s_5_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2320.INIT=32'hACACFF00;
  LUT5 desc2321(.I0(un4_v_high_s_4_56),.I1(un4_v_low_s_4_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2321.INIT=32'hACACFF00;
  LUT5 desc2322(.I0(un4_v_high_s_3_56),.I1(un4_v_low_s_3_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2322.INIT=32'hACACFF00;
  LUT5 desc2323(.I0(un4_v_high_s_2_56),.I1(un4_v_low_s_2_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2323.INIT=32'hACACFF00;
  LUT5 desc2324(.I0(un4_v_high_s_1_56),.I1(un4_v_low_s_1_56),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_44[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2324.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[44:44]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2325(.I0(acs_prob_tdata_24[0:0]),.I1(acs_prob_tdata_25[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2325.INIT=16'h9669;
  LUT2 desc2326(.I0(un4_v_high_s_1_56),.I1(un4_v_low_s_1_56),.O(v_diff_1_axb_1));
defparam desc2326.INIT=4'h9;
  LUT2 desc2327(.I0(un4_v_high_s_2_56),.I1(un4_v_low_s_2_56),.O(v_diff_1_axb_2));
defparam desc2327.INIT=4'h9;
  LUT2 desc2328(.I0(un4_v_high_s_3_56),.I1(un4_v_low_s_3_56),.O(v_diff_1_axb_3));
defparam desc2328.INIT=4'h9;
  LUT2 desc2329(.I0(un4_v_high_s_4_56),.I1(un4_v_low_s_4_56),.O(v_diff_1_axb_4));
defparam desc2329.INIT=4'h9;
  LUT2 desc2330(.I0(un4_v_high_s_5_56),.I1(un4_v_low_s_5_56),.O(v_diff_1_axb_5));
defparam desc2330.INIT=4'h9;
  LUT2 desc2331(.I0(un4_v_high_s_6_56),.I1(un4_v_low_s_6_56),.O(v_diff_1_axb_6));
defparam desc2331.INIT=4'h9;
  LUT2 desc2332(.I0(un4_v_high_s_7_56),.I1(un4_v_low_s_7_56),.O(v_diff_1_axb_7));
defparam desc2332.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_24[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_24[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_24[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_24[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_24[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_24[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_24[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_25[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_25[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_25[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_25[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_25[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_25[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_25[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_25[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2333(.I0(acs_prob_tdata_24[0:0]),.I1(acs_prob_tdata_25[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1228));
defparam desc2333.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_25[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_24[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2334(.I0(un4_v_high_s_8_56),.I1(un4_v_low_s_8_56),.O(v_diff_1_axb_8));
defparam desc2334.INIT=4'h9;
  LUT6 desc2335(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_3),.I2(write_ram_fsm_0_rep2),.I3(write_ram_fsm_0),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2335.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI27B91(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI27B91.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIK9GC1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIK9GC1));
defparam s_axis_inbranch_tlast_d_RNIK9GC1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_24[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIH6CV_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_56));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_56));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_25[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_56));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_25[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_56));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_25[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_56));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_25[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_56));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_25[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_56));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_25[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_56));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_25[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_25[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_56));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_56));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_24[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_56));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_24[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_56));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_24[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_56));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_24[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_56));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_24[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_56));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_24[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_56));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_24[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_24[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2336(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2337(.DI(un4_v_low_s_7_56),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2338(.DI(un4_v_low_s_6_56),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2339(.DI(un4_v_low_s_5_56),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2340(.DI(un4_v_low_s_4_56),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2341(.DI(un4_v_low_s_3_56),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2342(.DI(un4_v_low_s_2_56),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2343(.DI(un4_v_low_s_1_56),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2344(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2345(.Q(acs_prob_tdata_44[0:0]),.D(N_1228),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIK9GC1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2345_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2346(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIH6CV_O6));
defparam desc2346.INIT=16'hF4F0;
  LUT2 desc2347(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2347.INIT=4'h8;
endmodule
module acsZ0_57_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_49,acs_prob_tdata_48,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_56,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep1,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,N_1756_1,aresetn,p_desc2354_p_O_FD,p_desc2355_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2384_p_O_FDRE);
input branch_tlast ;
output [56:56] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_49 ;
input [8:0] acs_prob_tdata_48 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_56 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep1 ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep1 ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIQB181_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIQKS51 ;
wire un4_v_high_s_7_57 ;
wire un4_v_low_s_7_57 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_57 ;
wire un4_v_low_s_8_57 ;
wire un4_v_high_s_6_57 ;
wire un4_v_low_s_6_57 ;
wire un4_v_high_s_5_57 ;
wire un4_v_low_s_5_57 ;
wire un4_v_high_s_4_57 ;
wire un4_v_low_s_4_57 ;
wire un4_v_high_s_3_57 ;
wire un4_v_low_s_3_57 ;
wire un4_v_high_s_2_57 ;
wire un4_v_low_s_2_57 ;
wire un4_v_high_s_1_57 ;
wire un4_v_low_s_1_57 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1208 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc2354_p_O_FD ;
input p_desc2355_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2384_p_O_FDRE ;
// instances
  FDR desc2348(.Q(acs_prob_tdata_56[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  FDR desc2349(.Q(acs_prob_tdata_56[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  FDR desc2350(.Q(acs_prob_tdata_56[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  FDR desc2351(.Q(acs_prob_tdata_56[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  FDR desc2352(.Q(acs_prob_tdata_56[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  FDR desc2353(.Q(acs_prob_tdata_56[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51));
  p_O_FD desc2354(.Q(acs_prob_tdata_56[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2354_p_O_FD));
  p_O_FD desc2355(.Q(acs_prob_tdata_56[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2355_p_O_FD));
  LUT6 desc2356(.I0(un4_v_high_s_7_57),.I1(un4_v_low_s_7_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQKS51),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2356.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2357(.I0(un4_v_high_s_8_57),.I1(un4_v_low_s_8_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQKS51),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2357.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2358(.I0(un4_v_high_s_6_57),.I1(un4_v_low_s_6_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2358.INIT=32'hACACFF00;
  LUT5 desc2359(.I0(un4_v_high_s_5_57),.I1(un4_v_low_s_5_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2359.INIT=32'hACACFF00;
  LUT5 desc2360(.I0(un4_v_high_s_4_57),.I1(un4_v_low_s_4_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2360.INIT=32'hACACFF00;
  LUT5 desc2361(.I0(un4_v_high_s_3_57),.I1(un4_v_low_s_3_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2361.INIT=32'hACACFF00;
  LUT5 desc2362(.I0(un4_v_high_s_2_57),.I1(un4_v_low_s_2_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2362.INIT=32'hACACFF00;
  LUT5 desc2363(.I0(un4_v_high_s_1_57),.I1(un4_v_low_s_1_57),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_56[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2363.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[56:56]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_48[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_48[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_48[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_48[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_48[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_48[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_48[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_49[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_49[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_49[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_49[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_49[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_49[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_49[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_49[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc2364(.I0(acs_prob_tdata_48[0:0]),.I1(acs_prob_tdata_49[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2364.INIT=16'h9669;
  LUT2 desc2365(.I0(un4_v_high_s_1_57),.I1(un4_v_low_s_1_57),.O(v_diff_1_axb_1));
defparam desc2365.INIT=4'h9;
  LUT2 desc2366(.I0(un4_v_high_s_2_57),.I1(un4_v_low_s_2_57),.O(v_diff_1_axb_2));
defparam desc2366.INIT=4'h9;
  LUT2 desc2367(.I0(un4_v_high_s_3_57),.I1(un4_v_low_s_3_57),.O(v_diff_1_axb_3));
defparam desc2367.INIT=4'h9;
  LUT2 desc2368(.I0(un4_v_high_s_4_57),.I1(un4_v_low_s_4_57),.O(v_diff_1_axb_4));
defparam desc2368.INIT=4'h9;
  LUT2 desc2369(.I0(un4_v_high_s_5_57),.I1(un4_v_low_s_5_57),.O(v_diff_1_axb_5));
defparam desc2369.INIT=4'h9;
  LUT2 desc2370(.I0(un4_v_high_s_6_57),.I1(un4_v_low_s_6_57),.O(v_diff_1_axb_6));
defparam desc2370.INIT=4'h9;
  LUT2 desc2371(.I0(un4_v_high_s_7_57),.I1(un4_v_low_s_7_57),.O(v_diff_1_axb_7));
defparam desc2371.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2372(.I0(acs_prob_tdata_48[0:0]),.I1(acs_prob_tdata_49[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1208));
defparam desc2372.INIT=32'h3C3C55AA;
  LUT2 desc2373(.I0(un4_v_high_s_8_57),.I1(un4_v_low_s_8_57),.O(v_diff_1_axb_8));
defparam desc2373.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_49[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_48[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc2374(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2374.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI8IN21(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI8IN21.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIQKS51_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIQKS51));
defparam s_axis_inbranch_tlast_d_RNIQKS51_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_48[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIQB181_O6),.C(aclk),.R(aresetn_i));
  XORCY desc2375(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2376(.DI(un4_v_low_s_7_57),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2377(.DI(un4_v_low_s_6_57),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2378(.DI(un4_v_low_s_5_57),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2379(.DI(un4_v_low_s_4_57),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2380(.DI(un4_v_low_s_3_57),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2381(.DI(un4_v_low_s_2_57),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2382(.DI(un4_v_low_s_1_57),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2383(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_57));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_57));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_49[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_57));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_49[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_57));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_49[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_57));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_49[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_57));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_49[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_57));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_49[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_57));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_49[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_49[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_57));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_57));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_48[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_57));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_48[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_57));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_48[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_57));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_48[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_57));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_48[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_57));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_48[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_57));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_48[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_48[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc2384(.Q(acs_prob_tdata_56[0:0]),.D(N_1208),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQKS51),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2384_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2385(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIQB181_O6));
defparam desc2385.INIT=16'hF4F0;
  LUT2 desc2386(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2386.INIT=4'h8;
endmodule
module acsZ0_58_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_29,acs_prob_tdata_28,write_ram_fsm,branch_tvalid,branch_tdata_0_fast,acs_prob_tdata_14,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_3_0_rep1,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2393_p_O_FD,p_desc2394_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2423_p_O_FDRE);
input branch_tlast ;
output [14:14] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_29 ;
input [8:0] acs_prob_tdata_28 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_0_fast ;
output [8:0] acs_prob_tdata_14 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_3_0_rep1 ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_3_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI8RA71_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIEQTC1 ;
wire un4_v_high_s_7_58 ;
wire un4_v_low_s_7_58 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_58 ;
wire un4_v_low_s_8_58 ;
wire un4_v_high_s_6_58 ;
wire un4_v_low_s_6_58 ;
wire un4_v_high_s_5_58 ;
wire un4_v_low_s_5_58 ;
wire un4_v_high_s_4_58 ;
wire un4_v_low_s_4_58 ;
wire un4_v_high_s_3_58 ;
wire un4_v_low_s_3_58 ;
wire un4_v_high_s_2_58 ;
wire un4_v_low_s_2_58 ;
wire un4_v_high_s_1_58 ;
wire un4_v_low_s_1_58 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire N_1188 ;
wire v_diff_1_axb_8 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire un4_v_low_axb_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire N_1 ;
input p_desc2393_p_O_FD ;
input p_desc2394_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2423_p_O_FDRE ;
// instances
  FDR desc2387(.Q(acs_prob_tdata_14[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  FDR desc2388(.Q(acs_prob_tdata_14[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  FDR desc2389(.Q(acs_prob_tdata_14[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  FDR desc2390(.Q(acs_prob_tdata_14[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  FDR desc2391(.Q(acs_prob_tdata_14[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  FDR desc2392(.Q(acs_prob_tdata_14[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1));
  p_O_FD desc2393(.Q(acs_prob_tdata_14[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2393_p_O_FD));
  p_O_FD desc2394(.Q(acs_prob_tdata_14[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2394_p_O_FD));
  LUT6 desc2395(.I0(un4_v_high_s_7_58),.I1(un4_v_low_s_7_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIEQTC1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2395.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2396(.I0(un4_v_high_s_8_58),.I1(un4_v_low_s_8_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIEQTC1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2396.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2397(.I0(un4_v_high_s_6_58),.I1(un4_v_low_s_6_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2397.INIT=32'hACACFF00;
  LUT5 desc2398(.I0(un4_v_high_s_5_58),.I1(un4_v_low_s_5_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2398.INIT=32'hACACFF00;
  LUT5 desc2399(.I0(un4_v_high_s_4_58),.I1(un4_v_low_s_4_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2399.INIT=32'hACACFF00;
  LUT5 desc2400(.I0(un4_v_high_s_3_58),.I1(un4_v_low_s_3_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2400.INIT=32'hACACFF00;
  LUT5 desc2401(.I0(un4_v_high_s_2_58),.I1(un4_v_low_s_2_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2401.INIT=32'hACACFF00;
  LUT5 desc2402(.I0(un4_v_high_s_1_58),.I1(un4_v_low_s_1_58),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_14[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2402.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[14:14]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_28[1:1]),.I1(branch_tdata_0_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_28[2:2]),.I1(branch_tdata_0_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_28[3:3]),.I1(branch_tdata_0_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_28[4:4]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_28[5:5]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_28[6:6]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_28[7:7]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_29[0:0]),.I1(branch_tdata_3_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_29[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_29[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_29[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_29[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_29[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_29[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_29[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  LUT4 desc2403(.I0(acs_prob_tdata_28[0:0]),.I1(acs_prob_tdata_29[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2403.INIT=16'h9669;
  LUT2 desc2404(.I0(un4_v_high_s_1_58),.I1(un4_v_low_s_1_58),.O(v_diff_1_axb_1));
defparam desc2404.INIT=4'h9;
  LUT2 desc2405(.I0(un4_v_high_s_2_58),.I1(un4_v_low_s_2_58),.O(v_diff_1_axb_2));
defparam desc2405.INIT=4'h9;
  LUT2 desc2406(.I0(un4_v_high_s_3_58),.I1(un4_v_low_s_3_58),.O(v_diff_1_axb_3));
defparam desc2406.INIT=4'h9;
  LUT2 desc2407(.I0(un4_v_high_s_4_58),.I1(un4_v_low_s_4_58),.O(v_diff_1_axb_4));
defparam desc2407.INIT=4'h9;
  LUT2 desc2408(.I0(un4_v_high_s_5_58),.I1(un4_v_low_s_5_58),.O(v_diff_1_axb_5));
defparam desc2408.INIT=4'h9;
  LUT2 desc2409(.I0(un4_v_high_s_6_58),.I1(un4_v_low_s_6_58),.O(v_diff_1_axb_6));
defparam desc2409.INIT=4'h9;
  LUT2 desc2410(.I0(un4_v_high_s_7_58),.I1(un4_v_low_s_7_58),.O(v_diff_1_axb_7));
defparam desc2410.INIT=4'h9;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2411(.I0(acs_prob_tdata_28[0:0]),.I1(acs_prob_tdata_29[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1188));
defparam desc2411.INIT=32'h33CC5A5A;
  LUT2 desc2412(.I0(un4_v_high_s_8_58),.I1(un4_v_low_s_8_58),.O(v_diff_1_axb_8));
defparam desc2412.INIT=4'h9;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_29[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_28[8:8]),.I1(branch_tdata_0_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT6 desc2413(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2413.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNISNO91(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNISNO91.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIEQTC1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIEQTC1));
defparam s_axis_inbranch_tlast_d_RNIEQTC1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_28[0:0]),.I1(branch_tdata_0_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI8RA71_O6),.C(aclk),.R(aresetn_i));
  XORCY desc2414(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2415(.DI(un4_v_low_s_7_58),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2416(.DI(un4_v_low_s_6_58),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2417(.DI(un4_v_low_s_5_58),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2418(.DI(un4_v_low_s_4_58),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2419(.DI(un4_v_low_s_3_58),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2420(.DI(un4_v_low_s_2_58),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2421(.DI(un4_v_low_s_1_58),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2422(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_58));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_58));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_29[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_58));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_29[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_58));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_29[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_58));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_29[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_58));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_29[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_58));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_29[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_58));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_29[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_29[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_58));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_58));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_28[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_58));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_28[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_58));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_28[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_58));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_28[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_58));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_28[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_58));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_28[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_58));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_28[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_28[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  p_O_FDRE desc2423(.Q(acs_prob_tdata_14[0:0]),.D(N_1188),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIEQTC1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2423_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2424(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI8RA71_O6));
defparam desc2424.INIT=16'hF4F0;
  LUT2 desc2425(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2425.INIT=4'h8;
endmodule
module acsZ0_59_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_63,acs_prob_tdata_62,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_31,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2432_p_O_FD,p_desc2433_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2462_p_O_FDRE);
input branch_tlast ;
output [31:31] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_63 ;
input [8:0] acs_prob_tdata_62 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_31 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNI5BN31_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNICR0H1 ;
wire un4_v_high_s_7_59 ;
wire un4_v_low_s_7_59 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_59 ;
wire un4_v_low_s_8_59 ;
wire un4_v_high_s_6_59 ;
wire un4_v_low_s_6_59 ;
wire un4_v_high_s_5_59 ;
wire un4_v_low_s_5_59 ;
wire un4_v_high_s_4_59 ;
wire un4_v_low_s_4_59 ;
wire un4_v_high_s_3_59 ;
wire un4_v_low_s_3_59 ;
wire un4_v_high_s_2_59 ;
wire un4_v_low_s_2_59 ;
wire un4_v_high_s_1_59 ;
wire un4_v_low_s_1_59 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1168 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2432_p_O_FD ;
input p_desc2433_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2462_p_O_FDRE ;
// instances
  FDR desc2426(.Q(acs_prob_tdata_31[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  FDR desc2427(.Q(acs_prob_tdata_31[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  FDR desc2428(.Q(acs_prob_tdata_31[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  FDR desc2429(.Q(acs_prob_tdata_31[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  FDR desc2430(.Q(acs_prob_tdata_31[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  FDR desc2431(.Q(acs_prob_tdata_31[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1));
  p_O_FD desc2432(.Q(acs_prob_tdata_31[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2432_p_O_FD));
  p_O_FD desc2433(.Q(acs_prob_tdata_31[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2433_p_O_FD));
  LUT6 desc2434(.I0(un4_v_high_s_7_59),.I1(un4_v_low_s_7_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICR0H1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2434.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2435(.I0(un4_v_high_s_8_59),.I1(un4_v_low_s_8_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNICR0H1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2435.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2436(.I0(un4_v_high_s_6_59),.I1(un4_v_low_s_6_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2436.INIT=32'hACACFF00;
  LUT5 desc2437(.I0(un4_v_high_s_5_59),.I1(un4_v_low_s_5_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2437.INIT=32'hACACFF00;
  LUT5 desc2438(.I0(un4_v_high_s_4_59),.I1(un4_v_low_s_4_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2438.INIT=32'hACACFF00;
  LUT5 desc2439(.I0(un4_v_high_s_3_59),.I1(un4_v_low_s_3_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2439.INIT=32'hACACFF00;
  LUT5 desc2440(.I0(un4_v_high_s_2_59),.I1(un4_v_low_s_2_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2440.INIT=32'hACACFF00;
  LUT5 desc2441(.I0(un4_v_high_s_1_59),.I1(un4_v_low_s_1_59),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_31[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2441.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[31:31]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2442(.I0(acs_prob_tdata_62[0:0]),.I1(acs_prob_tdata_63[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2442.INIT=16'h9669;
  LUT2 desc2443(.I0(un4_v_high_s_1_59),.I1(un4_v_low_s_1_59),.O(v_diff_1_axb_1));
defparam desc2443.INIT=4'h9;
  LUT2 desc2444(.I0(un4_v_high_s_2_59),.I1(un4_v_low_s_2_59),.O(v_diff_1_axb_2));
defparam desc2444.INIT=4'h9;
  LUT2 desc2445(.I0(un4_v_high_s_3_59),.I1(un4_v_low_s_3_59),.O(v_diff_1_axb_3));
defparam desc2445.INIT=4'h9;
  LUT2 desc2446(.I0(un4_v_high_s_4_59),.I1(un4_v_low_s_4_59),.O(v_diff_1_axb_4));
defparam desc2446.INIT=4'h9;
  LUT2 desc2447(.I0(un4_v_high_s_5_59),.I1(un4_v_low_s_5_59),.O(v_diff_1_axb_5));
defparam desc2447.INIT=4'h9;
  LUT2 desc2448(.I0(un4_v_high_s_6_59),.I1(un4_v_low_s_6_59),.O(v_diff_1_axb_6));
defparam desc2448.INIT=4'h9;
  LUT2 desc2449(.I0(un4_v_high_s_7_59),.I1(un4_v_low_s_7_59),.O(v_diff_1_axb_7));
defparam desc2449.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_62[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_62[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_62[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_62[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_62[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_62[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_62[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_63[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_63[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_63[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_63[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_63[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_63[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_63[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_63[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2450(.I0(acs_prob_tdata_62[0:0]),.I1(acs_prob_tdata_63[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1168));
defparam desc2450.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_63[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_62[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2451(.I0(un4_v_high_s_8_59),.I1(un4_v_low_s_8_59),.O(v_diff_1_axb_8));
defparam desc2451.INIT=4'h9;
  LUT6 desc2452(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2452.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIQORD1(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIQORD1.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNICR0H1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNICR0H1));
defparam s_axis_inbranch_tlast_d_RNICR0H1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_62[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNI5BN31_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_59));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_59));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_63[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_59));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_63[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_59));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_63[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_59));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_63[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_59));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_63[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_59));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_63[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_59));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_63[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_63[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_59));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_59));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_62[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_59));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_62[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_59));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_62[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_59));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_62[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_59));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_62[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_59));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_62[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_59));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_62[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_62[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2453(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2454(.DI(un4_v_low_s_7_59),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2455(.DI(un4_v_low_s_6_59),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2456(.DI(un4_v_low_s_5_59),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2457(.DI(un4_v_low_s_4_59),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2458(.DI(un4_v_low_s_3_59),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2459(.DI(un4_v_low_s_2_59),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2460(.DI(un4_v_low_s_1_59),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2461(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2462(.Q(acs_prob_tdata_31[0:0]),.D(N_1168),.C(aclk),.R(s_axis_inbranch_tlast_d_RNICR0H1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2462_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2463(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNI5BN31_O6));
defparam desc2463.INIT=16'hF4F0;
  LUT2 desc2464(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2464.INIT=4'h8;
endmodule
module acsZ0_60_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_57,acs_prob_tdata_56,write_ram_fsm,branch_tvalid,branch_tdata_2_fast,acs_prob_tdata_28,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_1_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2471_p_O_FD,p_desc2472_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2501_p_O_FDRE);
input branch_tlast ;
output [28:28] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_57 ;
input [8:0] acs_prob_tdata_56 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_2_fast ;
output [8:0] acs_prob_tdata_28 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_1_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_1_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNINCV51_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIOBGA1 ;
wire un4_v_high_s_7_60 ;
wire un4_v_low_s_7_60 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_60 ;
wire un4_v_low_s_8_60 ;
wire un4_v_high_s_6_60 ;
wire un4_v_low_s_6_60 ;
wire un4_v_high_s_5_60 ;
wire un4_v_low_s_5_60 ;
wire un4_v_high_s_4_60 ;
wire un4_v_low_s_4_60 ;
wire un4_v_high_s_3_60 ;
wire un4_v_low_s_3_60 ;
wire un4_v_high_s_2_60 ;
wire un4_v_low_s_2_60 ;
wire un4_v_high_s_1_60 ;
wire un4_v_low_s_1_60 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1148 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2471_p_O_FD ;
input p_desc2472_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2501_p_O_FDRE ;
// instances
  FDR desc2465(.Q(acs_prob_tdata_28[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  FDR desc2466(.Q(acs_prob_tdata_28[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  FDR desc2467(.Q(acs_prob_tdata_28[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  FDR desc2468(.Q(acs_prob_tdata_28[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  FDR desc2469(.Q(acs_prob_tdata_28[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  FDR desc2470(.Q(acs_prob_tdata_28[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1));
  p_O_FD desc2471(.Q(acs_prob_tdata_28[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2471_p_O_FD));
  p_O_FD desc2472(.Q(acs_prob_tdata_28[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2472_p_O_FD));
  LUT6 desc2473(.I0(un4_v_high_s_7_60),.I1(un4_v_low_s_7_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOBGA1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2473.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2474(.I0(un4_v_high_s_8_60),.I1(un4_v_low_s_8_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIOBGA1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2474.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2475(.I0(un4_v_high_s_6_60),.I1(un4_v_low_s_6_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2475.INIT=32'hACACFF00;
  LUT5 desc2476(.I0(un4_v_high_s_5_60),.I1(un4_v_low_s_5_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2476.INIT=32'hACACFF00;
  LUT5 desc2477(.I0(un4_v_high_s_4_60),.I1(un4_v_low_s_4_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2477.INIT=32'hACACFF00;
  LUT5 desc2478(.I0(un4_v_high_s_3_60),.I1(un4_v_low_s_3_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2478.INIT=32'hACACFF00;
  LUT5 desc2479(.I0(un4_v_high_s_2_60),.I1(un4_v_low_s_2_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2479.INIT=32'hACACFF00;
  LUT5 desc2480(.I0(un4_v_high_s_1_60),.I1(un4_v_low_s_1_60),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_28[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2480.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[28:28]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2481(.I0(acs_prob_tdata_56[0:0]),.I1(acs_prob_tdata_57[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2481.INIT=16'h9669;
  LUT2 desc2482(.I0(un4_v_high_s_1_60),.I1(un4_v_low_s_1_60),.O(v_diff_1_axb_1));
defparam desc2482.INIT=4'h9;
  LUT2 desc2483(.I0(un4_v_high_s_2_60),.I1(un4_v_low_s_2_60),.O(v_diff_1_axb_2));
defparam desc2483.INIT=4'h9;
  LUT2 desc2484(.I0(un4_v_high_s_3_60),.I1(un4_v_low_s_3_60),.O(v_diff_1_axb_3));
defparam desc2484.INIT=4'h9;
  LUT2 desc2485(.I0(un4_v_high_s_4_60),.I1(un4_v_low_s_4_60),.O(v_diff_1_axb_4));
defparam desc2485.INIT=4'h9;
  LUT2 desc2486(.I0(un4_v_high_s_5_60),.I1(un4_v_low_s_5_60),.O(v_diff_1_axb_5));
defparam desc2486.INIT=4'h9;
  LUT2 desc2487(.I0(un4_v_high_s_6_60),.I1(un4_v_low_s_6_60),.O(v_diff_1_axb_6));
defparam desc2487.INIT=4'h9;
  LUT2 desc2488(.I0(un4_v_high_s_7_60),.I1(un4_v_low_s_7_60),.O(v_diff_1_axb_7));
defparam desc2488.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_56[1:1]),.I1(branch_tdata_2_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_56[2:2]),.I1(branch_tdata_2_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_56[3:3]),.I1(branch_tdata_2_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_56[4:4]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_56[5:5]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_56[6:6]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_56[7:7]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_57[0:0]),.I1(branch_tdata_1_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_57[1:1]),.I1(branch_tdata_1_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_57[2:2]),.I1(branch_tdata_1_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_57[3:3]),.I1(branch_tdata_1_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_57[4:4]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_57[5:5]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_57[6:6]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_57[7:7]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2489(.I0(acs_prob_tdata_56[0:0]),.I1(acs_prob_tdata_57[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1148));
defparam desc2489.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_57[8:8]),.I1(branch_tdata_1_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_56[8:8]),.I1(branch_tdata_2_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2490(.I0(un4_v_high_s_8_60),.I1(un4_v_low_s_8_60),.O(v_diff_1_axb_8));
defparam desc2490.INIT=4'h9;
  LUT6 desc2491(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2491.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI69B71(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI69B71.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIOBGA1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIOBGA1));
defparam s_axis_inbranch_tlast_d_RNIOBGA1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_56[0:0]),.I1(branch_tdata_2_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNINCV51_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_60));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_60));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_57[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_60));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_57[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_60));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_57[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_60));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_57[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_60));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_57[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_60));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_57[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_60));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_57[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_57[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_60));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_60));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_56[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_60));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_56[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_60));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_56[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_60));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_56[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_60));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_56[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_60));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_56[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_60));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_56[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_56[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2492(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2493(.DI(un4_v_low_s_7_60),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2494(.DI(un4_v_low_s_6_60),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2495(.DI(un4_v_low_s_5_60),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2496(.DI(un4_v_low_s_4_60),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2497(.DI(un4_v_low_s_3_60),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2498(.DI(un4_v_low_s_2_60),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2499(.DI(un4_v_low_s_1_60),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2500(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2501(.Q(acs_prob_tdata_28[0:0]),.D(N_1148),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIOBGA1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2501_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2502(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNINCV51_O6));
defparam desc2502.INIT=16'hF4F0;
  LUT2 desc2503(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2503.INIT=4'h8;
endmodule
module acsZ0_61_inj (branch_tlast,acs_dec_tdata,branch_tdata_0_1,branch_tdata_0_2,branch_tdata_0_3,branch_tdata_0_5,branch_tdata_0_0,branch_tdata_3,acs_prob_tdata_59,acs_prob_tdata_58,write_ram_fsm,branch_tvalid,branch_tdata_3_fast,acs_prob_tdata_29,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_0_0_rep2,branch_tdata_3_0_rep2,branch_tdata_0_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep2,N_1756_1,aresetn,p_desc2510_p_O_FD,p_desc2511_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2540_p_O_FDRE);
input branch_tlast ;
output [29:29] acs_dec_tdata ;
input branch_tdata_0_1 ;
input branch_tdata_0_2 ;
input branch_tdata_0_3 ;
input branch_tdata_0_5 ;
input branch_tdata_0_0 ;
input [5:0] branch_tdata_3 ;
input [8:0] acs_prob_tdata_59 ;
input [8:0] acs_prob_tdata_58 ;
input [1:1] write_ram_fsm ;
input branch_tvalid ;
input branch_tdata_3_fast ;
output [8:0] acs_prob_tdata_29 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_0_0_rep2 ;
input branch_tdata_3_0_rep2 ;
input branch_tdata_0_0_rep1 ;
input write_ram_fsm_0_rep2 ;
input write_ram_fsm_4_rep2 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_0_1 ;
wire branch_tdata_0_2 ;
wire branch_tdata_0_3 ;
wire branch_tdata_0_5 ;
wire branch_tdata_0_0 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_0_0_rep2 ;
wire branch_tdata_3_0_rep2 ;
wire branch_tdata_0_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep2 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIQ2V81_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIQEJC1 ;
wire un4_v_high_s_7_61 ;
wire un4_v_low_s_7_61 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_61 ;
wire un4_v_low_s_8_61 ;
wire un4_v_high_s_6_61 ;
wire un4_v_low_s_6_61 ;
wire un4_v_high_s_5_61 ;
wire un4_v_low_s_5_61 ;
wire un4_v_high_s_4_61 ;
wire un4_v_low_s_4_61 ;
wire un4_v_high_s_3_61 ;
wire un4_v_low_s_3_61 ;
wire un4_v_high_s_2_61 ;
wire un4_v_low_s_2_61 ;
wire un4_v_high_s_1_61 ;
wire un4_v_low_s_1_61 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1128 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2510_p_O_FD ;
input p_desc2511_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2540_p_O_FDRE ;
// instances
  FDR desc2504(.Q(acs_prob_tdata_29[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  FDR desc2505(.Q(acs_prob_tdata_29[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  FDR desc2506(.Q(acs_prob_tdata_29[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  FDR desc2507(.Q(acs_prob_tdata_29[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  FDR desc2508(.Q(acs_prob_tdata_29[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  FDR desc2509(.Q(acs_prob_tdata_29[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1));
  p_O_FD desc2510(.Q(acs_prob_tdata_29[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2510_p_O_FD));
  p_O_FD desc2511(.Q(acs_prob_tdata_29[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2511_p_O_FD));
  LUT6 desc2512(.I0(un4_v_high_s_7_61),.I1(un4_v_low_s_7_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQEJC1),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2512.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2513(.I0(un4_v_high_s_8_61),.I1(un4_v_low_s_8_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIQEJC1),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2513.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2514(.I0(un4_v_high_s_6_61),.I1(un4_v_low_s_6_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2514.INIT=32'hACACFF00;
  LUT5 desc2515(.I0(un4_v_high_s_5_61),.I1(un4_v_low_s_5_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2515.INIT=32'hACACFF00;
  LUT5 desc2516(.I0(un4_v_high_s_4_61),.I1(un4_v_low_s_4_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2516.INIT=32'hACACFF00;
  LUT5 desc2517(.I0(un4_v_high_s_3_61),.I1(un4_v_low_s_3_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2517.INIT=32'hACACFF00;
  LUT5 desc2518(.I0(un4_v_high_s_2_61),.I1(un4_v_low_s_2_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2518.INIT=32'hACACFF00;
  LUT5 desc2519(.I0(un4_v_high_s_1_61),.I1(un4_v_low_s_1_61),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_29[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2519.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[29:29]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2520(.I0(acs_prob_tdata_58[0:0]),.I1(acs_prob_tdata_59[0:0]),.I2(branch_tdata_0_0_rep2),.I3(branch_tdata_3_0_rep2),.O(v_diff_1_axb_0));
defparam desc2520.INIT=16'h9669;
  LUT2 desc2521(.I0(un4_v_high_s_1_61),.I1(un4_v_low_s_1_61),.O(v_diff_1_axb_1));
defparam desc2521.INIT=4'h9;
  LUT2 desc2522(.I0(un4_v_high_s_2_61),.I1(un4_v_low_s_2_61),.O(v_diff_1_axb_2));
defparam desc2522.INIT=4'h9;
  LUT2 desc2523(.I0(un4_v_high_s_3_61),.I1(un4_v_low_s_3_61),.O(v_diff_1_axb_3));
defparam desc2523.INIT=4'h9;
  LUT2 desc2524(.I0(un4_v_high_s_4_61),.I1(un4_v_low_s_4_61),.O(v_diff_1_axb_4));
defparam desc2524.INIT=4'h9;
  LUT2 desc2525(.I0(un4_v_high_s_5_61),.I1(un4_v_low_s_5_61),.O(v_diff_1_axb_5));
defparam desc2525.INIT=4'h9;
  LUT2 desc2526(.I0(un4_v_high_s_6_61),.I1(un4_v_low_s_6_61),.O(v_diff_1_axb_6));
defparam desc2526.INIT=4'h9;
  LUT2 desc2527(.I0(un4_v_high_s_7_61),.I1(un4_v_low_s_7_61),.O(v_diff_1_axb_7));
defparam desc2527.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_58[1:1]),.I1(branch_tdata_3[1:1]),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_58[2:2]),.I1(branch_tdata_3[2:2]),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_58[3:3]),.I1(branch_tdata_3[3:3]),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_58[4:4]),.I1(branch_tdata_3[4:4]),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_58[5:5]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_58[6:6]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_58[7:7]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_59[0:0]),.I1(branch_tdata_0_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_59[1:1]),.I1(branch_tdata_0_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_59[2:2]),.I1(branch_tdata_0_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_59[3:3]),.I1(branch_tdata_0_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_59[4:4]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_59[5:5]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_59[6:6]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_59[7:7]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2528(.I0(acs_prob_tdata_58[0:0]),.I1(acs_prob_tdata_59[0:0]),.I2(branch_tdata_0_0),.I3(branch_tdata_3[0:0]),.I4(v_diff_1[8:8]),.LO(N_1128));
defparam desc2528.INIT=32'h3C3C55AA;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_59[8:8]),.I1(branch_tdata_0_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_58[8:8]),.I1(branch_tdata_3[5:5]),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2529(.I0(un4_v_high_s_8_61),.I1(un4_v_low_s_8_61),.O(v_diff_1_axb_8));
defparam desc2529.INIT=4'h9;
  LUT6 desc2530(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_0_rep2),.I2(write_ram_fsm_4_rep2),.I3(write_ram_fsm[1:1]),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2530.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNI8CE91(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNI8CE91.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIQEJC1_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIQEJC1));
defparam s_axis_inbranch_tlast_d_RNIQEJC1_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_58[0:0]),.I1(branch_tdata_3_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIQ2V81_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_61));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_61));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_59[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_61));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_59[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_61));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_59[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_61));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_59[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_61));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_59[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_61));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_59[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_61));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_59[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_59[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_61));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_61));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_58[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_61));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_58[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_61));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_58[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_61));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_58[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_61));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_58[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_61));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_58[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_61));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_58[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_58[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2531(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2532(.DI(un4_v_low_s_7_61),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2533(.DI(un4_v_low_s_6_61),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2534(.DI(un4_v_low_s_5_61),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2535(.DI(un4_v_low_s_4_61),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2536(.DI(un4_v_low_s_3_61),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2537(.DI(un4_v_low_s_2_61),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2538(.DI(un4_v_low_s_1_61),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2539(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2540(.Q(acs_prob_tdata_29[0:0]),.D(N_1128),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIQEJC1),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2540_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2541(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIQ2V81_O6));
defparam desc2541.INIT=16'hF4F0;
  LUT2 desc2542(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2542.INIT=4'h8;
endmodule
module acsZ0_62_inj (branch_tlast,acs_dec_tdata,branch_tdata_1_1,branch_tdata_1_2,branch_tdata_1_3,branch_tdata_1_5,branch_tdata_1_0,branch_tdata_2_1,branch_tdata_2_2,branch_tdata_2_3,branch_tdata_2_5,branch_tdata_2_0,acs_prob_tdata_57,acs_prob_tdata_56,write_ram_fsm_4,write_ram_fsm_0,write_ram_fsm_1,branch_tvalid,branch_tdata_1_fast,acs_prob_tdata_60,un27_s_axis_input_tready_int,aclk,aresetn_i,branch_tdata_1_0_rep2,branch_tdata_2_0_rep2,branch_tdata_2_0_rep1,N_1756_1,aresetn,p_desc2549_p_O_FD,p_desc2550_p_O_FD,p_m_axis_outdec_tdata_Z_p_O_FDRE,p_desc2579_p_O_FDRE);
input branch_tlast ;
output [60:60] acs_dec_tdata ;
input branch_tdata_1_1 ;
input branch_tdata_1_2 ;
input branch_tdata_1_3 ;
input branch_tdata_1_5 ;
input branch_tdata_1_0 ;
input branch_tdata_2_1 ;
input branch_tdata_2_2 ;
input branch_tdata_2_3 ;
input branch_tdata_2_5 ;
input branch_tdata_2_0 ;
input [8:0] acs_prob_tdata_57 ;
input [8:0] acs_prob_tdata_56 ;
input write_ram_fsm_4 ;
input write_ram_fsm_0 ;
input write_ram_fsm_1 ;
input branch_tvalid ;
input branch_tdata_1_fast ;
output [8:0] acs_prob_tdata_60 ;
input un27_s_axis_input_tready_int ;
input aclk ;
input aresetn_i ;
input branch_tdata_1_0_rep2 ;
input branch_tdata_2_0_rep2 ;
input branch_tdata_2_0_rep1 ;
input N_1756_1 ;
input aresetn ;
wire branch_tdata_1_1 ;
wire branch_tdata_1_2 ;
wire branch_tdata_1_3 ;
wire branch_tdata_1_5 ;
wire branch_tdata_1_0 ;
wire branch_tdata_2_1 ;
wire branch_tdata_2_2 ;
wire branch_tdata_2_3 ;
wire branch_tdata_2_5 ;
wire branch_tdata_2_0 ;
wire write_ram_fsm_4 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_1 ;
wire un27_s_axis_input_tready_int ;
wire aclk ;
wire aresetn_i ;
wire branch_tdata_1_0_rep2 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_2_0_rep1 ;
wire N_1756_1 ;
wire aresetn ;
wire [6:1] m_axis_outprob_tdata_8_0 ;
wire [8:7] m_axis_outprob_tdata_8_0_e ;
wire [8:8] v_diff_1 ;
wire s_axis_inbranch_tlast_d ;
wire m_axis_outdec_tvalid_int ;
wire un1_s_axis_inbranch_tvalid ;
wire VCC ;
wire un1_s_axis_inbranch_tvalid_RNIB0PO_O6 ;
wire s_axis_inbranch_tlast_d_0 ;
wire s_axis_inbranch_tlast_d_RNIG7GU ;
wire un4_v_high_s_7_62 ;
wire un4_v_low_s_7_62 ;
wire s_axis_inbranch_tlast_d_1_sqmuxa_i ;
wire un4_v_high_s_8_62 ;
wire un4_v_low_s_8_62 ;
wire un4_v_high_s_6_62 ;
wire un4_v_low_s_6_62 ;
wire un4_v_high_s_5_62 ;
wire un4_v_low_s_5_62 ;
wire un4_v_high_s_4_62 ;
wire un4_v_low_s_4_62 ;
wire un4_v_high_s_3_62 ;
wire un4_v_low_s_3_62 ;
wire un4_v_high_s_2_62 ;
wire un4_v_low_s_2_62 ;
wire un4_v_high_s_1_62 ;
wire un4_v_low_s_1_62 ;
wire v_diff_1_axb_0 ;
wire v_diff_1_axb_1 ;
wire v_diff_1_axb_2 ;
wire v_diff_1_axb_3 ;
wire v_diff_1_axb_4 ;
wire v_diff_1_axb_5 ;
wire v_diff_1_axb_6 ;
wire v_diff_1_axb_7 ;
wire un4_v_low_axb_1 ;
wire un4_v_low_axb_2 ;
wire un4_v_low_axb_3 ;
wire un4_v_low_axb_4 ;
wire un4_v_low_axb_5 ;
wire un4_v_low_axb_6 ;
wire un4_v_low_axb_7 ;
wire un4_v_high_axb_0 ;
wire un4_v_high_axb_1 ;
wire un4_v_high_axb_2 ;
wire un4_v_high_axb_3 ;
wire un4_v_high_axb_4 ;
wire un4_v_high_axb_5 ;
wire un4_v_high_axb_6 ;
wire un4_v_high_axb_7 ;
wire N_1108 ;
wire un4_v_high_axb_8 ;
wire un4_v_low_axb_8 ;
wire v_diff_1_axb_8 ;
wire un4_v_low_axb_0 ;
wire un4_v_high_cry_7 ;
wire un4_v_high_cry_6 ;
wire un4_v_high_cry_5 ;
wire un4_v_high_cry_4 ;
wire un4_v_high_cry_3 ;
wire un4_v_high_cry_2 ;
wire un4_v_high_cry_1 ;
wire un4_v_high_cry_0 ;
wire GND ;
wire un4_v_low_cry_7 ;
wire un4_v_low_cry_6 ;
wire un4_v_low_cry_5 ;
wire un4_v_low_cry_4 ;
wire un4_v_low_cry_3 ;
wire un4_v_low_cry_2 ;
wire un4_v_low_cry_1 ;
wire un4_v_low_cry_0 ;
wire v_diff_1_cry_7 ;
wire v_diff_1_cry_6 ;
wire v_diff_1_cry_5 ;
wire v_diff_1_cry_4 ;
wire v_diff_1_cry_3 ;
wire v_diff_1_cry_2 ;
wire v_diff_1_cry_1 ;
wire v_diff_1_cry_0 ;
wire N_1 ;
input p_desc2549_p_O_FD ;
input p_desc2550_p_O_FD ;
input p_m_axis_outdec_tdata_Z_p_O_FDRE ;
input p_desc2579_p_O_FDRE ;
// instances
  FDR desc2543(.Q(acs_prob_tdata_60[1:1]),.D(m_axis_outprob_tdata_8_0[1:1]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  FDR desc2544(.Q(acs_prob_tdata_60[2:2]),.D(m_axis_outprob_tdata_8_0[2:2]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  FDR desc2545(.Q(acs_prob_tdata_60[3:3]),.D(m_axis_outprob_tdata_8_0[3:3]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  FDR desc2546(.Q(acs_prob_tdata_60[4:4]),.D(m_axis_outprob_tdata_8_0[4:4]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  FDR desc2547(.Q(acs_prob_tdata_60[5:5]),.D(m_axis_outprob_tdata_8_0[5:5]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  FDR desc2548(.Q(acs_prob_tdata_60[6:6]),.D(m_axis_outprob_tdata_8_0[6:6]),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU));
  p_O_FD desc2549(.Q(acs_prob_tdata_60[7:7]),.D(m_axis_outprob_tdata_8_0_e[7:7]),.C(aclk),.E(p_desc2549_p_O_FD));
  p_O_FD desc2550(.Q(acs_prob_tdata_60[8:8]),.D(m_axis_outprob_tdata_8_0_e[8:8]),.C(aclk),.E(p_desc2550_p_O_FD));
  LUT6 desc2551(.I0(un4_v_high_s_7_62),.I1(un4_v_low_s_7_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[7:7]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG7GU),.O(m_axis_outprob_tdata_8_0_e[7:7]));
defparam desc2551.INIT=64'hFFFFFFFFACACFF00;
  LUT6 desc2552(.I0(un4_v_high_s_8_62),.I1(un4_v_low_s_8_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[8:8]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.I5(s_axis_inbranch_tlast_d_RNIG7GU),.O(m_axis_outprob_tdata_8_0_e[8:8]));
defparam desc2552.INIT=64'hFFFFFFFFACACFF00;
  LUT5 desc2553(.I0(un4_v_high_s_6_62),.I1(un4_v_low_s_6_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[6:6]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[6:6]));
defparam desc2553.INIT=32'hACACFF00;
  LUT5 desc2554(.I0(un4_v_high_s_5_62),.I1(un4_v_low_s_5_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[5:5]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[5:5]));
defparam desc2554.INIT=32'hACACFF00;
  LUT5 desc2555(.I0(un4_v_high_s_4_62),.I1(un4_v_low_s_4_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[4:4]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[4:4]));
defparam desc2555.INIT=32'hACACFF00;
  LUT5 desc2556(.I0(un4_v_high_s_3_62),.I1(un4_v_low_s_3_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[3:3]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[3:3]));
defparam desc2556.INIT=32'hACACFF00;
  LUT5 desc2557(.I0(un4_v_high_s_2_62),.I1(un4_v_low_s_2_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[2:2]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[2:2]));
defparam desc2557.INIT=32'hACACFF00;
  LUT5 desc2558(.I0(un4_v_high_s_1_62),.I1(un4_v_low_s_1_62),.I2(v_diff_1[8:8]),.I3(acs_prob_tdata_60[1:1]),.I4(s_axis_inbranch_tlast_d_1_sqmuxa_i),.O(m_axis_outprob_tdata_8_0[1:1]));
defparam desc2558.INIT=32'hACACFF00;
  p_O_FDRE m_axis_outdec_tdata_Z(.Q(acs_dec_tdata[60:60]),.D(v_diff_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un1_s_axis_inbranch_tvalid),.E(p_m_axis_outdec_tdata_Z_p_O_FDRE));
  LUT4 desc2559(.I0(acs_prob_tdata_56[0:0]),.I1(acs_prob_tdata_57[0:0]),.I2(branch_tdata_1_0_rep2),.I3(branch_tdata_2_0_rep2),.O(v_diff_1_axb_0));
defparam desc2559.INIT=16'h9669;
  LUT2 desc2560(.I0(un4_v_high_s_1_62),.I1(un4_v_low_s_1_62),.O(v_diff_1_axb_1));
defparam desc2560.INIT=4'h9;
  LUT2 desc2561(.I0(un4_v_high_s_2_62),.I1(un4_v_low_s_2_62),.O(v_diff_1_axb_2));
defparam desc2561.INIT=4'h9;
  LUT2 desc2562(.I0(un4_v_high_s_3_62),.I1(un4_v_low_s_3_62),.O(v_diff_1_axb_3));
defparam desc2562.INIT=4'h9;
  LUT2 desc2563(.I0(un4_v_high_s_4_62),.I1(un4_v_low_s_4_62),.O(v_diff_1_axb_4));
defparam desc2563.INIT=4'h9;
  LUT2 desc2564(.I0(un4_v_high_s_5_62),.I1(un4_v_low_s_5_62),.O(v_diff_1_axb_5));
defparam desc2564.INIT=4'h9;
  LUT2 desc2565(.I0(un4_v_high_s_6_62),.I1(un4_v_low_s_6_62),.O(v_diff_1_axb_6));
defparam desc2565.INIT=4'h9;
  LUT2 desc2566(.I0(un4_v_high_s_7_62),.I1(un4_v_low_s_7_62),.O(v_diff_1_axb_7));
defparam desc2566.INIT=4'h9;
  LUT2 un4_v_low_axb_1_cZ(.I0(acs_prob_tdata_56[1:1]),.I1(branch_tdata_1_1),.O(un4_v_low_axb_1));
defparam un4_v_low_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_2_cZ(.I0(acs_prob_tdata_56[2:2]),.I1(branch_tdata_1_2),.O(un4_v_low_axb_2));
defparam un4_v_low_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_3_cZ(.I0(acs_prob_tdata_56[3:3]),.I1(branch_tdata_1_3),.O(un4_v_low_axb_3));
defparam un4_v_low_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_4_cZ(.I0(acs_prob_tdata_56[4:4]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_4));
defparam un4_v_low_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_5_cZ(.I0(acs_prob_tdata_56[5:5]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_5));
defparam un4_v_low_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_6_cZ(.I0(acs_prob_tdata_56[6:6]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_6));
defparam un4_v_low_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_7_cZ(.I0(acs_prob_tdata_56[7:7]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_7));
defparam un4_v_low_axb_7_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_0_cZ(.I0(acs_prob_tdata_57[0:0]),.I1(branch_tdata_2_0_rep1),.O(un4_v_high_axb_0));
defparam un4_v_high_axb_0_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_1_cZ(.I0(acs_prob_tdata_57[1:1]),.I1(branch_tdata_2_1),.O(un4_v_high_axb_1));
defparam un4_v_high_axb_1_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_2_cZ(.I0(acs_prob_tdata_57[2:2]),.I1(branch_tdata_2_2),.O(un4_v_high_axb_2));
defparam un4_v_high_axb_2_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_3_cZ(.I0(acs_prob_tdata_57[3:3]),.I1(branch_tdata_2_3),.O(un4_v_high_axb_3));
defparam un4_v_high_axb_3_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_4_cZ(.I0(acs_prob_tdata_57[4:4]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_4));
defparam un4_v_high_axb_4_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_5_cZ(.I0(acs_prob_tdata_57[5:5]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_5));
defparam un4_v_high_axb_5_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_6_cZ(.I0(acs_prob_tdata_57[6:6]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_6));
defparam un4_v_high_axb_6_cZ.INIT=4'h6;
  LUT2 un4_v_high_axb_7_cZ(.I0(acs_prob_tdata_57[7:7]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_7));
defparam un4_v_high_axb_7_cZ.INIT=4'h6;
  FDR s_axis_inbranch_tlast_d_Z(.Q(s_axis_inbranch_tlast_d),.D(s_axis_inbranch_tlast_d_0),.C(aclk),.R(aresetn_i));
  LUT5_L desc2567(.I0(acs_prob_tdata_56[0:0]),.I1(acs_prob_tdata_57[0:0]),.I2(branch_tdata_1_0),.I3(branch_tdata_2_0),.I4(v_diff_1[8:8]),.LO(N_1108));
defparam desc2567.INIT=32'h33CC5A5A;
  LUT2 un4_v_high_axb_8_cZ(.I0(acs_prob_tdata_57[8:8]),.I1(branch_tdata_2_5),.O(un4_v_high_axb_8));
defparam un4_v_high_axb_8_cZ.INIT=4'h6;
  LUT2 un4_v_low_axb_8_cZ(.I0(acs_prob_tdata_56[8:8]),.I1(branch_tdata_1_5),.O(un4_v_low_axb_8));
defparam un4_v_low_axb_8_cZ.INIT=4'h6;
  LUT2 desc2568(.I0(un4_v_high_s_8_62),.I1(un4_v_low_s_8_62),.O(v_diff_1_axb_8));
defparam desc2568.INIT=4'h9;
  LUT6 desc2569(.I0(m_axis_outdec_tvalid_int),.I1(write_ram_fsm_4),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(branch_tvalid),.I5(N_1756_1),.O(un1_s_axis_inbranch_tvalid));
defparam desc2569.INIT=64'h5557000055550000;
  LUT4 s_axis_inbranch_tlast_d_RNIU4BR(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(branch_tvalid),.I3(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_1_sqmuxa_i));
defparam s_axis_inbranch_tlast_d_RNIU4BR.INIT=16'hBAFA;
  LUT5 s_axis_inbranch_tlast_d_RNIG7GU_cZ(.I0(aresetn),.I1(s_axis_inbranch_tlast_d),.I2(m_axis_outdec_tvalid_int),.I3(branch_tvalid),.I4(un27_s_axis_input_tready_int),.O(s_axis_inbranch_tlast_d_RNIG7GU));
defparam s_axis_inbranch_tlast_d_RNIG7GU_cZ.INIT=32'hD5DD55DD;
  LUT2 un4_v_low_axb_0_cZ(.I0(acs_prob_tdata_56[0:0]),.I1(branch_tdata_1_fast),.O(un4_v_low_axb_0));
defparam un4_v_low_axb_0_cZ.INIT=4'h6;
  FDR m_axis_outdec_tvalid_int_Z(.Q(m_axis_outdec_tvalid_int),.D(un1_s_axis_inbranch_tvalid_RNIB0PO_O6),.C(aclk),.R(aresetn_i));
  XORCY un4_v_high_s_8(.LI(un4_v_high_axb_8),.CI(un4_v_high_cry_7),.O(un4_v_high_s_8_62));
  XORCY un4_v_high_s_7(.LI(un4_v_high_axb_7),.CI(un4_v_high_cry_6),.O(un4_v_high_s_7_62));
  MUXCY_L un4_v_high_cry_7_cZ(.DI(acs_prob_tdata_57[7:7]),.CI(un4_v_high_cry_6),.S(un4_v_high_axb_7),.LO(un4_v_high_cry_7));
  XORCY un4_v_high_s_6(.LI(un4_v_high_axb_6),.CI(un4_v_high_cry_5),.O(un4_v_high_s_6_62));
  MUXCY_L un4_v_high_cry_6_cZ(.DI(acs_prob_tdata_57[6:6]),.CI(un4_v_high_cry_5),.S(un4_v_high_axb_6),.LO(un4_v_high_cry_6));
  XORCY un4_v_high_s_5(.LI(un4_v_high_axb_5),.CI(un4_v_high_cry_4),.O(un4_v_high_s_5_62));
  MUXCY_L un4_v_high_cry_5_cZ(.DI(acs_prob_tdata_57[5:5]),.CI(un4_v_high_cry_4),.S(un4_v_high_axb_5),.LO(un4_v_high_cry_5));
  XORCY un4_v_high_s_4(.LI(un4_v_high_axb_4),.CI(un4_v_high_cry_3),.O(un4_v_high_s_4_62));
  MUXCY_L un4_v_high_cry_4_cZ(.DI(acs_prob_tdata_57[4:4]),.CI(un4_v_high_cry_3),.S(un4_v_high_axb_4),.LO(un4_v_high_cry_4));
  XORCY un4_v_high_s_3(.LI(un4_v_high_axb_3),.CI(un4_v_high_cry_2),.O(un4_v_high_s_3_62));
  MUXCY_L un4_v_high_cry_3_cZ(.DI(acs_prob_tdata_57[3:3]),.CI(un4_v_high_cry_2),.S(un4_v_high_axb_3),.LO(un4_v_high_cry_3));
  XORCY un4_v_high_s_2(.LI(un4_v_high_axb_2),.CI(un4_v_high_cry_1),.O(un4_v_high_s_2_62));
  MUXCY_L un4_v_high_cry_2_cZ(.DI(acs_prob_tdata_57[2:2]),.CI(un4_v_high_cry_1),.S(un4_v_high_axb_2),.LO(un4_v_high_cry_2));
  XORCY un4_v_high_s_1(.LI(un4_v_high_axb_1),.CI(un4_v_high_cry_0),.O(un4_v_high_s_1_62));
  MUXCY_L un4_v_high_cry_1_cZ(.DI(acs_prob_tdata_57[1:1]),.CI(un4_v_high_cry_0),.S(un4_v_high_axb_1),.LO(un4_v_high_cry_1));
  MUXCY_L un4_v_high_cry_0_cZ(.DI(acs_prob_tdata_57[0:0]),.CI(GND),.S(un4_v_high_axb_0),.LO(un4_v_high_cry_0));
  XORCY un4_v_low_s_8(.LI(un4_v_low_axb_8),.CI(un4_v_low_cry_7),.O(un4_v_low_s_8_62));
  XORCY un4_v_low_s_7(.LI(un4_v_low_axb_7),.CI(un4_v_low_cry_6),.O(un4_v_low_s_7_62));
  MUXCY_L un4_v_low_cry_7_cZ(.DI(acs_prob_tdata_56[7:7]),.CI(un4_v_low_cry_6),.S(un4_v_low_axb_7),.LO(un4_v_low_cry_7));
  XORCY un4_v_low_s_6(.LI(un4_v_low_axb_6),.CI(un4_v_low_cry_5),.O(un4_v_low_s_6_62));
  MUXCY_L un4_v_low_cry_6_cZ(.DI(acs_prob_tdata_56[6:6]),.CI(un4_v_low_cry_5),.S(un4_v_low_axb_6),.LO(un4_v_low_cry_6));
  XORCY un4_v_low_s_5(.LI(un4_v_low_axb_5),.CI(un4_v_low_cry_4),.O(un4_v_low_s_5_62));
  MUXCY_L un4_v_low_cry_5_cZ(.DI(acs_prob_tdata_56[5:5]),.CI(un4_v_low_cry_4),.S(un4_v_low_axb_5),.LO(un4_v_low_cry_5));
  XORCY un4_v_low_s_4(.LI(un4_v_low_axb_4),.CI(un4_v_low_cry_3),.O(un4_v_low_s_4_62));
  MUXCY_L un4_v_low_cry_4_cZ(.DI(acs_prob_tdata_56[4:4]),.CI(un4_v_low_cry_3),.S(un4_v_low_axb_4),.LO(un4_v_low_cry_4));
  XORCY un4_v_low_s_3(.LI(un4_v_low_axb_3),.CI(un4_v_low_cry_2),.O(un4_v_low_s_3_62));
  MUXCY_L un4_v_low_cry_3_cZ(.DI(acs_prob_tdata_56[3:3]),.CI(un4_v_low_cry_2),.S(un4_v_low_axb_3),.LO(un4_v_low_cry_3));
  XORCY un4_v_low_s_2(.LI(un4_v_low_axb_2),.CI(un4_v_low_cry_1),.O(un4_v_low_s_2_62));
  MUXCY_L un4_v_low_cry_2_cZ(.DI(acs_prob_tdata_56[2:2]),.CI(un4_v_low_cry_1),.S(un4_v_low_axb_2),.LO(un4_v_low_cry_2));
  XORCY un4_v_low_s_1(.LI(un4_v_low_axb_1),.CI(un4_v_low_cry_0),.O(un4_v_low_s_1_62));
  MUXCY_L un4_v_low_cry_1_cZ(.DI(acs_prob_tdata_56[1:1]),.CI(un4_v_low_cry_0),.S(un4_v_low_axb_1),.LO(un4_v_low_cry_1));
  MUXCY_L un4_v_low_cry_0_cZ(.DI(acs_prob_tdata_56[0:0]),.CI(GND),.S(un4_v_low_axb_0),.LO(un4_v_low_cry_0));
  XORCY desc2570(.LI(v_diff_1_axb_8),.CI(v_diff_1_cry_7),.O(v_diff_1[8:8]));
  MUXCY_L desc2571(.DI(un4_v_low_s_7_62),.CI(v_diff_1_cry_6),.S(v_diff_1_axb_7),.LO(v_diff_1_cry_7));
  MUXCY_L desc2572(.DI(un4_v_low_s_6_62),.CI(v_diff_1_cry_5),.S(v_diff_1_axb_6),.LO(v_diff_1_cry_6));
  MUXCY_L desc2573(.DI(un4_v_low_s_5_62),.CI(v_diff_1_cry_4),.S(v_diff_1_axb_5),.LO(v_diff_1_cry_5));
  MUXCY_L desc2574(.DI(un4_v_low_s_4_62),.CI(v_diff_1_cry_3),.S(v_diff_1_axb_4),.LO(v_diff_1_cry_4));
  MUXCY_L desc2575(.DI(un4_v_low_s_3_62),.CI(v_diff_1_cry_2),.S(v_diff_1_axb_3),.LO(v_diff_1_cry_3));
  MUXCY_L desc2576(.DI(un4_v_low_s_2_62),.CI(v_diff_1_cry_1),.S(v_diff_1_axb_2),.LO(v_diff_1_cry_2));
  MUXCY_L desc2577(.DI(un4_v_low_s_1_62),.CI(v_diff_1_cry_0),.S(v_diff_1_axb_1),.LO(v_diff_1_cry_1));
  MUXCY_L desc2578(.DI(un4_v_low_axb_0),.CI(VCC),.S(v_diff_1_axb_0),.LO(v_diff_1_cry_0));
  p_O_FDRE desc2579(.Q(acs_prob_tdata_60[0:0]),.D(N_1108),.C(aclk),.R(s_axis_inbranch_tlast_d_RNIG7GU),.CE(s_axis_inbranch_tlast_d_1_sqmuxa_i),.E(p_desc2579_p_O_FDRE));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc2580(.I0(s_axis_inbranch_tlast_d),.I1(m_axis_outdec_tvalid_int),.I2(un1_s_axis_inbranch_tvalid),.I3(un27_s_axis_input_tready_int),.O(un1_s_axis_inbranch_tvalid_RNIB0PO_O6));
defparam desc2580.INIT=16'hF4F0;
  LUT2 desc2581(.I0(branch_tlast),.I1(un1_s_axis_inbranch_tvalid),.O(s_axis_inbranch_tlast_d_0));
defparam desc2581.INIT=4'h8;
endmodule
module generic_sp_ram_inj (q_reg_1,addr_1,acs_dec_tdata,wen_ram,aclk);
output [63:0] q_reg_1 ;
input [6:0] addr_1 ;
input [63:0] acs_dec_tdata ;
input [1:1] wen_ram ;
input aclk ;
wire aclk ;
wire [3:0] sp_ram_sp_ram_0_0_DOPADOP ;
wire [3:0] sp_ram_sp_ram_0_0_DOPBDOP ;
wire VCC ;
wire GND ;
wire NC0 ;
wire NC1 ;
wire NC2 ;
wire NC3 ;
wire NC4 ;
wire NC5 ;
wire NC6 ;
wire NC7 ;
wire NC8 ;
wire NC9 ;
wire NC10 ;
wire NC11 ;
wire NC12 ;
wire NC13 ;
wire NC14 ;
wire NC15 ;
wire NC16 ;
wire NC17 ;
wire NC18 ;
wire NC19 ;
wire NC20 ;
// instances
  RAMB36E1 sp_ram_sp_ram_0_0(.DOADO({q_reg_1[47:47],q_reg_1[15:15],q_reg_1[46:46],q_reg_1[14:14],q_reg_1[45:45],q_reg_1[13:13],q_reg_1[44:44],q_reg_1[12:12],q_reg_1[43:43],q_reg_1[11:11],q_reg_1[42:42],q_reg_1[10:10],q_reg_1[41:41],q_reg_1[9:9],q_reg_1[40:40],q_reg_1[8:8],q_reg_1[39:39],q_reg_1[7:7],q_reg_1[38:38],q_reg_1[6:6],q_reg_1[37:37],q_reg_1[5:5],q_reg_1[36:36],q_reg_1[4:4],q_reg_1[35:35],q_reg_1[3:3],q_reg_1[34:34],q_reg_1[2:2],q_reg_1[33:33],q_reg_1[1:1],q_reg_1[32:32],q_reg_1[0:0]}),.DOBDO({q_reg_1[63:63],q_reg_1[31:31],q_reg_1[62:62],q_reg_1[30:30],q_reg_1[61:61],q_reg_1[29:29],q_reg_1[60:60],q_reg_1[28:28],q_reg_1[59:59],q_reg_1[27:27],q_reg_1[58:58],q_reg_1[26:26],q_reg_1[57:57],q_reg_1[25:25],q_reg_1[56:56],q_reg_1[24:24],q_reg_1[55:55],q_reg_1[23:23],q_reg_1[54:54],q_reg_1[22:22],q_reg_1[53:53],q_reg_1[21:21],q_reg_1[52:52],q_reg_1[20:20],q_reg_1[51:51],q_reg_1[19:19],q_reg_1[50:50],q_reg_1[18:18],q_reg_1[49:49],q_reg_1[17:17],q_reg_1[48:48],q_reg_1[16:16]}),.DOPADOP(sp_ram_sp_ram_0_0_DOPADOP[3:0]),.DOPBDOP(sp_ram_sp_ram_0_0_DOPBDOP[3:0]),.ECCPARITY({NC10,NC9,NC8,NC7,NC6,NC5,NC4,NC3}),.RDADDRECC({NC19,NC18,NC17,NC16,NC15,NC14,NC13,NC12,NC11}),.ADDRARDADDR({VCC,GND,GND,addr_1[6:0],GND,VCC,VCC,VCC,VCC,VCC}),.ADDRBWRADDR({VCC,GND,GND,addr_1[6:0],VCC,VCC,VCC,VCC,VCC,VCC}),.CASCADEINA(GND),.CASCADEINB(GND),.CLKARDCLK(aclk),.CLKBWRCLK(aclk),.DIADI({acs_dec_tdata[47:47],acs_dec_tdata[15:15],acs_dec_tdata[46:46],acs_dec_tdata[14:14],acs_dec_tdata[45:45],acs_dec_tdata[13:13],acs_dec_tdata[44:44],acs_dec_tdata[12:12],acs_dec_tdata[43:43],acs_dec_tdata[11:11],acs_dec_tdata[42:42],acs_dec_tdata[10:10],acs_dec_tdata[41:41],acs_dec_tdata[9:9],acs_dec_tdata[40:40],acs_dec_tdata[8:8],acs_dec_tdata[39:39],acs_dec_tdata[7:7],acs_dec_tdata[38:38],acs_dec_tdata[6:6],acs_dec_tdata[37:37],acs_dec_tdata[5:5],acs_dec_tdata[36:36],acs_dec_tdata[4:4],acs_dec_tdata[35:35],acs_dec_tdata[3:3],acs_dec_tdata[34:34],acs_dec_tdata[2:2],acs_dec_tdata[33:33],acs_dec_tdata[1:1],acs_dec_tdata[32:32],acs_dec_tdata[0:0]}),.DIBDI({acs_dec_tdata[63:63],acs_dec_tdata[31:31],acs_dec_tdata[62:62],acs_dec_tdata[30:30],acs_dec_tdata[61:61],acs_dec_tdata[29:29],acs_dec_tdata[60:60],acs_dec_tdata[28:28],acs_dec_tdata[59:59],acs_dec_tdata[27:27],acs_dec_tdata[58:58],acs_dec_tdata[26:26],acs_dec_tdata[57:57],acs_dec_tdata[25:25],acs_dec_tdata[56:56],acs_dec_tdata[24:24],acs_dec_tdata[55:55],acs_dec_tdata[23:23],acs_dec_tdata[54:54],acs_dec_tdata[22:22],acs_dec_tdata[53:53],acs_dec_tdata[21:21],acs_dec_tdata[52:52],acs_dec_tdata[20:20],acs_dec_tdata[51:51],acs_dec_tdata[19:19],acs_dec_tdata[50:50],acs_dec_tdata[18:18],acs_dec_tdata[49:49],acs_dec_tdata[17:17],acs_dec_tdata[48:48],acs_dec_tdata[16:16]}),.DIPADIP({GND,GND,GND,GND}),.DIPBDIP({GND,GND,GND,GND}),.ENARDEN(VCC),.ENBWREN(VCC),.INJECTDBITERR(GND),.INJECTSBITERR(GND),.REGCEAREGCE(GND),.REGCEB(GND),.RSTRAMARSTRAM(GND),.RSTRAMB(GND),.RSTREGARSTREG(GND),.RSTREGB(GND),.WEA({wen_ram[1:1],wen_ram[1:1],wen_ram[1:1],wen_ram[1:1]}),.WEBWE({GND,GND,GND,GND,wen_ram[1:1],wen_ram[1:1],wen_ram[1:1],wen_ram[1:1]}));
defparam sp_ram_sp_ram_0_0.RAM_MODE="TDP";
defparam sp_ram_sp_ram_0_0.READ_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.READ_WIDTH_B=36;
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_A="REGCE";
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_B="REGCE";
defparam sp_ram_sp_ram_0_0.SRVAL_A=36'h000000000;
defparam sp_ram_sp_ram_0_0.SRVAL_B=36'h000000000;
defparam sp_ram_sp_ram_0_0.WRITE_MODE_A="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_MODE_B="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_B=36;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module generic_sp_ram_1_inj (q_reg_2,addr_2,acs_dec_tdata,wen_ram,aclk);
output [63:0] q_reg_2 ;
input [6:0] addr_2 ;
input [63:0] acs_dec_tdata ;
input [2:2] wen_ram ;
input aclk ;
wire aclk ;
wire [3:0] sp_ram_sp_ram_0_0_DOPADOP_0 ;
wire [3:0] sp_ram_sp_ram_0_0_DOPBDOP_0 ;
wire VCC ;
wire GND ;
wire NC0 ;
wire NC1 ;
wire NC2 ;
wire NC3 ;
wire NC4 ;
wire NC5 ;
wire NC6 ;
wire NC7 ;
wire NC8 ;
wire NC9 ;
wire NC10 ;
wire NC11 ;
wire NC12 ;
wire NC13 ;
wire NC14 ;
wire NC15 ;
wire NC16 ;
wire NC17 ;
wire NC18 ;
wire NC19 ;
wire NC20 ;
// instances
  RAMB36E1 sp_ram_sp_ram_0_0(.DOADO({q_reg_2[47:47],q_reg_2[15:15],q_reg_2[46:46],q_reg_2[14:14],q_reg_2[45:45],q_reg_2[13:13],q_reg_2[44:44],q_reg_2[12:12],q_reg_2[43:43],q_reg_2[11:11],q_reg_2[42:42],q_reg_2[10:10],q_reg_2[41:41],q_reg_2[9:9],q_reg_2[40:40],q_reg_2[8:8],q_reg_2[39:39],q_reg_2[7:7],q_reg_2[38:38],q_reg_2[6:6],q_reg_2[37:37],q_reg_2[5:5],q_reg_2[36:36],q_reg_2[4:4],q_reg_2[35:35],q_reg_2[3:3],q_reg_2[34:34],q_reg_2[2:2],q_reg_2[33:33],q_reg_2[1:1],q_reg_2[32:32],q_reg_2[0:0]}),.DOBDO({q_reg_2[63:63],q_reg_2[31:31],q_reg_2[62:62],q_reg_2[30:30],q_reg_2[61:61],q_reg_2[29:29],q_reg_2[60:60],q_reg_2[28:28],q_reg_2[59:59],q_reg_2[27:27],q_reg_2[58:58],q_reg_2[26:26],q_reg_2[57:57],q_reg_2[25:25],q_reg_2[56:56],q_reg_2[24:24],q_reg_2[55:55],q_reg_2[23:23],q_reg_2[54:54],q_reg_2[22:22],q_reg_2[53:53],q_reg_2[21:21],q_reg_2[52:52],q_reg_2[20:20],q_reg_2[51:51],q_reg_2[19:19],q_reg_2[50:50],q_reg_2[18:18],q_reg_2[49:49],q_reg_2[17:17],q_reg_2[48:48],q_reg_2[16:16]}),.DOPADOP(sp_ram_sp_ram_0_0_DOPADOP_0[3:0]),.DOPBDOP(sp_ram_sp_ram_0_0_DOPBDOP_0[3:0]),.ECCPARITY({NC10,NC9,NC8,NC7,NC6,NC5,NC4,NC3}),.RDADDRECC({NC19,NC18,NC17,NC16,NC15,NC14,NC13,NC12,NC11}),.ADDRARDADDR({VCC,GND,GND,addr_2[6:0],GND,VCC,VCC,VCC,VCC,VCC}),.ADDRBWRADDR({VCC,GND,GND,addr_2[6:0],VCC,VCC,VCC,VCC,VCC,VCC}),.CASCADEINA(GND),.CASCADEINB(GND),.CLKARDCLK(aclk),.CLKBWRCLK(aclk),.DIADI({acs_dec_tdata[47:47],acs_dec_tdata[15:15],acs_dec_tdata[46:46],acs_dec_tdata[14:14],acs_dec_tdata[45:45],acs_dec_tdata[13:13],acs_dec_tdata[44:44],acs_dec_tdata[12:12],acs_dec_tdata[43:43],acs_dec_tdata[11:11],acs_dec_tdata[42:42],acs_dec_tdata[10:10],acs_dec_tdata[41:41],acs_dec_tdata[9:9],acs_dec_tdata[40:40],acs_dec_tdata[8:8],acs_dec_tdata[39:39],acs_dec_tdata[7:7],acs_dec_tdata[38:38],acs_dec_tdata[6:6],acs_dec_tdata[37:37],acs_dec_tdata[5:5],acs_dec_tdata[36:36],acs_dec_tdata[4:4],acs_dec_tdata[35:35],acs_dec_tdata[3:3],acs_dec_tdata[34:34],acs_dec_tdata[2:2],acs_dec_tdata[33:33],acs_dec_tdata[1:1],acs_dec_tdata[32:32],acs_dec_tdata[0:0]}),.DIBDI({acs_dec_tdata[63:63],acs_dec_tdata[31:31],acs_dec_tdata[62:62],acs_dec_tdata[30:30],acs_dec_tdata[61:61],acs_dec_tdata[29:29],acs_dec_tdata[60:60],acs_dec_tdata[28:28],acs_dec_tdata[59:59],acs_dec_tdata[27:27],acs_dec_tdata[58:58],acs_dec_tdata[26:26],acs_dec_tdata[57:57],acs_dec_tdata[25:25],acs_dec_tdata[56:56],acs_dec_tdata[24:24],acs_dec_tdata[55:55],acs_dec_tdata[23:23],acs_dec_tdata[54:54],acs_dec_tdata[22:22],acs_dec_tdata[53:53],acs_dec_tdata[21:21],acs_dec_tdata[52:52],acs_dec_tdata[20:20],acs_dec_tdata[51:51],acs_dec_tdata[19:19],acs_dec_tdata[50:50],acs_dec_tdata[18:18],acs_dec_tdata[49:49],acs_dec_tdata[17:17],acs_dec_tdata[48:48],acs_dec_tdata[16:16]}),.DIPADIP({GND,GND,GND,GND}),.DIPBDIP({GND,GND,GND,GND}),.ENARDEN(VCC),.ENBWREN(VCC),.INJECTDBITERR(GND),.INJECTSBITERR(GND),.REGCEAREGCE(GND),.REGCEB(GND),.RSTRAMARSTRAM(GND),.RSTRAMB(GND),.RSTREGARSTREG(GND),.RSTREGB(GND),.WEA({wen_ram[2:2],wen_ram[2:2],wen_ram[2:2],wen_ram[2:2]}),.WEBWE({GND,GND,GND,GND,wen_ram[2:2],wen_ram[2:2],wen_ram[2:2],wen_ram[2:2]}));
defparam sp_ram_sp_ram_0_0.RAM_MODE="TDP";
defparam sp_ram_sp_ram_0_0.READ_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.READ_WIDTH_B=36;
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_A="REGCE";
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_B="REGCE";
defparam sp_ram_sp_ram_0_0.SRVAL_A=36'h000000000;
defparam sp_ram_sp_ram_0_0.SRVAL_B=36'h000000000;
defparam sp_ram_sp_ram_0_0.WRITE_MODE_A="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_MODE_B="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_B=36;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module generic_sp_ram_2_inj (q_reg_3,addr_3,acs_dec_tdata,wen_ram,aclk);
output [63:0] q_reg_3 ;
input [6:0] addr_3 ;
input [63:0] acs_dec_tdata ;
input [3:3] wen_ram ;
input aclk ;
wire aclk ;
wire [3:0] sp_ram_sp_ram_0_0_DOPADOP_1 ;
wire [3:0] sp_ram_sp_ram_0_0_DOPBDOP_1 ;
wire VCC ;
wire GND ;
wire NC0 ;
wire NC1 ;
wire NC2 ;
wire NC3 ;
wire NC4 ;
wire NC5 ;
wire NC6 ;
wire NC7 ;
wire NC8 ;
wire NC9 ;
wire NC10 ;
wire NC11 ;
wire NC12 ;
wire NC13 ;
wire NC14 ;
wire NC15 ;
wire NC16 ;
wire NC17 ;
wire NC18 ;
wire NC19 ;
wire NC20 ;
// instances
  RAMB36E1 sp_ram_sp_ram_0_0(.DOADO({q_reg_3[47:47],q_reg_3[15:15],q_reg_3[46:46],q_reg_3[14:14],q_reg_3[45:45],q_reg_3[13:13],q_reg_3[44:44],q_reg_3[12:12],q_reg_3[43:43],q_reg_3[11:11],q_reg_3[42:42],q_reg_3[10:10],q_reg_3[41:41],q_reg_3[9:9],q_reg_3[40:40],q_reg_3[8:8],q_reg_3[39:39],q_reg_3[7:7],q_reg_3[38:38],q_reg_3[6:6],q_reg_3[37:37],q_reg_3[5:5],q_reg_3[36:36],q_reg_3[4:4],q_reg_3[35:35],q_reg_3[3:3],q_reg_3[34:34],q_reg_3[2:2],q_reg_3[33:33],q_reg_3[1:1],q_reg_3[32:32],q_reg_3[0:0]}),.DOBDO({q_reg_3[63:63],q_reg_3[31:31],q_reg_3[62:62],q_reg_3[30:30],q_reg_3[61:61],q_reg_3[29:29],q_reg_3[60:60],q_reg_3[28:28],q_reg_3[59:59],q_reg_3[27:27],q_reg_3[58:58],q_reg_3[26:26],q_reg_3[57:57],q_reg_3[25:25],q_reg_3[56:56],q_reg_3[24:24],q_reg_3[55:55],q_reg_3[23:23],q_reg_3[54:54],q_reg_3[22:22],q_reg_3[53:53],q_reg_3[21:21],q_reg_3[52:52],q_reg_3[20:20],q_reg_3[51:51],q_reg_3[19:19],q_reg_3[50:50],q_reg_3[18:18],q_reg_3[49:49],q_reg_3[17:17],q_reg_3[48:48],q_reg_3[16:16]}),.DOPADOP(sp_ram_sp_ram_0_0_DOPADOP_1[3:0]),.DOPBDOP(sp_ram_sp_ram_0_0_DOPBDOP_1[3:0]),.ECCPARITY({NC10,NC9,NC8,NC7,NC6,NC5,NC4,NC3}),.RDADDRECC({NC19,NC18,NC17,NC16,NC15,NC14,NC13,NC12,NC11}),.ADDRARDADDR({VCC,GND,GND,addr_3[6:0],GND,VCC,VCC,VCC,VCC,VCC}),.ADDRBWRADDR({VCC,GND,GND,addr_3[6:0],VCC,VCC,VCC,VCC,VCC,VCC}),.CASCADEINA(GND),.CASCADEINB(GND),.CLKARDCLK(aclk),.CLKBWRCLK(aclk),.DIADI({acs_dec_tdata[47:47],acs_dec_tdata[15:15],acs_dec_tdata[46:46],acs_dec_tdata[14:14],acs_dec_tdata[45:45],acs_dec_tdata[13:13],acs_dec_tdata[44:44],acs_dec_tdata[12:12],acs_dec_tdata[43:43],acs_dec_tdata[11:11],acs_dec_tdata[42:42],acs_dec_tdata[10:10],acs_dec_tdata[41:41],acs_dec_tdata[9:9],acs_dec_tdata[40:40],acs_dec_tdata[8:8],acs_dec_tdata[39:39],acs_dec_tdata[7:7],acs_dec_tdata[38:38],acs_dec_tdata[6:6],acs_dec_tdata[37:37],acs_dec_tdata[5:5],acs_dec_tdata[36:36],acs_dec_tdata[4:4],acs_dec_tdata[35:35],acs_dec_tdata[3:3],acs_dec_tdata[34:34],acs_dec_tdata[2:2],acs_dec_tdata[33:33],acs_dec_tdata[1:1],acs_dec_tdata[32:32],acs_dec_tdata[0:0]}),.DIBDI({acs_dec_tdata[63:63],acs_dec_tdata[31:31],acs_dec_tdata[62:62],acs_dec_tdata[30:30],acs_dec_tdata[61:61],acs_dec_tdata[29:29],acs_dec_tdata[60:60],acs_dec_tdata[28:28],acs_dec_tdata[59:59],acs_dec_tdata[27:27],acs_dec_tdata[58:58],acs_dec_tdata[26:26],acs_dec_tdata[57:57],acs_dec_tdata[25:25],acs_dec_tdata[56:56],acs_dec_tdata[24:24],acs_dec_tdata[55:55],acs_dec_tdata[23:23],acs_dec_tdata[54:54],acs_dec_tdata[22:22],acs_dec_tdata[53:53],acs_dec_tdata[21:21],acs_dec_tdata[52:52],acs_dec_tdata[20:20],acs_dec_tdata[51:51],acs_dec_tdata[19:19],acs_dec_tdata[50:50],acs_dec_tdata[18:18],acs_dec_tdata[49:49],acs_dec_tdata[17:17],acs_dec_tdata[48:48],acs_dec_tdata[16:16]}),.DIPADIP({GND,GND,GND,GND}),.DIPBDIP({GND,GND,GND,GND}),.ENARDEN(VCC),.ENBWREN(VCC),.INJECTDBITERR(GND),.INJECTSBITERR(GND),.REGCEAREGCE(GND),.REGCEB(GND),.RSTRAMARSTRAM(GND),.RSTRAMB(GND),.RSTREGARSTREG(GND),.RSTREGB(GND),.WEA({wen_ram[3:3],wen_ram[3:3],wen_ram[3:3],wen_ram[3:3]}),.WEBWE({GND,GND,GND,GND,wen_ram[3:3],wen_ram[3:3],wen_ram[3:3],wen_ram[3:3]}));
defparam sp_ram_sp_ram_0_0.RAM_MODE="TDP";
defparam sp_ram_sp_ram_0_0.READ_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.READ_WIDTH_B=36;
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_A="REGCE";
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_B="REGCE";
defparam sp_ram_sp_ram_0_0.SRVAL_A=36'h000000000;
defparam sp_ram_sp_ram_0_0.SRVAL_B=36'h000000000;
defparam sp_ram_sp_ram_0_0.WRITE_MODE_A="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_MODE_B="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_B=36;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module generic_sp_ram_3_inj (q_reg_0,addr_0,acs_dec_tdata,wen_ram,aclk);
output [63:0] q_reg_0 ;
input [6:0] addr_0 ;
input [63:0] acs_dec_tdata ;
input wen_ram ;
input aclk ;
wire aclk ;
wire [3:0] sp_ram_sp_ram_0_0_DOPADOP_2 ;
wire [3:0] sp_ram_sp_ram_0_0_DOPBDOP_2 ;
wire VCC ;
wire GND ;
wire NC0 ;
wire NC1 ;
wire NC2 ;
wire NC3 ;
wire NC4 ;
wire NC5 ;
wire NC6 ;
wire NC7 ;
wire NC8 ;
wire NC9 ;
wire NC10 ;
wire NC11 ;
wire NC12 ;
wire NC13 ;
wire NC14 ;
wire NC15 ;
wire NC16 ;
wire NC17 ;
wire NC18 ;
wire NC19 ;
wire NC20 ;
// instances
  RAMB36E1 sp_ram_sp_ram_0_0(.DOADO({q_reg_0[47:47],q_reg_0[15:15],q_reg_0[46:46],q_reg_0[14:14],q_reg_0[45:45],q_reg_0[13:13],q_reg_0[44:44],q_reg_0[12:12],q_reg_0[43:43],q_reg_0[11:11],q_reg_0[42:42],q_reg_0[10:10],q_reg_0[41:41],q_reg_0[9:9],q_reg_0[40:40],q_reg_0[8:8],q_reg_0[39:39],q_reg_0[7:7],q_reg_0[38:38],q_reg_0[6:6],q_reg_0[37:37],q_reg_0[5:5],q_reg_0[36:36],q_reg_0[4:4],q_reg_0[35:35],q_reg_0[3:3],q_reg_0[34:34],q_reg_0[2:2],q_reg_0[33:33],q_reg_0[1:1],q_reg_0[32:32],q_reg_0[0:0]}),.DOBDO({q_reg_0[63:63],q_reg_0[31:31],q_reg_0[62:62],q_reg_0[30:30],q_reg_0[61:61],q_reg_0[29:29],q_reg_0[60:60],q_reg_0[28:28],q_reg_0[59:59],q_reg_0[27:27],q_reg_0[58:58],q_reg_0[26:26],q_reg_0[57:57],q_reg_0[25:25],q_reg_0[56:56],q_reg_0[24:24],q_reg_0[55:55],q_reg_0[23:23],q_reg_0[54:54],q_reg_0[22:22],q_reg_0[53:53],q_reg_0[21:21],q_reg_0[52:52],q_reg_0[20:20],q_reg_0[51:51],q_reg_0[19:19],q_reg_0[50:50],q_reg_0[18:18],q_reg_0[49:49],q_reg_0[17:17],q_reg_0[48:48],q_reg_0[16:16]}),.DOPADOP(sp_ram_sp_ram_0_0_DOPADOP_2[3:0]),.DOPBDOP(sp_ram_sp_ram_0_0_DOPBDOP_2[3:0]),.ECCPARITY({NC10,NC9,NC8,NC7,NC6,NC5,NC4,NC3}),.RDADDRECC({NC19,NC18,NC17,NC16,NC15,NC14,NC13,NC12,NC11}),.ADDRARDADDR({VCC,GND,GND,addr_0[6:0],GND,VCC,VCC,VCC,VCC,VCC}),.ADDRBWRADDR({VCC,GND,GND,addr_0[6:0],VCC,VCC,VCC,VCC,VCC,VCC}),.CASCADEINA(GND),.CASCADEINB(GND),.CLKARDCLK(aclk),.CLKBWRCLK(aclk),.DIADI({acs_dec_tdata[47:47],acs_dec_tdata[15:15],acs_dec_tdata[46:46],acs_dec_tdata[14:14],acs_dec_tdata[45:45],acs_dec_tdata[13:13],acs_dec_tdata[44:44],acs_dec_tdata[12:12],acs_dec_tdata[43:43],acs_dec_tdata[11:11],acs_dec_tdata[42:42],acs_dec_tdata[10:10],acs_dec_tdata[41:41],acs_dec_tdata[9:9],acs_dec_tdata[40:40],acs_dec_tdata[8:8],acs_dec_tdata[39:39],acs_dec_tdata[7:7],acs_dec_tdata[38:38],acs_dec_tdata[6:6],acs_dec_tdata[37:37],acs_dec_tdata[5:5],acs_dec_tdata[36:36],acs_dec_tdata[4:4],acs_dec_tdata[35:35],acs_dec_tdata[3:3],acs_dec_tdata[34:34],acs_dec_tdata[2:2],acs_dec_tdata[33:33],acs_dec_tdata[1:1],acs_dec_tdata[32:32],acs_dec_tdata[0:0]}),.DIBDI({acs_dec_tdata[63:63],acs_dec_tdata[31:31],acs_dec_tdata[62:62],acs_dec_tdata[30:30],acs_dec_tdata[61:61],acs_dec_tdata[29:29],acs_dec_tdata[60:60],acs_dec_tdata[28:28],acs_dec_tdata[59:59],acs_dec_tdata[27:27],acs_dec_tdata[58:58],acs_dec_tdata[26:26],acs_dec_tdata[57:57],acs_dec_tdata[25:25],acs_dec_tdata[56:56],acs_dec_tdata[24:24],acs_dec_tdata[55:55],acs_dec_tdata[23:23],acs_dec_tdata[54:54],acs_dec_tdata[22:22],acs_dec_tdata[53:53],acs_dec_tdata[21:21],acs_dec_tdata[52:52],acs_dec_tdata[20:20],acs_dec_tdata[51:51],acs_dec_tdata[19:19],acs_dec_tdata[50:50],acs_dec_tdata[18:18],acs_dec_tdata[49:49],acs_dec_tdata[17:17],acs_dec_tdata[48:48],acs_dec_tdata[16:16]}),.DIPADIP({GND,GND,GND,GND}),.DIPBDIP({GND,GND,GND,GND}),.ENARDEN(VCC),.ENBWREN(VCC),.INJECTDBITERR(GND),.INJECTSBITERR(GND),.REGCEAREGCE(GND),.REGCEB(GND),.RSTRAMARSTRAM(GND),.RSTRAMB(GND),.RSTREGARSTREG(GND),.RSTREGB(GND),.WEA({wen_ram,wen_ram,wen_ram,wen_ram}),.WEBWE({GND,GND,GND,GND,wen_ram,wen_ram,wen_ram,wen_ram}));
defparam sp_ram_sp_ram_0_0.RAM_MODE="TDP";
defparam sp_ram_sp_ram_0_0.READ_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.READ_WIDTH_B=36;
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_A="REGCE";
defparam sp_ram_sp_ram_0_0.RSTREG_PRIORITY_B="REGCE";
defparam sp_ram_sp_ram_0_0.SRVAL_A=36'h000000000;
defparam sp_ram_sp_ram_0_0.SRVAL_B=36'h000000000;
defparam sp_ram_sp_ram_0_0.WRITE_MODE_A="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_MODE_B="NO_CHANGE";
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_A=36;
defparam sp_ram_sp_ram_0_0.WRITE_WIDTH_B=36;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module ram_ctrl_inj (acs_tlast,acs_tvalid,write_ram_fsm_1,write_ram_fsm_0,write_ram_fsm_4,ram_tlast,ram_last_tuser,s_axis_ctrl_tdata_16,s_axis_ctrl_tdata_17,s_axis_ctrl_tdata_18,s_axis_ctrl_tdata_19,s_axis_ctrl_tdata_20,s_axis_ctrl_tdata_21,s_axis_ctrl_tdata_22,s_axis_ctrl_tdata_0,s_axis_ctrl_tdata_1,s_axis_ctrl_tdata_2,s_axis_ctrl_tdata_3,s_axis_ctrl_tdata_4,s_axis_ctrl_tdata_5,s_axis_ctrl_tdata_6,ram_buffer_full,traceback_tvalid,ram_tvalid,ram_buffer_1_1,ram_buffer_0_2,ram_window_tuser,reorder_tvalid_fast,ram_buffer_0,ram_buffer_1,acs_dec_tdata,aresetn,reorder_tvalid_1_rep1,un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5,un1_s_axis_input_tvalid,aclk,write_ram_fsm_0_rep1,write_ram_fsm_0_rep2,write_ram_fsm_4_rep1,write_ram_fsm_4_rep2,aresetn_i,N_1756_1,reorder_tvalid_0_rep1,reorder_tvalid_0_rep2,N_99,s_axis_ctrl_tvalid,s_axis_ctrl_tready,un27_s_axis_input_tready_int);
input acs_tlast ;
input acs_tvalid ;
output write_ram_fsm_1 ;
output write_ram_fsm_0 ;
output write_ram_fsm_4 ;
output [1:0] ram_tlast ;
output [1:0] ram_last_tuser ;
input s_axis_ctrl_tdata_16 ;
input s_axis_ctrl_tdata_17 ;
input s_axis_ctrl_tdata_18 ;
input s_axis_ctrl_tdata_19 ;
input s_axis_ctrl_tdata_20 ;
input s_axis_ctrl_tdata_21 ;
input s_axis_ctrl_tdata_22 ;
input s_axis_ctrl_tdata_0 ;
input s_axis_ctrl_tdata_1 ;
input s_axis_ctrl_tdata_2 ;
input s_axis_ctrl_tdata_3 ;
input s_axis_ctrl_tdata_4 ;
input s_axis_ctrl_tdata_5 ;
input s_axis_ctrl_tdata_6 ;
output [1:0] ram_buffer_full ;
input [1:0] traceback_tvalid ;
output [1:0] ram_tvalid ;
output [63:0] ram_buffer_1_1 ;
output [63:0] ram_buffer_0_2 ;
output [1:0] ram_window_tuser ;
input [1:0] reorder_tvalid_fast ;
output [63:0] ram_buffer_0 ;
output [63:0] ram_buffer_1 ;
input [63:0] acs_dec_tdata ;
input aresetn ;
input reorder_tvalid_1_rep1 ;
output un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ;
input un1_s_axis_input_tvalid ;
input aclk ;
output write_ram_fsm_0_rep1 ;
output write_ram_fsm_0_rep2 ;
output write_ram_fsm_4_rep1 ;
output write_ram_fsm_4_rep2 ;
output aresetn_i ;
output N_1756_1 ;
input reorder_tvalid_0_rep1 ;
input reorder_tvalid_0_rep2 ;
input N_99 ;
input s_axis_ctrl_tvalid ;
output s_axis_ctrl_tready ;
output un27_s_axis_input_tready_int ;
wire write_ram_fsm_1 ;
wire write_ram_fsm_0 ;
wire write_ram_fsm_4 ;
wire s_axis_ctrl_tdata_16 ;
wire s_axis_ctrl_tdata_17 ;
wire s_axis_ctrl_tdata_18 ;
wire s_axis_ctrl_tdata_19 ;
wire s_axis_ctrl_tdata_20 ;
wire s_axis_ctrl_tdata_21 ;
wire s_axis_ctrl_tdata_22 ;
wire s_axis_ctrl_tdata_0 ;
wire s_axis_ctrl_tdata_1 ;
wire s_axis_ctrl_tdata_2 ;
wire s_axis_ctrl_tdata_3 ;
wire s_axis_ctrl_tdata_4 ;
wire s_axis_ctrl_tdata_5 ;
wire s_axis_ctrl_tdata_6 ;
wire aresetn ;
wire reorder_tvalid_1_rep1 ;
wire un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ;
wire un1_s_axis_input_tvalid ;
wire aclk ;
wire write_ram_fsm_0_rep1 ;
wire write_ram_fsm_0_rep2 ;
wire write_ram_fsm_4_rep1 ;
wire write_ram_fsm_4_rep2 ;
wire aresetn_i ;
wire N_1756_1 ;
wire reorder_tvalid_0_rep1 ;
wire reorder_tvalid_0_rep2 ;
wire N_99 ;
wire s_axis_ctrl_tvalid ;
wire s_axis_ctrl_tready ;
wire un27_s_axis_input_tready_int ;
wire un2_write_ram_ptr_3_iv_1_RNI880U2_O6 ;
wire un2_write_ram_ptr_2_iv_1_RNIGNT55_O6 ;
wire [1:0] read_ram_fsm_1 ;
wire next_traceback ;
wire [1:0] write_ram_ptr ;
wire [3:2] write_ram_fsm ;
wire [1:0] write_ram_ptr_fast ;
wire [3:3] read_ram_fsm_0_d_i_0 ;
wire [4:0] write_ram_fsm_fast ;
wire [1:0] read_ram_fsm_0 ;
wire [4:0] write_ram_fsm_srsts_0_e ;
wire [4:0] write_ram_fsm_srsts_fast_0_e ;
wire [4:0] write_ram_fsm_srsts_rep1_0_e ;
wire [4:0] write_ram_fsm_srsts_rep2_0_e ;
wire [4:4] write_ram_fsm_ns_i_0 ;
wire [2:0] write_ram_fsm_ns_0_0 ;
wire [3:3] write_ram_fsm_ns_i_o4_0_0 ;
wire [3:3] write_ram_fsm_nss_0 ;
wire [2:1] write_ram_fsm_nss ;
wire acquisition_length_fast ;
wire [4:0] window_length_fast ;
wire [6:0] acquisition_length ;
wire [6:0] window_length ;
wire [6:0] read_addr_ptr_1 ;
wire [6:0] read_addr_ptr_0 ;
wire [6:1] un64_m_axis_output_tready_a_5 ;
wire [6:1] un18_m_axis_output_tready ;
wire [1:0] m_axis_output_tlast_int ;
wire [1:0] m_axis_output_last_tuser_int ;
wire [1:0] read_ram_ptr_0 ;
wire read_ram_ptr_0_RNO ;
wire [1:0] read_ram_ptr_1 ;
wire read_ram_ptr_1_RNO ;
wire [1:0] ram_buffer_full_nss ;
wire [1:0] read_ram_fsm_0_nss ;
wire [1:0] read_ram_fsm_1_nss ;
wire [6:0] write_addr_ptr ;
wire [3:0] wen_ram ;
wire [3:0] wen_ramd_0 ;
wire [1:0] read_ram_ptr_0_fast ;
wire [1:0] read_ram_ptr_1_fast ;
wire [1:0] read_ram_fsm_1_fast ;
wire [1:0] read_ram_fsm_1_nss_fast ;
wire [1:0] read_ram_fsm_1_nss_rep1 ;
wire [1:0] read_ram_fsm_0_fast ;
wire [1:0] read_ram_fsm_0_nss_fast ;
wire [1:0] read_ram_fsm_0_nss_rep1 ;
wire [1:0] un9_s_axis_input_tvalid_0_data_tmp ;
wire [1:0] un30_m_axis_output_tready_0_data_tmp ;
wire [1:0] un64_m_axis_output_tready_0_data_tmp ;
wire [1:0] un23_m_axis_output_tready_0_data_tmp ;
wire [1:0] un57_m_axis_output_tready_0_data_tmp ;
wire [1:1] un2_write_ram_ptr_2_1 ;
wire [1:1] un2_write_ram_ptr_3_1 ;
wire [2:2] write_ram_fsm_ns_0_a4_0_0 ;
wire write_ram_fsm_ns_0_a4_2_1 ;
wire [6:6] un1_read_addr_ptr_0_1_sqmuxa_2_f1 ;
wire [6:0] read_last_addr_ptr ;
wire [6:0] read_last_addr_ptr_m ;
wire [6:0] read_last_addr_ptr_m_0 ;
wire [6:6] un1_read_addr_ptr_1_1_sqmuxa_2_f0_0 ;
wire [5:5] read_addr_ptr_0_m ;
wire [6:6] un1_read_addr_ptr_0_1_sqmuxa_2_f0_0 ;
wire [6:6] un1_read_addr_ptr_1_1_sqmuxa_2_f1 ;
wire [1:0] read_ram_ptr_d_1 ;
wire [63:0] q_reg_0 ;
wire [63:0] q_reg_1 ;
wire [63:0] q_reg_2 ;
wire [63:0] q_reg_3 ;
wire [1:0] read_ram_ptr_d_0 ;
wire [1:0] m_axis_output_window_tuser_int_RNO ;
wire m_axis_output_tvalid_int_RNO ;
wire [6:0] addr_1 ;
wire [6:0] addr_0 ;
wire [6:0] addr_3 ;
wire [6:0] addr_2 ;
wire [5:5] window_length_m_0 ;
wire [5:5] read_addr_ptr_1_m ;
wire [6:0] un1_write_addr_ptr_11 ;
wire [6:0] un1_write_addr_ptr_10 ;
wire [6:6] un1_write_addr_ptr_2 ;
wire [1:1] write_ram_fsm_ns_0_a4_0_RNI314E ;
wire [1:1] write_ram_fsm_ns_0_a4_0_RNI424E ;
wire [1:1] write_ram_fsm_ns_0_a4_0_RNI534E ;
wire [1:1] write_ram_fsm_ns_0_a4_0_RNITR4E ;
wire [1:1] write_ram_fsm_ns_0_a4_0_RNIUS4E ;
wire CO0_3 ;
wire SUM1_3_0 ;
wire GND ;
wire VCC ;
wire N_426_fast ;
wire CO0_4 ;
wire SUM1_4_0 ;
wire N_430_fast ;
wire write_window_complete ;
wire write_window_complete_RNIV26T_O6 ;
wire N_941s ;
wire un21_m_axis_output_tvalid_int ;
wire read_ram_fsm_1_1_rep1 ;
wire read_ram_fsm_1_0_rep1 ;
wire N_720 ;
wire N_1733 ;
wire write_last_window_complete ;
wire un44_m_axis_output_tready ;
wire N_745 ;
wire N_13 ;
wire N_709 ;
wire un106_addr ;
wire un42_addr ;
wire un3_addr ;
wire un74_addr ;
wire last_of_block ;
wire m_axis_output_tlast_int_0_sqmuxa_0 ;
wire last_of_block_0 ;
wire un1_write_ram_ptr_0_sqmuxa ;
wire un9_s_axis_input_tvalid ;
wire N_1740 ;
wire N_2332_i_fast_0 ;
wire read_ram_fsm_0_0_rep1 ;
wire read_ram_fsm_0_1_rep1 ;
wire read_addr_ptr_0_1_sqmuxa_1 ;
wire un13_write_last_window_complete ;
wire un1_m_axis_output_window_tuser_int_0_sqmuxa_set_0 ;
wire un1_write_ram_ptr_0_sqmuxa_sx ;
wire N_1739 ;
wire N_1731 ;
wire write_ram_fsm_1_sqmuxa ;
wire SUM1_5 ;
wire N_2332_i_0 ;
wire SUM1_5_fast ;
wire N_1743 ;
wire un3_s_axis_input_tready_int_li ;
wire un64_m_axis_output_tready_a_5_cry_0_RNO ;
wire un64_m_axis_output_tready_a_5_axb_1 ;
wire un64_m_axis_output_tready_a_5_axb_2 ;
wire un64_m_axis_output_tready_a_5_axb_3 ;
wire un64_m_axis_output_tready_a_5_axb_4 ;
wire un64_m_axis_output_tready_a_5_axb_5 ;
wire un18_m_axis_output_tready_cry_0_RNO ;
wire un18_m_axis_output_tready_axb_1 ;
wire un18_m_axis_output_tready_axb_2 ;
wire un18_m_axis_output_tready_axb_3 ;
wire un18_m_axis_output_tready_axb_4 ;
wire un18_m_axis_output_tready_axb_5 ;
wire un21_m_axis_output_tready_axb_1 ;
wire un21_m_axis_output_tready_axb_2 ;
wire un21_m_axis_output_tready_axb_3 ;
wire un21_m_axis_output_tready_axb_4 ;
wire un21_m_axis_output_tready_axb_5 ;
wire read_ram_fsm_1_0_sqmuxa_1_scy ;
wire un21_m_axis_output_tready_s_6 ;
wire un57_m_axis_output_tready_0_N_3_i ;
wire un23_m_axis_output_tready_0_N_3_i ;
wire un64_m_axis_output_tready_0_N_3_i ;
wire un30_m_axis_output_tready_0_N_3_i ;
wire write_window_complete_0 ;
wire write_last_window_complete_0 ;
wire wen_ram_0_sqmuxa_3 ;
wire un1_read_addr_ptr_0_2_axb_0 ;
wire un1_read_addr_ptr_0_2_s_1 ;
wire un1_read_addr_ptr_0_2_s_2 ;
wire un1_read_addr_ptr_0_2_s_3 ;
wire un1_read_addr_ptr_0_2_s_4 ;
wire un1_read_addr_ptr_0_2_s_5 ;
wire un1_read_addr_ptr_0_2_s_6 ;
wire un1_read_addr_ptr_1_2_axb_0 ;
wire un1_read_addr_ptr_1_2_s_1 ;
wire un1_read_addr_ptr_1_2_s_2 ;
wire un1_read_addr_ptr_1_2_s_3 ;
wire un1_read_addr_ptr_1_2_s_4 ;
wire un1_read_addr_ptr_1_2_s_5 ;
wire un1_read_addr_ptr_1_2_s_6 ;
wire N_1785 ;
wire un9_s_axis_input_tvalid_0_I_19_RNIUQCT ;
wire N_1786 ;
wire N_1787 ;
wire N_1788 ;
wire N_1789 ;
wire N_1790 ;
wire N_1791 ;
wire N_425_fast ;
wire N_429_fast ;
wire un9_s_axis_input_tvalid_0_I_19_RNO ;
wire un30_m_axis_output_tready ;
wire un64_m_axis_output_tready ;
wire un23_m_axis_output_tready ;
wire un57_m_axis_output_tready ;
wire read_ram_fsm_1_0_sqmuxa_1 ;
wire read_ram_fsm_0_0_sqmuxa ;
wire N_54_mux ;
wire un10_m_axis_output_tready ;
wire N_13_0 ;
wire N_54_mux_0 ;
wire N_41_mux ;
wire g5_0_0_0 ;
wire g5_0_0 ;
wire un15_s_axis_input_tready_int_li ;
wire N_1872 ;
wire un9_s_axis_input_tvalid_0_I_19_RNIN8NO ;
wire un1_wen_ram_1_sqmuxa_1_i ;
wire N_1875 ;
wire N_1874 ;
wire N_1873 ;
wire N_1747 ;
wire m33_0_0 ;
wire m33_0 ;
wire un1_read_ram_ptr_1_1_sqmuxa_0 ;
wire read_ram_fsm_0_2_sqmuxa_0 ;
wire read_addr_ptr_0_1_sqmuxa_3 ;
wire read_addr_ptr_0_2_sqmuxa_1 ;
wire un1_read_addr_ptr_0_1_sqmuxa_1_1 ;
wire un16_addr ;
wire un87_addr ;
wire un55_addr ;
wire un119_addr ;
wire m_axis_output_tlast_int_0_sqmuxa_1_1 ;
wire un5_m_axis_output_tvalid_int ;
wire read_addr_ptr_0_1_sqmuxa_3_RNIVHT32 ;
wire un1_read_addr_ptr_1_1_sqmuxa_0 ;
wire read_addr_ptr_1_2_sqmuxa_1 ;
wire read_addr_ptr_1_1_sqmuxa_3 ;
wire read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ ;
wire un1_read_addr_ptr_0_2_axb_5 ;
wire un1_ram_buffer_05_4 ;
wire un1_read_addr_ptr_1_2_axb_1 ;
wire un1_read_addr_ptr_1_2_cry_0_RNO ;
wire un1_read_addr_ptr_1_2_axb_3 ;
wire un1_read_addr_ptr_1_2_axb_4 ;
wire un1_read_addr_ptr_1_2_axb_6 ;
wire un1_read_addr_ptr_1_2_axb_2 ;
wire un1_ram_buffer_05_5 ;
wire un1_read_addr_ptr_0_2_axb_4 ;
wire un1_read_addr_ptr_0_2_axb_6 ;
wire un1_read_addr_ptr_0_2_cry_0_RNO ;
wire un1_read_addr_ptr_0_2_axb_1 ;
wire un1_read_addr_ptr_0_2_axb_2 ;
wire un1_read_addr_ptr_0_2_axb_3 ;
wire un1_write_addr_ptr_cry_0_cy ;
wire wen_ram_0_sqmuxa_3_ci ;
wire un1_write_addr_ptr_0_cry_0_cy ;
wire read_ram_fsm_1_2_sqmuxa_i_a2_0 ;
wire un21_m_axis_output_tready_axb_6 ;
wire un21_m_axis_output_tready_axb_0 ;
wire un18_m_axis_output_tready_axb_6 ;
wire un64_m_axis_output_tready_a_5_axb_6 ;
wire m33_1 ;
wire m33_0_2 ;
wire un6_m_axis_output_tready_3 ;
wire un30_m_axis_output_tready_0_N_14 ;
wire un64_m_axis_output_tready_a_5_axb_0 ;
wire un64_m_axis_output_tready_0_N_11 ;
wire N_743 ;
wire un21_m_axis_output_tready_s_3 ;
wire un21_m_axis_output_tready_s_4 ;
wire un21_m_axis_output_tready_s_5 ;
wire un57_m_axis_output_tready_0_N_4 ;
wire un23_m_axis_output_tready_0_N_4 ;
wire un64_m_axis_output_tready_0_N_4 ;
wire un30_m_axis_output_tready_0_N_4 ;
wire un21_m_axis_output_tready_s_1 ;
wire un21_m_axis_output_tready_s_2 ;
wire un57_m_axis_output_tready_0_N_11 ;
wire un23_m_axis_output_tready_0_N_11 ;
wire un30_m_axis_output_tready_0_N_11 ;
wire un9_s_axis_input_tvalid_0_N_11 ;
wire N_1754 ;
wire m33_2 ;
wire N_2339 ;
wire un9_s_axis_input_tvalid_a_4_c4 ;
wire un1_read_ram_ptr_0_1_sqmuxa_1 ;
wire un1_read_addr_ptr_1_1_sqmuxa_1_1 ;
wire write_ram_ptr_0_sqmuxa_1 ;
wire un1_write_addr_ptr_0_axb_6 ;
wire un1_write_addr_ptr_axb_6 ;
wire un1_write_addr_ptr_axb_5 ;
wire un1_write_addr_ptr_axb_4 ;
wire un1_write_addr_ptr_axb_3 ;
wire un1_write_addr_ptr_axb_2 ;
wire un1_write_addr_ptr_axb_1 ;
wire un9_s_axis_input_tvalid_0_N_4 ;
wire un1_write_addr_ptr_axb_0 ;
wire un1_write_addr_ptr_0_axb_0 ;
wire un1_write_addr_ptr_0_cry_0_RNO ;
wire un1_write_addr_ptr_0_axb_1 ;
wire un1_write_addr_ptr_0_axb_2 ;
wire un1_write_addr_ptr_0_axb_3 ;
wire un1_write_addr_ptr_0_axb_4 ;
wire un1_write_addr_ptr_0_axb_5 ;
wire un1_read_addr_ptr_1_2_axb_5 ;
wire un21_m_axis_output_tready_cry_5 ;
wire un21_m_axis_output_tready_cry_4 ;
wire un21_m_axis_output_tready_cry_3 ;
wire un21_m_axis_output_tready_cry_2 ;
wire un21_m_axis_output_tready_cry_1 ;
wire un21_m_axis_output_tready_cry_0 ;
wire un1_read_addr_ptr_0_2_cry_5 ;
wire un1_read_addr_ptr_0_2_cry_4 ;
wire un1_read_addr_ptr_0_2_cry_3 ;
wire un1_read_addr_ptr_0_2_cry_2 ;
wire un1_read_addr_ptr_0_2_cry_1 ;
wire un1_read_addr_ptr_0_2_cry_0 ;
wire un1_read_addr_ptr_1_2_cry_5 ;
wire un1_read_addr_ptr_1_2_cry_4 ;
wire un1_read_addr_ptr_1_2_cry_3 ;
wire un1_read_addr_ptr_1_2_cry_2 ;
wire un1_read_addr_ptr_1_2_cry_1 ;
wire un1_read_addr_ptr_1_2_cry_0 ;
wire un18_m_axis_output_tready_cry_5 ;
wire un18_m_axis_output_tready_cry_4 ;
wire un18_m_axis_output_tready_cry_3 ;
wire un18_m_axis_output_tready_cry_2 ;
wire un18_m_axis_output_tready_cry_1 ;
wire un18_m_axis_output_tready_cry_0 ;
wire un1_write_addr_ptr_0_cry_5 ;
wire un1_write_addr_ptr_0_cry_4 ;
wire un1_write_addr_ptr_0_cry_3 ;
wire un1_write_addr_ptr_0_cry_2 ;
wire un1_write_addr_ptr_0_cry_1 ;
wire un1_write_addr_ptr_0_cry_0 ;
wire un1_write_addr_ptr_cry_5 ;
wire un1_write_addr_ptr_cry_4 ;
wire un1_write_addr_ptr_cry_3 ;
wire un1_write_addr_ptr_cry_2 ;
wire un1_write_addr_ptr_cry_1 ;
wire un1_write_addr_ptr_cry_0 ;
wire un64_m_axis_output_tready_a_5_cry_5 ;
wire un64_m_axis_output_tready_a_5_cry_4 ;
wire un64_m_axis_output_tready_a_5_cry_3 ;
wire un64_m_axis_output_tready_a_5_cry_2 ;
wire un64_m_axis_output_tready_a_5_cry_1 ;
wire un64_m_axis_output_tready_a_5_cry_0 ;
wire N_1105 ;
wire N_1104 ;
wire N_1103 ;
wire N_1102 ;
wire N_968 ;
wire N_967 ;
wire N_966 ;
wire N_965 ;
wire N_964 ;
wire N_936 ;
wire N_935 ;
wire N_751 ;
wire N_750 ;
wire N_749 ;
wire N_748 ;
wire N_464 ;
wire N_463 ;
wire N_462 ;
wire N_461 ;
// instances
  LUT6_2 desc2582(.I0(write_window_complete),.I1(write_last_window_complete),.I2(next_traceback),.I3(un44_m_axis_output_tready),.I4(N_745),.I5(read_ram_fsm_1[0:0]),.O6(N_13),.O5(N_709));
defparam desc2582.INIT=64'hFF0000001F1F1F1F;
  FD desc2583(.Q(write_ram_fsm_0),.D(write_ram_fsm_srsts_0_e[0:0]),.C(aclk));
defparam desc2583.INIT=1'b0;
  FD desc2584(.Q(write_ram_fsm_fast[0:0]),.D(write_ram_fsm_srsts_fast_0_e[0:0]),.C(aclk));
defparam desc2584.INIT=1'b0;
  FD write_ram_fsm_0_rep1_Z(.Q(write_ram_fsm_0_rep1),.D(write_ram_fsm_srsts_rep1_0_e[0:0]),.C(aclk));
defparam write_ram_fsm_0_rep1_Z.INIT=1'b0;
  FD write_ram_fsm_0_rep2_Z(.Q(write_ram_fsm_0_rep2),.D(write_ram_fsm_srsts_rep2_0_e[0:0]),.C(aclk));
defparam write_ram_fsm_0_rep2_Z.INIT=1'b0;
  FD desc2585(.Q(write_ram_fsm_4),.D(write_ram_fsm_srsts_0_e[4:4]),.C(aclk));
defparam desc2585.INIT=1'b1;
  FD desc2586(.Q(write_ram_fsm_fast[4:4]),.D(write_ram_fsm_srsts_fast_0_e[4:4]),.C(aclk));
defparam desc2586.INIT=1'b1;
  FD write_ram_fsm_4_rep1_Z(.Q(write_ram_fsm_4_rep1),.D(write_ram_fsm_srsts_rep1_0_e[4:4]),.C(aclk));
defparam write_ram_fsm_4_rep1_Z.INIT=1'b1;
  FD write_ram_fsm_4_rep2_Z(.Q(write_ram_fsm_4_rep2),.D(write_ram_fsm_srsts_rep2_0_e[4:4]),.C(aclk));
defparam write_ram_fsm_4_rep2_Z.INIT=1'b1;
  FDR desc2587(.Q(write_ram_ptr[0:0]),.D(N_2332_i_0),.C(aclk),.R(aresetn_i));
  FDR desc2588(.Q(write_ram_ptr[1:1]),.D(SUM1_5),.C(aclk),.R(aresetn_i));
  FDR desc2589(.Q(write_ram_ptr_fast[0:0]),.D(N_2332_i_fast_0),.C(aclk),.R(aresetn_i));
  FDR desc2590(.Q(write_ram_ptr_fast[1:1]),.D(SUM1_5_fast),.C(aclk),.R(aresetn_i));
  LUT6 write_ram_fsm_0_rep2_RNO(.I0(acs_tlast),.I1(aresetn),.I2(N_1731),.I3(write_ram_fsm[2:2]),.I4(write_ram_fsm_0_rep2),.I5(write_ram_fsm_ns_i_0[4:4]),.O(write_ram_fsm_srsts_rep2_0_e[0:0]));
defparam write_ram_fsm_0_rep2_RNO.INIT=64'h000000000C0C8800;
  LUT6 write_ram_fsm_0_rep1_RNO(.I0(acs_tlast),.I1(aresetn),.I2(N_1731),.I3(write_ram_fsm[2:2]),.I4(write_ram_fsm_0_rep1),.I5(write_ram_fsm_ns_i_0[4:4]),.O(write_ram_fsm_srsts_rep1_0_e[0:0]));
defparam write_ram_fsm_0_rep1_RNO.INIT=64'h000000000C0C8800;
  LUT6 desc2591(.I0(acs_tlast),.I1(aresetn),.I2(N_1731),.I3(write_ram_fsm[2:2]),.I4(write_ram_fsm_fast[0:0]),.I5(write_ram_fsm_ns_i_0[4:4]),.O(write_ram_fsm_srsts_fast_0_e[0:0]));
defparam desc2591.INIT=64'h000000000C0C8800;
  LUT6 desc2592(.I0(acs_tlast),.I1(aresetn),.I2(N_1731),.I3(write_ram_fsm_0),.I4(write_ram_fsm[2:2]),.I5(write_ram_fsm_ns_i_0[4:4]),.O(write_ram_fsm_srsts_0_e[0:0]));
defparam desc2592.INIT=64'h000000000C880C00;
  LUT6 write_ram_fsm_4_rep2_RNO(.I0(aresetn),.I1(N_1731),.I2(N_1743),.I3(write_ram_fsm_0),.I4(write_ram_fsm_4_rep2),.I5(write_ram_fsm_ns_0_0[0:0]),.O(write_ram_fsm_srsts_rep2_0_e[4:4]));
defparam write_ram_fsm_4_rep2_RNO.INIT=64'hFFFFFFFFFDF5DD55;
  LUT6 write_ram_fsm_4_rep1_RNO(.I0(aresetn),.I1(N_1731),.I2(N_1743),.I3(write_ram_fsm_0),.I4(write_ram_fsm_4_rep1),.I5(write_ram_fsm_ns_0_0[0:0]),.O(write_ram_fsm_srsts_rep1_0_e[4:4]));
defparam write_ram_fsm_4_rep1_RNO.INIT=64'hFFFFFFFFFDF5DD55;
  LUT6 desc2593(.I0(aresetn),.I1(N_1731),.I2(N_1743),.I3(write_ram_fsm_0),.I4(write_ram_fsm_fast[4:4]),.I5(write_ram_fsm_ns_0_0[0:0]),.O(write_ram_fsm_srsts_fast_0_e[4:4]));
defparam desc2593.INIT=64'hFFFFFFFFFDF5DD55;
  LUT6 desc2594(.I0(aresetn),.I1(N_1731),.I2(N_1743),.I3(write_ram_fsm_0),.I4(write_ram_fsm_4),.I5(write_ram_fsm_ns_0_0[0:0]),.O(write_ram_fsm_srsts_0_e[4:4]));
defparam desc2594.INIT=64'hFFFFFFFFFDF5DD55;
  LUT5 desc2595(.I0(un1_s_axis_input_tvalid),.I1(un9_s_axis_input_tvalid),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(write_ram_ptr_fast[1:1]),.I4(write_ram_ptr[0:0]),.O(SUM1_5_fast));
defparam desc2595.INIT=32'h758AFF00;
  LUT6 desc2596(.I0(aresetn),.I1(N_1731),.I2(N_1740),.I3(un3_s_axis_input_tready_int_li),.I4(write_ram_fsm_1),.I5(write_ram_fsm_ns_i_o4_0_0[3:3]),.O(write_ram_fsm_nss_0[3:3]));
defparam desc2596.INIT=64'h2222000022220200;
  FD desc2597(.Q(write_ram_fsm[2:2]),.D(write_ram_fsm_nss[2:2]),.C(aclk));
defparam desc2597.INIT=1'b0;
  FD desc2598(.Q(write_ram_fsm_1),.D(write_ram_fsm_nss_0[3:3]),.C(aclk));
defparam desc2598.INIT=1'b0;
  FD desc2599(.Q(write_ram_fsm[3:3]),.D(write_ram_fsm_nss[1:1]),.C(aclk));
defparam desc2599.INIT=1'b0;
  LUT2 desc2600(.I0(acquisition_length_fast),.I1(window_length_fast[0:0]),.O(un64_m_axis_output_tready_a_5_cry_0_RNO));
defparam desc2600.INIT=4'h9;
  LUT2 desc2601(.I0(acquisition_length[1:1]),.I1(window_length_fast[1:1]),.O(un64_m_axis_output_tready_a_5_axb_1));
defparam desc2601.INIT=4'h9;
  LUT2 desc2602(.I0(acquisition_length[2:2]),.I1(window_length_fast[2:2]),.O(un64_m_axis_output_tready_a_5_axb_2));
defparam desc2602.INIT=4'h9;
  LUT2 desc2603(.I0(acquisition_length[3:3]),.I1(window_length_fast[3:3]),.O(un64_m_axis_output_tready_a_5_axb_3));
defparam desc2603.INIT=4'h9;
  LUT2 desc2604(.I0(acquisition_length[4:4]),.I1(window_length_fast[4:4]),.O(un64_m_axis_output_tready_a_5_axb_4));
defparam desc2604.INIT=4'h9;
  LUT2 desc2605(.I0(acquisition_length[5:5]),.I1(window_length[5:5]),.O(un64_m_axis_output_tready_a_5_axb_5));
defparam desc2605.INIT=4'h9;
  LUT2 desc2606(.I0(acquisition_length[0:0]),.I1(window_length_fast[0:0]),.O(un18_m_axis_output_tready_cry_0_RNO));
defparam desc2606.INIT=4'h9;
  LUT2 desc2607(.I0(acquisition_length[1:1]),.I1(window_length[1:1]),.O(un18_m_axis_output_tready_axb_1));
defparam desc2607.INIT=4'h9;
  LUT2 desc2608(.I0(acquisition_length[2:2]),.I1(window_length[2:2]),.O(un18_m_axis_output_tready_axb_2));
defparam desc2608.INIT=4'h9;
  LUT2 desc2609(.I0(acquisition_length[3:3]),.I1(window_length[3:3]),.O(un18_m_axis_output_tready_axb_3));
defparam desc2609.INIT=4'h9;
  LUT2 desc2610(.I0(acquisition_length[4:4]),.I1(window_length[4:4]),.O(un18_m_axis_output_tready_axb_4));
defparam desc2610.INIT=4'h9;
  LUT2 desc2611(.I0(acquisition_length[5:5]),.I1(window_length[5:5]),.O(un18_m_axis_output_tready_axb_5));
defparam desc2611.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_1_cZ(.I0(acquisition_length[1:1]),.I1(window_length[1:1]),.O(un21_m_axis_output_tready_axb_1));
defparam un21_m_axis_output_tready_axb_1_cZ.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_2_cZ(.I0(acquisition_length[2:2]),.I1(window_length[2:2]),.O(un21_m_axis_output_tready_axb_2));
defparam un21_m_axis_output_tready_axb_2_cZ.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_3_cZ(.I0(acquisition_length[3:3]),.I1(window_length[3:3]),.O(un21_m_axis_output_tready_axb_3));
defparam un21_m_axis_output_tready_axb_3_cZ.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_4_cZ(.I0(acquisition_length[4:4]),.I1(window_length[4:4]),.O(un21_m_axis_output_tready_axb_4));
defparam un21_m_axis_output_tready_axb_4_cZ.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_5_cZ(.I0(acquisition_length[5:5]),.I1(window_length[5:5]),.O(un21_m_axis_output_tready_axb_5));
defparam un21_m_axis_output_tready_axb_5_cZ.INIT=4'h9;
  LUT4 read_ram_fsm_1_0_sqmuxa_1_scy_cZ(.I0(read_ram_fsm_1_0_rep1),.I1(read_ram_fsm_1_1_rep1),.I2(reorder_tvalid_fast[1:1]),.I3(traceback_tvalid[1:1]),.O(read_ram_fsm_1_0_sqmuxa_1_scy));
defparam read_ram_fsm_1_0_sqmuxa_1_scy_cZ.INIT=16'h0888;
  LUT2 desc2612(.I0(read_addr_ptr_1[6:6]),.I1(un21_m_axis_output_tready_s_6),.O(un57_m_axis_output_tready_0_N_3_i));
defparam desc2612.INIT=4'h9;
  LUT2 desc2613(.I0(read_addr_ptr_0[6:6]),.I1(un21_m_axis_output_tready_s_6),.O(un23_m_axis_output_tready_0_N_3_i));
defparam desc2613.INIT=4'h9;
  LUT2 desc2614(.I0(un64_m_axis_output_tready_a_5[6:6]),.I1(read_addr_ptr_1[6:6]),.O(un64_m_axis_output_tready_0_N_3_i));
defparam desc2614.INIT=4'h9;
  LUT2 desc2615(.I0(un18_m_axis_output_tready[6:6]),.I1(read_addr_ptr_0[6:6]),.O(un30_m_axis_output_tready_0_N_3_i));
defparam desc2615.INIT=4'h9;
  INV aresetn_i_c(.I(aresetn),.O(aresetn_i));
  FDR desc2616(.Q(ram_tlast[1:1]),.D(m_axis_output_tlast_int[1:1]),.C(aclk),.R(aresetn_i));
  FDR desc2617(.Q(ram_tlast[0:0]),.D(m_axis_output_tlast_int[0:0]),.C(aclk),.R(aresetn_i));
  FDR desc2618(.Q(ram_last_tuser[1:1]),.D(m_axis_output_last_tuser_int[1:1]),.C(aclk),.R(aresetn_i));
  FDR desc2619(.Q(ram_last_tuser[0:0]),.D(m_axis_output_last_tuser_int[0:0]),.C(aclk),.R(aresetn_i));
  FDR write_window_complete_Z(.Q(write_window_complete),.D(write_window_complete_0),.C(aclk),.R(aresetn_i));
  FDR write_last_window_complete_Z(.Q(write_last_window_complete),.D(write_last_window_complete_0),.C(aclk),.R(aresetn_i));
  FDE desc2620(.Q(window_length[0:0]),.D(s_axis_ctrl_tdata_16),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2621(.Q(window_length[1:1]),.D(s_axis_ctrl_tdata_17),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2622(.Q(window_length[2:2]),.D(s_axis_ctrl_tdata_18),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2623(.Q(window_length[3:3]),.D(s_axis_ctrl_tdata_19),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2624(.Q(window_length[4:4]),.D(s_axis_ctrl_tdata_20),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2625(.Q(window_length[5:5]),.D(s_axis_ctrl_tdata_21),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2626(.Q(window_length[6:6]),.D(s_axis_ctrl_tdata_22),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2627(.Q(acquisition_length[0:0]),.D(s_axis_ctrl_tdata_0),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2628(.Q(acquisition_length[1:1]),.D(s_axis_ctrl_tdata_1),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2629(.Q(acquisition_length[2:2]),.D(s_axis_ctrl_tdata_2),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2630(.Q(acquisition_length[3:3]),.D(s_axis_ctrl_tdata_3),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2631(.Q(acquisition_length[4:4]),.D(s_axis_ctrl_tdata_4),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2632(.Q(acquisition_length[5:5]),.D(s_axis_ctrl_tdata_5),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2633(.Q(acquisition_length[6:6]),.D(s_axis_ctrl_tdata_6),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FD desc2634(.Q(read_addr_ptr_0[0:0]),.D(un1_read_addr_ptr_0_2_axb_0),.C(aclk));
  FD desc2635(.Q(read_addr_ptr_0[1:1]),.D(un1_read_addr_ptr_0_2_s_1),.C(aclk));
  FD desc2636(.Q(read_addr_ptr_0[2:2]),.D(un1_read_addr_ptr_0_2_s_2),.C(aclk));
  FD desc2637(.Q(read_addr_ptr_0[3:3]),.D(un1_read_addr_ptr_0_2_s_3),.C(aclk));
  FD desc2638(.Q(read_addr_ptr_0[4:4]),.D(un1_read_addr_ptr_0_2_s_4),.C(aclk));
  FD desc2639(.Q(read_addr_ptr_0[5:5]),.D(un1_read_addr_ptr_0_2_s_5),.C(aclk));
  FD desc2640(.Q(read_addr_ptr_0[6:6]),.D(un1_read_addr_ptr_0_2_s_6),.C(aclk));
  FD desc2641(.Q(read_addr_ptr_1[0:0]),.D(un1_read_addr_ptr_1_2_axb_0),.C(aclk));
  FD desc2642(.Q(read_addr_ptr_1[1:1]),.D(un1_read_addr_ptr_1_2_s_1),.C(aclk));
  FD desc2643(.Q(read_addr_ptr_1[2:2]),.D(un1_read_addr_ptr_1_2_s_2),.C(aclk));
  FD desc2644(.Q(read_addr_ptr_1[3:3]),.D(un1_read_addr_ptr_1_2_s_3),.C(aclk));
  FD desc2645(.Q(read_addr_ptr_1[4:4]),.D(un1_read_addr_ptr_1_2_s_4),.C(aclk));
  FD desc2646(.Q(read_addr_ptr_1[5:5]),.D(un1_read_addr_ptr_1_2_s_5),.C(aclk));
  FD desc2647(.Q(read_addr_ptr_1[6:6]),.D(un1_read_addr_ptr_1_2_s_6),.C(aclk));
  FD desc2648(.Q(read_ram_ptr_0[0:0]),.D(read_ram_ptr_0_RNO),.C(aclk));
  FD desc2649(.Q(read_ram_ptr_0[1:1]),.D(un2_write_ram_ptr_3_iv_1_RNI880U2_O6),.C(aclk));
  FD desc2650(.Q(read_ram_ptr_1[0:0]),.D(read_ram_ptr_1_RNO),.C(aclk));
  FD desc2651(.Q(read_ram_ptr_1[1:1]),.D(un2_write_ram_ptr_2_iv_1_RNIGNT55_O6),.C(aclk));
  FD desc2652(.Q(ram_buffer_full[0:0]),.D(ram_buffer_full_nss[0:0]),.C(aclk));
  FD desc2653(.Q(ram_buffer_full[1:1]),.D(ram_buffer_full_nss[1:1]),.C(aclk));
  FD desc2654(.Q(next_traceback),.D(N_941s),.C(aclk));
  FD desc2655(.Q(read_ram_fsm_0[0:0]),.D(read_ram_fsm_0_nss[0:0]),.C(aclk));
  FD desc2656(.Q(read_ram_fsm_0[1:1]),.D(read_ram_fsm_0_nss[1:1]),.C(aclk));
  FD desc2657(.Q(read_ram_fsm_1[0:0]),.D(read_ram_fsm_1_nss[0:0]),.C(aclk));
  FD desc2658(.Q(read_ram_fsm_1[1:1]),.D(read_ram_fsm_1_nss[1:1]),.C(aclk));
  FDR last_of_block_Z(.Q(last_of_block),.D(last_of_block_0),.C(aclk),.R(aresetn_i));
  FDR desc2659(.Q(write_addr_ptr[0:0]),.D(N_1785),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2660(.Q(write_addr_ptr[1:1]),.D(N_1786),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2661(.Q(write_addr_ptr[2:2]),.D(N_1787),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2662(.Q(write_addr_ptr[3:3]),.D(N_1788),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2663(.Q(write_addr_ptr[4:4]),.D(N_1789),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2664(.Q(write_addr_ptr[5:5]),.D(N_1790),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FDR desc2665(.Q(write_addr_ptr[6:6]),.D(N_1791),.C(aclk),.R(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
  FD desc2666(.Q(wen_ram[0:0]),.D(wen_ramd_0[0:0]),.C(aclk));
  FD desc2667(.Q(wen_ram[1:1]),.D(wen_ramd_0[1:1]),.C(aclk));
  FD desc2668(.Q(wen_ram[2:2]),.D(wen_ramd_0[2:2]),.C(aclk));
  FD desc2669(.Q(wen_ram[3:3]),.D(wen_ramd_0[3:3]),.C(aclk));
  FD desc2670(.Q(read_ram_ptr_0_fast[0:0]),.D(N_425_fast),.C(aclk));
  FD desc2671(.Q(read_ram_ptr_0_fast[1:1]),.D(N_426_fast),.C(aclk));
  FDE desc2672(.Q(window_length_fast[0:0]),.D(s_axis_ctrl_tdata_16),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FD desc2673(.Q(read_ram_ptr_1_fast[1:1]),.D(N_430_fast),.C(aclk));
  FD desc2674(.Q(read_ram_ptr_1_fast[0:0]),.D(N_429_fast),.C(aclk));
  FDE desc2675(.Q(acquisition_length_fast),.D(s_axis_ctrl_tdata_0),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2676(.Q(window_length_fast[1:1]),.D(s_axis_ctrl_tdata_17),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2677(.Q(window_length_fast[2:2]),.D(s_axis_ctrl_tdata_18),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2678(.Q(window_length_fast[3:3]),.D(s_axis_ctrl_tdata_19),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FDE desc2679(.Q(window_length_fast[4:4]),.D(s_axis_ctrl_tdata_20),.C(aclk),.CE(wen_ram_0_sqmuxa_3));
  FD desc2680(.Q(read_ram_fsm_1_fast[1:1]),.D(read_ram_fsm_1_nss_fast[1:1]),.C(aclk));
  FD read_ram_fsm_1_1_rep1_Z(.Q(read_ram_fsm_1_1_rep1),.D(read_ram_fsm_1_nss_rep1[1:1]),.C(aclk));
  FD desc2681(.Q(read_ram_fsm_1_fast[0:0]),.D(read_ram_fsm_1_nss_fast[0:0]),.C(aclk));
  FD read_ram_fsm_1_0_rep1_Z(.Q(read_ram_fsm_1_0_rep1),.D(read_ram_fsm_1_nss_rep1[0:0]),.C(aclk));
  FD desc2682(.Q(read_ram_fsm_0_fast[0:0]),.D(read_ram_fsm_0_nss_fast[0:0]),.C(aclk));
  FD read_ram_fsm_0_0_rep1_Z(.Q(read_ram_fsm_0_0_rep1),.D(read_ram_fsm_0_nss_rep1[0:0]),.C(aclk));
  FD desc2683(.Q(read_ram_fsm_0_fast[1:1]),.D(read_ram_fsm_0_nss_fast[1:1]),.C(aclk));
  FD read_ram_fsm_0_1_rep1_Z(.Q(read_ram_fsm_0_1_rep1),.D(read_ram_fsm_0_nss_rep1[1:1]),.C(aclk));
  MUXCY desc2684(.DI(GND),.CI(un9_s_axis_input_tvalid_0_data_tmp[1:1]),.S(un9_s_axis_input_tvalid_0_I_19_RNO),.O(un9_s_axis_input_tvalid));
  MUXCY desc2685(.DI(GND),.CI(un30_m_axis_output_tready_0_data_tmp[1:1]),.S(un30_m_axis_output_tready_0_N_3_i),.O(un30_m_axis_output_tready));
  MUXCY desc2686(.DI(GND),.CI(un64_m_axis_output_tready_0_data_tmp[1:1]),.S(un64_m_axis_output_tready_0_N_3_i),.O(un64_m_axis_output_tready));
  MUXCY desc2687(.DI(GND),.CI(un23_m_axis_output_tready_0_data_tmp[1:1]),.S(un23_m_axis_output_tready_0_N_3_i),.O(un23_m_axis_output_tready));
  MUXCY desc2688(.DI(GND),.CI(un57_m_axis_output_tready_0_data_tmp[1:1]),.S(un57_m_axis_output_tready_0_N_3_i),.O(un57_m_axis_output_tready));
  LUT4 un1_write_ram_ptr_0_sqmuxa_cZ(.I0(acs_tvalid),.I1(write_ram_fsm_1),.I2(un1_write_ram_ptr_0_sqmuxa_sx),.I3(N_1756_1),.O(un1_write_ram_ptr_0_sqmuxa));
defparam un1_write_ram_ptr_0_sqmuxa_cZ.INIT=16'h0200;
  MUXCY read_ram_fsm_1_0_sqmuxa_1_cZ(.DI(GND),.CI(un64_m_axis_output_tready),.S(read_ram_fsm_1_0_sqmuxa_1_scy),.O(read_ram_fsm_1_0_sqmuxa_1));
  LUT5_L read_ram_fsm_0_1_rep1_RNO(.I0(aresetn),.I1(read_ram_fsm_0_1_rep1),.I2(read_ram_fsm_0[0:0]),.I3(read_ram_fsm_0_0_sqmuxa),.I4(N_54_mux),.LO(read_ram_fsm_0_nss_rep1[1:1]));
defparam read_ram_fsm_0_1_rep1_RNO.INIT=32'h2808A888;
  LUT5_L desc2689(.I0(aresetn),.I1(read_ram_fsm_0_fast[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(read_ram_fsm_0_0_sqmuxa),.I4(N_54_mux),.LO(read_ram_fsm_0_nss_fast[1:1]));
defparam desc2689.INIT=32'h2808A888;
  LUT6_L read_ram_fsm_0_0_rep1_RNO(.I0(aresetn),.I1(read_ram_fsm_0_0_rep1),.I2(read_ram_fsm_0[1:1]),.I3(un10_m_axis_output_tready),.I4(N_13_0),.I5(N_54_mux),.LO(read_ram_fsm_0_nss_rep1[0:0]));
defparam read_ram_fsm_0_0_rep1_RNO.INIT=64'h00200A2A80A08AAA;
  LUT6_L desc2690(.I0(aresetn),.I1(read_ram_fsm_0_fast[0:0]),.I2(read_ram_fsm_0[1:1]),.I3(un10_m_axis_output_tready),.I4(N_13_0),.I5(N_54_mux),.LO(read_ram_fsm_0_nss_fast[0:0]));
defparam desc2690.INIT=64'h00200A2A80A08AAA;
  LUT6_L read_ram_fsm_1_0_rep1_RNO(.I0(aresetn),.I1(read_ram_fsm_1_0_rep1),.I2(read_ram_fsm_1[1:1]),.I3(un44_m_axis_output_tready),.I4(N_13),.I5(N_54_mux_0),.LO(read_ram_fsm_1_nss_rep1[0:0]));
defparam read_ram_fsm_1_0_rep1_RNO.INIT=64'h00200A2A80A08AAA;
  LUT6_L desc2691(.I0(aresetn),.I1(read_ram_fsm_1_fast[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(un44_m_axis_output_tready),.I4(N_13),.I5(N_54_mux_0),.LO(read_ram_fsm_1_nss_fast[0:0]));
defparam desc2691.INIT=64'h00200A2A80A08AAA;
  LUT5_L read_ram_fsm_1_1_rep1_RNO(.I0(aresetn),.I1(read_ram_fsm_1_1_rep1),.I2(read_ram_fsm_1[0:0]),.I3(N_745),.I4(N_54_mux_0),.LO(read_ram_fsm_1_nss_rep1[1:1]));
defparam read_ram_fsm_1_1_rep1_RNO.INIT=32'h2808A888;
  LUT5_L desc2692(.I0(aresetn),.I1(read_ram_fsm_1_fast[1:1]),.I2(read_ram_fsm_1[0:0]),.I3(N_745),.I4(N_54_mux_0),.LO(read_ram_fsm_1_nss_fast[1:1]));
defparam desc2692.INIT=32'h2808A888;
  LUT6_L desc2693(.I0(aresetn),.I1(read_ram_ptr_1_fast[0:0]),.I2(write_ram_ptr[0:0]),.I3(N_1733),.I4(N_709),.I5(un2_write_ram_ptr_2_1[1:1]),.LO(N_429_fast));
defparam desc2693.INIT=64'h775F775588A0880A;
  LUT6_L desc2694(.I0(aresetn),.I1(read_ram_ptr_0_fast[0:0]),.I2(write_ram_ptr[0:0]),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(N_41_mux),.I5(un2_write_ram_ptr_3_1[1:1]),.LO(N_425_fast));
defparam desc2694.INIT=64'h7755775F880A88A0;
  LUT4 desc2695(.I0(read_ram_ptr_1_fast[1:1]),.I1(read_ram_ptr_1_fast[0:0]),.I2(write_ram_ptr_fast[0:0]),.I3(write_ram_ptr_fast[1:1]),.O(g5_0_0_0));
defparam desc2695.INIT=16'h7DBE;
  LUT4 desc2696(.I0(read_ram_ptr_0_fast[1:1]),.I1(read_ram_ptr_0_fast[0:0]),.I2(write_ram_ptr_fast[0:0]),.I3(write_ram_ptr_fast[1:1]),.O(g5_0_0));
defparam desc2696.INIT=16'h7DBE;
  LUT4 desc2697(.I0(read_ram_ptr_1[1:1]),.I1(read_ram_ptr_1[0:0]),.I2(write_ram_ptr[1:1]),.I3(write_ram_ptr[0:0]),.O(un3_s_axis_input_tready_int_li));
defparam desc2697.INIT=16'h7BDE;
  LUT6 desc2698(.I0(read_ram_fsm_0_fast[0:0]),.I1(read_ram_fsm_0_fast[1:1]),.I2(read_ram_fsm_1_fast[0:0]),.I3(read_ram_fsm_1_fast[1:1]),.I4(g5_0_0),.I5(g5_0_0_0),.O(N_1756_1));
defparam desc2698.INIT=64'hFFFF1111000F0001;
  LUT4 desc2699(.I0(read_ram_ptr_0[1:1]),.I1(read_ram_ptr_0[0:0]),.I2(write_ram_ptr[1:1]),.I3(write_ram_ptr[0:0]),.O(un15_s_axis_input_tready_int_li));
defparam desc2699.INIT=16'h7BDE;
  LUT4_L desc2700(.I0(wen_ram[0:0]),.I1(N_1872),.I2(un9_s_axis_input_tvalid_0_I_19_RNIN8NO),.I3(un1_wen_ram_1_sqmuxa_1_i),.LO(wen_ramd_0[0:0]));
defparam desc2700.INIT=16'h0C0A;
  LUT4_L desc2701(.I0(wen_ram[3:3]),.I1(N_1875),.I2(un9_s_axis_input_tvalid_0_I_19_RNIN8NO),.I3(un1_wen_ram_1_sqmuxa_1_i),.LO(wen_ramd_0[3:3]));
defparam desc2701.INIT=16'h0C0A;
  LUT4_L desc2702(.I0(wen_ram[2:2]),.I1(N_1874),.I2(un9_s_axis_input_tvalid_0_I_19_RNIN8NO),.I3(un1_wen_ram_1_sqmuxa_1_i),.LO(wen_ramd_0[2:2]));
defparam desc2702.INIT=16'h0C0A;
  LUT4_L desc2703(.I0(wen_ram[1:1]),.I1(N_1873),.I2(un9_s_axis_input_tvalid_0_I_19_RNIN8NO),.I3(un1_wen_ram_1_sqmuxa_1_i),.LO(wen_ramd_0[1:1]));
defparam desc2703.INIT=16'h0C0A;
  LUT5 desc2704(.I0(read_ram_fsm_0[1:1]),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(read_ram_fsm_0[0:0]),.I4(un9_s_axis_input_tvalid),.O(N_1747));
defparam desc2704.INIT=32'h0357FFFF;
  LUT6 desc2705(.I0(write_ram_fsm[3:3]),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(un3_s_axis_input_tready_int_li),.I5(un15_s_axis_input_tready_int_li),.O(write_ram_fsm_ns_0_a4_0_0[2:2]));
defparam desc2705.INIT=64'hAAAA020200AA0002;
  LUT6 desc2706(.I0(read_ram_fsm_1[0:0]),.I1(read_ram_fsm_1[1:1]),.I2(write_ram_fsm_ns_0_a4_2_1),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(un3_s_axis_input_tready_int_li),.I5(un15_s_axis_input_tready_int_li),.O(write_ram_fsm_ns_0_0[0:0]));
defparam desc2706.INIT=64'h10F0101000F00010;
  LUT6_L desc2707(.I0(acquisition_length[0:0]),.I1(window_length[0:0]),.I2(read_addr_ptr_1[0:0]),.I3(traceback_tvalid[1:1]),.I4(reorder_tvalid_1_rep1),.I5(m33_0_0),.LO(m33_0));
defparam desc2707.INIT=64'h0069696900000000;
  LUT6 desc2708(.I0(write_window_complete),.I1(write_last_window_complete),.I2(read_ram_fsm_0[0:0]),.I3(next_traceback),.I4(un10_m_axis_output_tready),.I5(read_ram_fsm_0_0_sqmuxa),.O(N_13_0));
defparam desc2708.INIT=64'hFFF10F010F010F01;
  LUT6 un1_read_ram_ptr_1_1_sqmuxa_0_cZ(.I0(read_ram_fsm_1_1_rep1),.I1(read_ram_fsm_1_0_rep1),.I2(write_window_complete),.I3(write_last_window_complete),.I4(next_traceback),.I5(un44_m_axis_output_tready),.O(un1_read_ram_ptr_1_1_sqmuxa_0));
defparam un1_read_ram_ptr_1_1_sqmuxa_0_cZ.INIT=64'h0001111122233333;
  LUT6 desc2709(.I0(traceback_tvalid[0:0]),.I1(reorder_tvalid_0_rep1),.I2(read_addr_ptr_0_1_sqmuxa_1),.I3(read_ram_fsm_0_2_sqmuxa_0),.I4(read_addr_ptr_0_1_sqmuxa_3),.I5(read_addr_ptr_0_2_sqmuxa_1),.O(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]));
defparam desc2709.INIT=64'hFFFFFFFFFFFFF7F0;
  LUT6 un1_read_addr_ptr_0_1_sqmuxa_1_1_cZ(.I0(traceback_tvalid[0:0]),.I1(reorder_tvalid_0_rep1),.I2(read_ram_fsm_0[1:1]),.I3(read_ram_fsm_0[0:0]),.I4(un10_m_axis_output_tready),.I5(un30_m_axis_output_tready),.O(un1_read_addr_ptr_0_1_sqmuxa_1_1));
defparam un1_read_addr_ptr_0_1_sqmuxa_1_1_cZ.INIT=64'h88F08800F8F0F800;
  LUT6 un1_read_addr_ptr_0_2_axb_4_RNO(.I0(aresetn),.I1(read_last_addr_ptr[4:4]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[4:4]));
defparam un1_read_addr_ptr_0_2_axb_4_RNO.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_1_2_axb_4_RNO(.I0(aresetn),.I1(read_last_addr_ptr[4:4]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[4:4]));
defparam un1_read_addr_ptr_1_2_axb_4_RNO.INIT=64'h0000008000000000;
  LUT6 desc2710(.I0(aresetn),.I1(read_last_addr_ptr[0:0]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[0:0]));
defparam desc2710.INIT=64'h0000008000000000;
  LUT6 desc2711(.I0(aresetn),.I1(read_last_addr_ptr[5:5]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[5:5]));
defparam desc2711.INIT=64'h0000008000000000;
  LUT6 desc2712(.I0(read_ram_fsm_0_0_rep1),.I1(read_ram_ptr_0[1:1]),.I2(read_ram_ptr_0[0:0]),.I3(write_window_complete),.I4(read_ram_fsm_0[1:1]),.I5(next_traceback),.O(un16_addr));
defparam desc2712.INIT=64'h0303020203030302;
  LUT6 desc2713(.I0(aresetn),.I1(read_last_addr_ptr[0:0]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[0:0]));
defparam desc2713.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_0_2_axb_1_RNO(.I0(aresetn),.I1(read_last_addr_ptr[1:1]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[1:1]));
defparam un1_read_addr_ptr_0_2_axb_1_RNO.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_0_2_axb_2_RNO(.I0(aresetn),.I1(read_last_addr_ptr[2:2]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[2:2]));
defparam un1_read_addr_ptr_0_2_axb_2_RNO.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_0_2_axb_3_RNO(.I0(aresetn),.I1(read_last_addr_ptr[3:3]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[3:3]));
defparam un1_read_addr_ptr_0_2_axb_3_RNO.INIT=64'h0000000000000080;
  LUT6 desc2714(.I0(aresetn),.I1(read_last_addr_ptr[5:5]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[5:5]));
defparam desc2714.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_0_2_axb_6_RNO(.I0(aresetn),.I1(read_last_addr_ptr[6:6]),.I2(write_last_window_complete),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(read_last_addr_ptr_m[6:6]));
defparam un1_read_addr_ptr_0_2_axb_6_RNO.INIT=64'h0000000000000080;
  LUT6 un1_read_addr_ptr_1_2_axb_1_RNO(.I0(aresetn),.I1(read_last_addr_ptr[1:1]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[1:1]));
defparam un1_read_addr_ptr_1_2_axb_1_RNO.INIT=64'h0000008000000000;
  LUT6 un1_read_addr_ptr_1_2_axb_2_RNO(.I0(aresetn),.I1(read_last_addr_ptr[2:2]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[2:2]));
defparam un1_read_addr_ptr_1_2_axb_2_RNO.INIT=64'h0000008000000000;
  LUT6 un1_read_addr_ptr_1_2_axb_3_RNO(.I0(aresetn),.I1(read_last_addr_ptr[3:3]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[3:3]));
defparam un1_read_addr_ptr_1_2_axb_3_RNO.INIT=64'h0000008000000000;
  LUT6 un1_read_addr_ptr_1_2_axb_6_RNO(.I0(aresetn),.I1(read_last_addr_ptr[6:6]),.I2(write_last_window_complete),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(next_traceback),.O(read_last_addr_ptr_m_0[6:6]));
defparam un1_read_addr_ptr_1_2_axb_6_RNO.INIT=64'h0000008000000000;
  LUT6 desc2715(.I0(read_ram_fsm_0_1_rep1),.I1(read_ram_ptr_0[1:1]),.I2(read_ram_ptr_0[0:0]),.I3(write_window_complete),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(un87_addr));
defparam desc2715.INIT=64'h0C0C08080C0C0C08;
  LUT6 desc2716(.I0(read_ram_fsm_0_1_rep1),.I1(read_ram_ptr_0[1:1]),.I2(read_ram_ptr_0[0:0]),.I3(write_window_complete),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(un55_addr));
defparam desc2716.INIT=64'h3030202030303020;
  LUT6 desc2717(.I0(read_ram_fsm_0_1_rep1),.I1(read_ram_ptr_0[1:1]),.I2(read_ram_ptr_0[0:0]),.I3(write_window_complete),.I4(read_ram_fsm_0[0:0]),.I5(next_traceback),.O(un119_addr));
defparam desc2717.INIT=64'hC0C08080C0C0C080;
  LUT5 m_axis_output_tlast_int_0_sqmuxa_1_1_cZ(.I0(last_of_block),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep1),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.O(m_axis_output_tlast_int_0_sqmuxa_1_1));
defparam m_axis_output_tlast_int_0_sqmuxa_1_1_cZ.INIT=32'h0000002A;
  LUT5 desc2718(.I0(aresetn),.I1(write_last_window_complete),.I2(read_ram_fsm_1[0:0]),.I3(read_ram_fsm_1[1:1]),.I4(next_traceback),.O(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]));
defparam desc2718.INIT=32'hAAA2AAAA;
  LUT6 read_addr_ptr_0_1_sqmuxa_3_cZ(.I0(ram_tvalid[0:0]),.I1(traceback_tvalid[0:0]),.I2(reorder_tvalid_0_rep1),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(un30_m_axis_output_tready),.O(read_addr_ptr_0_1_sqmuxa_3));
defparam read_addr_ptr_0_1_sqmuxa_3_cZ.INIT=64'h400000007F000000;
  LUT6_L desc2719(.I0(ram_last_tuser[0:0]),.I1(traceback_tvalid[0:0]),.I2(reorder_tvalid_0_rep1),.I3(read_ram_fsm_0[1:1]),.I4(read_ram_fsm_0[0:0]),.I5(un30_m_axis_output_tready),.LO(m_axis_output_last_tuser_int[0:0]));
defparam desc2719.INIT=64'hBF00AA00AA00AA00;
  LUT6 desc2720(.I0(acs_tlast),.I1(read_ram_ptr_0[1:1]),.I2(read_ram_ptr_0[0:0]),.I3(write_ram_fsm[2:2]),.I4(write_ram_ptr[1:1]),.I5(write_ram_ptr[0:0]),.O(write_ram_fsm_ns_i_o4_0_0[3:3]));
defparam desc2720.INIT=64'hEAFFBAFFAEFFABFF;
  LUT5_L desc2721(.I0(aresetn),.I1(ram_tvalid[0:0]),.I2(traceback_tvalid[0:0]),.I3(ram_buffer_full[0:0]),.I4(reorder_tvalid_0_rep2),.LO(ram_buffer_full_nss[0:0]));
defparam desc2721.INIT=32'hA2802200;
  LUT4 desc2722(.I0(ram_tvalid[0:0]),.I1(traceback_tvalid[0:0]),.I2(reorder_tvalid_0_rep1),.I3(ram_buffer_full[0:0]),.O(un5_m_axis_output_tvalid_int));
defparam desc2722.INIT=16'h0080;
  LUT5 un1_read_addr_ptr_0_1_sqmuxa_1_1_RNIVUDO(.I0(aresetn),.I1(read_addr_ptr_0[5:5]),.I2(read_addr_ptr_0_1_sqmuxa_1),.I3(read_ram_fsm_0_2_sqmuxa_0),.I4(un1_read_addr_ptr_0_1_sqmuxa_1_1),.O(read_addr_ptr_0_m[5:5]));
defparam un1_read_addr_ptr_0_1_sqmuxa_1_1_RNIVUDO.INIT=32'h88888880;
  LUT6 read_addr_ptr_0_1_sqmuxa_3_RNIVHT32_cZ(.I0(N_99),.I1(read_addr_ptr_0_1_sqmuxa_1),.I2(read_ram_fsm_0_2_sqmuxa_0),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(read_addr_ptr_0_1_sqmuxa_3),.I5(read_addr_ptr_0_2_sqmuxa_1),.O(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32));
defparam read_addr_ptr_0_1_sqmuxa_3_RNIVHT32_cZ.INIT=64'hFF00FF00FF00DC00;
  LUT4 read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ_cZ(.I0(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I1(un1_read_addr_ptr_1_1_sqmuxa_0),.I2(read_addr_ptr_1_2_sqmuxa_1),.I3(read_addr_ptr_1_1_sqmuxa_3),.O(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ));
defparam read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ_cZ.INIT=16'hAAA8;
  LUT6_L read_addr_ptr_0_2_sqmuxa_1_RNI630O2(.I0(window_length[5:5]),.I1(read_last_addr_ptr_m[5:5]),.I2(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I3(read_addr_ptr_0_2_sqmuxa_1),.I4(read_addr_ptr_0_m[5:5]),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_5));
defparam read_addr_ptr_0_2_sqmuxa_1_RNI630O2.INIT=64'h0F0F1E3CFFFFEECC;
  LUT6_L un1_read_addr_ptr_1_2_axb_0_cZ(.I0(window_length[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(read_last_addr_ptr_m_0[0:0]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_0));
defparam un1_read_addr_ptr_1_2_axb_0_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_1_2_axb_1_cZ(.I0(window_length[1:1]),.I1(read_addr_ptr_1[1:1]),.I2(read_last_addr_ptr_m_0[1:1]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_1));
defparam un1_read_addr_ptr_1_2_axb_1_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6 un1_read_addr_ptr_1_2_cry_0_RNO_cZ(.I0(window_length[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(read_last_addr_ptr_m_0[0:0]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.O(un1_read_addr_ptr_1_2_cry_0_RNO));
defparam un1_read_addr_ptr_1_2_cry_0_RNO_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_1_2_axb_3_cZ(.I0(window_length[3:3]),.I1(read_addr_ptr_1[3:3]),.I2(read_last_addr_ptr_m_0[3:3]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_3));
defparam un1_read_addr_ptr_1_2_axb_3_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_1_2_axb_4_cZ(.I0(window_length[4:4]),.I1(read_addr_ptr_1[4:4]),.I2(read_last_addr_ptr_m_0[4:4]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_4));
defparam un1_read_addr_ptr_1_2_axb_4_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_1_2_axb_6_cZ(.I0(window_length[6:6]),.I1(read_addr_ptr_1[6:6]),.I2(read_last_addr_ptr_m_0[6:6]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_6));
defparam un1_read_addr_ptr_1_2_axb_6_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_1_2_axb_2_cZ(.I0(window_length[2:2]),.I1(read_addr_ptr_1[2:2]),.I2(read_last_addr_ptr_m_0[2:2]),.I3(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_4),.I5(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_2));
defparam un1_read_addr_ptr_1_2_axb_2_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_0_cZ(.I0(window_length[0:0]),.I1(read_addr_ptr_0[0:0]),.I2(read_last_addr_ptr_m[0:0]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_0));
defparam un1_read_addr_ptr_0_2_axb_0_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_4_cZ(.I0(window_length[4:4]),.I1(read_addr_ptr_0[4:4]),.I2(read_last_addr_ptr_m[4:4]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_4));
defparam un1_read_addr_ptr_0_2_axb_4_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_6_cZ(.I0(window_length[6:6]),.I1(read_addr_ptr_0[6:6]),.I2(read_last_addr_ptr_m[6:6]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_6));
defparam un1_read_addr_ptr_0_2_axb_6_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6 un1_read_addr_ptr_0_2_cry_0_RNO_cZ(.I0(window_length[0:0]),.I1(read_addr_ptr_0[0:0]),.I2(read_last_addr_ptr_m[0:0]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.O(un1_read_addr_ptr_0_2_cry_0_RNO));
defparam un1_read_addr_ptr_0_2_cry_0_RNO_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_1_cZ(.I0(window_length[1:1]),.I1(read_addr_ptr_0[1:1]),.I2(read_last_addr_ptr_m[1:1]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_1));
defparam un1_read_addr_ptr_0_2_axb_1_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_2_cZ(.I0(window_length[2:2]),.I1(read_addr_ptr_0[2:2]),.I2(read_last_addr_ptr_m[2:2]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_2));
defparam un1_read_addr_ptr_0_2_axb_2_cZ.INIT=64'h03FC05F0FCFCF0F0;
  LUT6_L un1_read_addr_ptr_0_2_axb_3_cZ(.I0(window_length[3:3]),.I1(read_addr_ptr_0[3:3]),.I2(read_last_addr_ptr_m[3:3]),.I3(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]),.I4(un1_ram_buffer_05_5),.I5(un1_read_addr_ptr_0_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_0_2_axb_3));
defparam un1_read_addr_ptr_0_2_axb_3_cZ.INIT=64'h03FC05F0FCFCF0F0;
  MUXCY_L un1_write_addr_ptr_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(wen_ram_0_sqmuxa_3),.LO(un1_write_addr_ptr_cry_0_cy));
  MUXCY_L un1_write_addr_ptr_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(wen_ram_0_sqmuxa_3_ci),.LO(un1_write_addr_ptr_0_cry_0_cy));
  LUT6 wen_ram_0_sqmuxa_3_ci_cZ(.I0(aresetn),.I1(s_axis_ctrl_tvalid),.I2(write_ram_fsm_4_rep1),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(read_ram_fsm_0_d_i_0[3:3]),.O(wen_ram_0_sqmuxa_3_ci));
defparam wen_ram_0_sqmuxa_3_ci_cZ.INIT=64'h0000000000000080;
  LUT4 un1_ram_buffer_05_5_cZ(.I0(aresetn),.I1(read_addr_ptr_0_1_sqmuxa_1),.I2(read_ram_fsm_0_2_sqmuxa_0),.I3(un1_read_addr_ptr_0_1_sqmuxa_1_1),.O(un1_ram_buffer_05_5));
defparam un1_ram_buffer_05_5_cZ.INIT=16'hAAA8;
  LUT5 un9_s_axis_ctrl_tready_int(.I0(read_ram_fsm_0[0:0]),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_1[0:0]),.I3(read_ram_fsm_1[1:1]),.I4(write_ram_fsm_4),.O(s_axis_ctrl_tready));
defparam un9_s_axis_ctrl_tready_int.INIT=32'h00010000;
  LUT2_L read_ram_fsm_1_2_sqmuxa_i_a2_0_cZ(.I0(read_addr_ptr_1[3:3]),.I1(read_addr_ptr_1[4:4]),.LO(read_ram_fsm_1_2_sqmuxa_i_a2_0));
defparam read_ram_fsm_1_2_sqmuxa_i_a2_0_cZ.INIT=4'h1;
  LUT2 un21_m_axis_output_tready_axb_6_cZ(.I0(acquisition_length[6:6]),.I1(window_length[6:6]),.O(un21_m_axis_output_tready_axb_6));
defparam un21_m_axis_output_tready_axb_6_cZ.INIT=4'h9;
  LUT2 un21_m_axis_output_tready_axb_0_cZ(.I0(acquisition_length[0:0]),.I1(window_length[0:0]),.O(un21_m_axis_output_tready_axb_0));
defparam un21_m_axis_output_tready_axb_0_cZ.INIT=4'h9;
  LUT2 desc2723(.I0(acquisition_length[6:6]),.I1(window_length[6:6]),.O(un18_m_axis_output_tready_axb_6));
defparam desc2723.INIT=4'h9;
  LUT2 desc2724(.I0(acquisition_length[6:6]),.I1(window_length[6:6]),.O(un64_m_axis_output_tready_a_5_axb_6));
defparam desc2724.INIT=4'h9;
  LUT4 desc2725(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_0[2:2]),.I2(un18_m_axis_output_tready[2:2]),.I3(un18_m_axis_output_tready[3:3]),.O(m33_1));
defparam desc2725.INIT=16'h8241;
  LUT4 desc2726(.I0(read_addr_ptr_1[5:5]),.I1(read_addr_ptr_1[6:6]),.I2(un18_m_axis_output_tready[5:5]),.I3(un18_m_axis_output_tready[6:6]),.O(m33_0_2));
defparam desc2726.INIT=16'h8421;
  LUT4_L desc2727(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_1[2:2]),.I2(un18_m_axis_output_tready[1:1]),.I3(un18_m_axis_output_tready[2:2]),.LO(m33_0_0));
defparam desc2727.INIT=16'h8421;
  LUT4 desc2728(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_0[4:4]),.I2(read_addr_ptr_0[5:5]),.I3(read_addr_ptr_0[6:6]),.O(un6_m_axis_output_tready_3));
defparam desc2728.INIT=16'h0001;
  LUT4 desc2729(.I0(acs_tlast),.I1(write_ram_fsm[2:2]),.I2(write_window_complete),.I3(acs_tvalid),.O(write_ram_fsm_ns_0_a4_2_1));
defparam desc2729.INIT=16'h0800;
  LUT3 desc2730(.I0(acquisition_length[0:0]),.I1(window_length[0:0]),.I2(read_addr_ptr_0[0:0]),.O(un30_m_axis_output_tready_0_N_14));
defparam desc2730.INIT=8'h96;
  LUT6 desc2731(.I0(read_ram_ptr_1[1:1]),.I1(read_ram_ptr_1[0:0]),.I2(read_ram_fsm_1_1_rep1),.I3(read_ram_ptr_0[1:1]),.I4(read_ram_fsm_1_0_rep1),.I5(read_ram_ptr_0[0:0]),.O(un10_m_axis_output_tready));
defparam desc2731.INIT=64'h0201000004080000;
  LUT6 desc2732(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_1[2:2]),.I2(read_addr_ptr_1[0:0]),.I3(un64_m_axis_output_tready_a_5_axb_0),.I4(un64_m_axis_output_tready_a_5[1:1]),.I5(un64_m_axis_output_tready_a_5[2:2]),.O(un64_m_axis_output_tready_0_N_11));
defparam desc2732.INIT=64'h0880044002200110;
  LUT6 read_ram_fsm_1_2_sqmuxa_i_a2(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_1[2:2]),.I2(read_addr_ptr_1[5:5]),.I3(read_addr_ptr_1[6:6]),.I4(read_addr_ptr_1[0:0]),.I5(read_ram_fsm_1_2_sqmuxa_i_a2_0),.O(N_743));
defparam read_ram_fsm_1_2_sqmuxa_i_a2.INIT=64'h0000000100000000;
  LUT6 desc2733(.I0(read_addr_ptr_1[3:3]),.I1(read_addr_ptr_1[4:4]),.I2(read_addr_ptr_1[5:5]),.I3(un21_m_axis_output_tready_s_3),.I4(un21_m_axis_output_tready_s_4),.I5(un21_m_axis_output_tready_s_5),.O(un57_m_axis_output_tready_0_N_4));
defparam desc2733.INIT=64'h8040201008040201;
  LUT6 desc2734(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_0[4:4]),.I2(read_addr_ptr_0[5:5]),.I3(un21_m_axis_output_tready_s_3),.I4(un21_m_axis_output_tready_s_4),.I5(un21_m_axis_output_tready_s_5),.O(un23_m_axis_output_tready_0_N_4));
defparam desc2734.INIT=64'h8040201008040201;
  LUT6 desc2735(.I0(read_addr_ptr_1[3:3]),.I1(read_addr_ptr_1[4:4]),.I2(read_addr_ptr_1[5:5]),.I3(un64_m_axis_output_tready_a_5[3:3]),.I4(un64_m_axis_output_tready_a_5[4:4]),.I5(un64_m_axis_output_tready_a_5[5:5]),.O(un64_m_axis_output_tready_0_N_4));
defparam desc2735.INIT=64'h8040201008040201;
  LUT5 desc2736(.I0(s_axis_ctrl_tvalid),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_1[0:0]),.I3(read_ram_fsm_1[1:1]),.I4(read_ram_fsm_0[0:0]),.O(N_1743));
defparam desc2736.INIT=32'hFFFFFFFD;
  LUT6 desc2737(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_0[4:4]),.I2(read_addr_ptr_0[5:5]),.I3(un18_m_axis_output_tready[3:3]),.I4(un18_m_axis_output_tready[4:4]),.I5(un18_m_axis_output_tready[5:5]),.O(un30_m_axis_output_tready_0_N_4));
defparam desc2737.INIT=64'h8040201008040201;
  LUT6 desc2738(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[0:0]),.I3(q_reg_1[0:0]),.I4(q_reg_2[0:0]),.I5(q_reg_3[0:0]),.O(ram_buffer_1_1[0:0]));
defparam desc2738.INIT=64'hFEDCBA9876543210;
  LUT6 desc2739(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[0:0]),.I3(q_reg_1[0:0]),.I4(q_reg_2[0:0]),.I5(q_reg_3[0:0]),.O(ram_buffer_0_2[0:0]));
defparam desc2739.INIT=64'hFEDCBA9876543210;
  LUT6 desc2740(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[1:1]),.I3(q_reg_1[1:1]),.I4(q_reg_2[1:1]),.I5(q_reg_3[1:1]),.O(ram_buffer_1_1[1:1]));
defparam desc2740.INIT=64'hFEDCBA9876543210;
  LUT6 desc2741(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[1:1]),.I3(q_reg_1[1:1]),.I4(q_reg_2[1:1]),.I5(q_reg_3[1:1]),.O(ram_buffer_0_2[1:1]));
defparam desc2741.INIT=64'hFEDCBA9876543210;
  LUT6 desc2742(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[2:2]),.I3(q_reg_1[2:2]),.I4(q_reg_2[2:2]),.I5(q_reg_3[2:2]),.O(ram_buffer_1_1[2:2]));
defparam desc2742.INIT=64'hFEDCBA9876543210;
  LUT6 desc2743(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[2:2]),.I3(q_reg_1[2:2]),.I4(q_reg_2[2:2]),.I5(q_reg_3[2:2]),.O(ram_buffer_0_2[2:2]));
defparam desc2743.INIT=64'hFEDCBA9876543210;
  LUT6 desc2744(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[3:3]),.I3(q_reg_1[3:3]),.I4(q_reg_2[3:3]),.I5(q_reg_3[3:3]),.O(ram_buffer_1_1[3:3]));
defparam desc2744.INIT=64'hFEDCBA9876543210;
  LUT6 desc2745(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[3:3]),.I3(q_reg_1[3:3]),.I4(q_reg_2[3:3]),.I5(q_reg_3[3:3]),.O(ram_buffer_0_2[3:3]));
defparam desc2745.INIT=64'hFEDCBA9876543210;
  LUT6 desc2746(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[4:4]),.I3(q_reg_1[4:4]),.I4(q_reg_2[4:4]),.I5(q_reg_3[4:4]),.O(ram_buffer_1_1[4:4]));
defparam desc2746.INIT=64'hFEDCBA9876543210;
  LUT6 desc2747(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[4:4]),.I3(q_reg_1[4:4]),.I4(q_reg_2[4:4]),.I5(q_reg_3[4:4]),.O(ram_buffer_0_2[4:4]));
defparam desc2747.INIT=64'hFEDCBA9876543210;
  LUT6 desc2748(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[5:5]),.I3(q_reg_1[5:5]),.I4(q_reg_2[5:5]),.I5(q_reg_3[5:5]),.O(ram_buffer_1_1[5:5]));
defparam desc2748.INIT=64'hFEDCBA9876543210;
  LUT6 desc2749(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[5:5]),.I3(q_reg_1[5:5]),.I4(q_reg_2[5:5]),.I5(q_reg_3[5:5]),.O(ram_buffer_0_2[5:5]));
defparam desc2749.INIT=64'hFEDCBA9876543210;
  LUT6 desc2750(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[6:6]),.I3(q_reg_1[6:6]),.I4(q_reg_2[6:6]),.I5(q_reg_3[6:6]),.O(ram_buffer_1_1[6:6]));
defparam desc2750.INIT=64'hFEDCBA9876543210;
  LUT6 desc2751(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[6:6]),.I3(q_reg_1[6:6]),.I4(q_reg_2[6:6]),.I5(q_reg_3[6:6]),.O(ram_buffer_0_2[6:6]));
defparam desc2751.INIT=64'hFEDCBA9876543210;
  LUT6 desc2752(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[7:7]),.I3(q_reg_1[7:7]),.I4(q_reg_2[7:7]),.I5(q_reg_3[7:7]),.O(ram_buffer_1_1[7:7]));
defparam desc2752.INIT=64'hFEDCBA9876543210;
  LUT6 desc2753(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[7:7]),.I3(q_reg_1[7:7]),.I4(q_reg_2[7:7]),.I5(q_reg_3[7:7]),.O(ram_buffer_0_2[7:7]));
defparam desc2753.INIT=64'hFEDCBA9876543210;
  LUT6 desc2754(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[8:8]),.I3(q_reg_1[8:8]),.I4(q_reg_2[8:8]),.I5(q_reg_3[8:8]),.O(ram_buffer_1_1[8:8]));
defparam desc2754.INIT=64'hFEDCBA9876543210;
  LUT6 desc2755(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[8:8]),.I3(q_reg_1[8:8]),.I4(q_reg_2[8:8]),.I5(q_reg_3[8:8]),.O(ram_buffer_0_2[8:8]));
defparam desc2755.INIT=64'hFEDCBA9876543210;
  LUT6 desc2756(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[9:9]),.I3(q_reg_1[9:9]),.I4(q_reg_2[9:9]),.I5(q_reg_3[9:9]),.O(ram_buffer_1_1[9:9]));
defparam desc2756.INIT=64'hFEDCBA9876543210;
  LUT6 desc2757(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[9:9]),.I3(q_reg_1[9:9]),.I4(q_reg_2[9:9]),.I5(q_reg_3[9:9]),.O(ram_buffer_0_2[9:9]));
defparam desc2757.INIT=64'hFEDCBA9876543210;
  LUT6 desc2758(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[10:10]),.I3(q_reg_1[10:10]),.I4(q_reg_2[10:10]),.I5(q_reg_3[10:10]),.O(ram_buffer_1_1[10:10]));
defparam desc2758.INIT=64'hFEDCBA9876543210;
  LUT6 desc2759(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[10:10]),.I3(q_reg_1[10:10]),.I4(q_reg_2[10:10]),.I5(q_reg_3[10:10]),.O(ram_buffer_0_2[10:10]));
defparam desc2759.INIT=64'hFEDCBA9876543210;
  LUT6 desc2760(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[11:11]),.I3(q_reg_1[11:11]),.I4(q_reg_2[11:11]),.I5(q_reg_3[11:11]),.O(ram_buffer_1_1[11:11]));
defparam desc2760.INIT=64'hFEDCBA9876543210;
  LUT6 desc2761(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[11:11]),.I3(q_reg_1[11:11]),.I4(q_reg_2[11:11]),.I5(q_reg_3[11:11]),.O(ram_buffer_0_2[11:11]));
defparam desc2761.INIT=64'hFEDCBA9876543210;
  LUT6 desc2762(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[12:12]),.I3(q_reg_1[12:12]),.I4(q_reg_2[12:12]),.I5(q_reg_3[12:12]),.O(ram_buffer_1_1[12:12]));
defparam desc2762.INIT=64'hFEDCBA9876543210;
  LUT6 desc2763(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[12:12]),.I3(q_reg_1[12:12]),.I4(q_reg_2[12:12]),.I5(q_reg_3[12:12]),.O(ram_buffer_0_2[12:12]));
defparam desc2763.INIT=64'hFEDCBA9876543210;
  LUT6 desc2764(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[13:13]),.I3(q_reg_1[13:13]),.I4(q_reg_2[13:13]),.I5(q_reg_3[13:13]),.O(ram_buffer_1_1[13:13]));
defparam desc2764.INIT=64'hFEDCBA9876543210;
  LUT6 desc2765(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[13:13]),.I3(q_reg_1[13:13]),.I4(q_reg_2[13:13]),.I5(q_reg_3[13:13]),.O(ram_buffer_0_2[13:13]));
defparam desc2765.INIT=64'hFEDCBA9876543210;
  LUT6 desc2766(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[14:14]),.I3(q_reg_1[14:14]),.I4(q_reg_2[14:14]),.I5(q_reg_3[14:14]),.O(ram_buffer_1_1[14:14]));
defparam desc2766.INIT=64'hFEDCBA9876543210;
  LUT6 desc2767(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[14:14]),.I3(q_reg_1[14:14]),.I4(q_reg_2[14:14]),.I5(q_reg_3[14:14]),.O(ram_buffer_0_2[14:14]));
defparam desc2767.INIT=64'hFEDCBA9876543210;
  LUT6 desc2768(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[15:15]),.I3(q_reg_1[15:15]),.I4(q_reg_2[15:15]),.I5(q_reg_3[15:15]),.O(ram_buffer_1_1[15:15]));
defparam desc2768.INIT=64'hFEDCBA9876543210;
  LUT6 desc2769(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[15:15]),.I3(q_reg_1[15:15]),.I4(q_reg_2[15:15]),.I5(q_reg_3[15:15]),.O(ram_buffer_0_2[15:15]));
defparam desc2769.INIT=64'hFEDCBA9876543210;
  LUT6 desc2770(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[16:16]),.I3(q_reg_1[16:16]),.I4(q_reg_2[16:16]),.I5(q_reg_3[16:16]),.O(ram_buffer_1_1[16:16]));
defparam desc2770.INIT=64'hFEDCBA9876543210;
  LUT6 desc2771(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[16:16]),.I3(q_reg_1[16:16]),.I4(q_reg_2[16:16]),.I5(q_reg_3[16:16]),.O(ram_buffer_0_2[16:16]));
defparam desc2771.INIT=64'hFEDCBA9876543210;
  LUT6 desc2772(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[17:17]),.I3(q_reg_1[17:17]),.I4(q_reg_2[17:17]),.I5(q_reg_3[17:17]),.O(ram_buffer_1_1[17:17]));
defparam desc2772.INIT=64'hFEDCBA9876543210;
  LUT6 desc2773(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[17:17]),.I3(q_reg_1[17:17]),.I4(q_reg_2[17:17]),.I5(q_reg_3[17:17]),.O(ram_buffer_0_2[17:17]));
defparam desc2773.INIT=64'hFEDCBA9876543210;
  LUT6 desc2774(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[18:18]),.I3(q_reg_1[18:18]),.I4(q_reg_2[18:18]),.I5(q_reg_3[18:18]),.O(ram_buffer_1_1[18:18]));
defparam desc2774.INIT=64'hFEDCBA9876543210;
  LUT6 desc2775(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[18:18]),.I3(q_reg_1[18:18]),.I4(q_reg_2[18:18]),.I5(q_reg_3[18:18]),.O(ram_buffer_0_2[18:18]));
defparam desc2775.INIT=64'hFEDCBA9876543210;
  LUT6 desc2776(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[19:19]),.I3(q_reg_1[19:19]),.I4(q_reg_2[19:19]),.I5(q_reg_3[19:19]),.O(ram_buffer_1_1[19:19]));
defparam desc2776.INIT=64'hFEDCBA9876543210;
  LUT6 desc2777(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[19:19]),.I3(q_reg_1[19:19]),.I4(q_reg_2[19:19]),.I5(q_reg_3[19:19]),.O(ram_buffer_0_2[19:19]));
defparam desc2777.INIT=64'hFEDCBA9876543210;
  LUT6 desc2778(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[20:20]),.I3(q_reg_1[20:20]),.I4(q_reg_2[20:20]),.I5(q_reg_3[20:20]),.O(ram_buffer_1_1[20:20]));
defparam desc2778.INIT=64'hFEDCBA9876543210;
  LUT6 desc2779(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[20:20]),.I3(q_reg_1[20:20]),.I4(q_reg_2[20:20]),.I5(q_reg_3[20:20]),.O(ram_buffer_0_2[20:20]));
defparam desc2779.INIT=64'hFEDCBA9876543210;
  LUT6 desc2780(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[21:21]),.I3(q_reg_1[21:21]),.I4(q_reg_2[21:21]),.I5(q_reg_3[21:21]),.O(ram_buffer_1_1[21:21]));
defparam desc2780.INIT=64'hFEDCBA9876543210;
  LUT6 desc2781(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[21:21]),.I3(q_reg_1[21:21]),.I4(q_reg_2[21:21]),.I5(q_reg_3[21:21]),.O(ram_buffer_0_2[21:21]));
defparam desc2781.INIT=64'hFEDCBA9876543210;
  LUT6 desc2782(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[22:22]),.I3(q_reg_1[22:22]),.I4(q_reg_2[22:22]),.I5(q_reg_3[22:22]),.O(ram_buffer_1_1[22:22]));
defparam desc2782.INIT=64'hFEDCBA9876543210;
  LUT6 desc2783(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[22:22]),.I3(q_reg_1[22:22]),.I4(q_reg_2[22:22]),.I5(q_reg_3[22:22]),.O(ram_buffer_0_2[22:22]));
defparam desc2783.INIT=64'hFEDCBA9876543210;
  LUT6 desc2784(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[23:23]),.I3(q_reg_1[23:23]),.I4(q_reg_2[23:23]),.I5(q_reg_3[23:23]),.O(ram_buffer_1_1[23:23]));
defparam desc2784.INIT=64'hFEDCBA9876543210;
  LUT6 desc2785(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[23:23]),.I3(q_reg_1[23:23]),.I4(q_reg_2[23:23]),.I5(q_reg_3[23:23]),.O(ram_buffer_0_2[23:23]));
defparam desc2785.INIT=64'hFEDCBA9876543210;
  LUT6 desc2786(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[24:24]),.I3(q_reg_1[24:24]),.I4(q_reg_2[24:24]),.I5(q_reg_3[24:24]),.O(ram_buffer_1_1[24:24]));
defparam desc2786.INIT=64'hFEDCBA9876543210;
  LUT6 desc2787(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[24:24]),.I3(q_reg_1[24:24]),.I4(q_reg_2[24:24]),.I5(q_reg_3[24:24]),.O(ram_buffer_0_2[24:24]));
defparam desc2787.INIT=64'hFEDCBA9876543210;
  LUT6 desc2788(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[25:25]),.I3(q_reg_1[25:25]),.I4(q_reg_2[25:25]),.I5(q_reg_3[25:25]),.O(ram_buffer_1_1[25:25]));
defparam desc2788.INIT=64'hFEDCBA9876543210;
  LUT6 desc2789(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[25:25]),.I3(q_reg_1[25:25]),.I4(q_reg_2[25:25]),.I5(q_reg_3[25:25]),.O(ram_buffer_0_2[25:25]));
defparam desc2789.INIT=64'hFEDCBA9876543210;
  LUT6 desc2790(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[26:26]),.I3(q_reg_1[26:26]),.I4(q_reg_2[26:26]),.I5(q_reg_3[26:26]),.O(ram_buffer_1_1[26:26]));
defparam desc2790.INIT=64'hFEDCBA9876543210;
  LUT6 desc2791(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[26:26]),.I3(q_reg_1[26:26]),.I4(q_reg_2[26:26]),.I5(q_reg_3[26:26]),.O(ram_buffer_0_2[26:26]));
defparam desc2791.INIT=64'hFEDCBA9876543210;
  LUT6 desc2792(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[27:27]),.I3(q_reg_1[27:27]),.I4(q_reg_2[27:27]),.I5(q_reg_3[27:27]),.O(ram_buffer_1_1[27:27]));
defparam desc2792.INIT=64'hFEDCBA9876543210;
  LUT6 desc2793(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[27:27]),.I3(q_reg_1[27:27]),.I4(q_reg_2[27:27]),.I5(q_reg_3[27:27]),.O(ram_buffer_0_2[27:27]));
defparam desc2793.INIT=64'hFEDCBA9876543210;
  LUT6 desc2794(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[28:28]),.I3(q_reg_1[28:28]),.I4(q_reg_2[28:28]),.I5(q_reg_3[28:28]),.O(ram_buffer_1_1[28:28]));
defparam desc2794.INIT=64'hFEDCBA9876543210;
  LUT6 desc2795(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[28:28]),.I3(q_reg_1[28:28]),.I4(q_reg_2[28:28]),.I5(q_reg_3[28:28]),.O(ram_buffer_0_2[28:28]));
defparam desc2795.INIT=64'hFEDCBA9876543210;
  LUT6 desc2796(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[29:29]),.I3(q_reg_1[29:29]),.I4(q_reg_2[29:29]),.I5(q_reg_3[29:29]),.O(ram_buffer_1_1[29:29]));
defparam desc2796.INIT=64'hFEDCBA9876543210;
  LUT6 desc2797(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[29:29]),.I3(q_reg_1[29:29]),.I4(q_reg_2[29:29]),.I5(q_reg_3[29:29]),.O(ram_buffer_0_2[29:29]));
defparam desc2797.INIT=64'hFEDCBA9876543210;
  LUT6 desc2798(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[30:30]),.I3(q_reg_1[30:30]),.I4(q_reg_2[30:30]),.I5(q_reg_3[30:30]),.O(ram_buffer_1_1[30:30]));
defparam desc2798.INIT=64'hFEDCBA9876543210;
  LUT6 desc2799(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[30:30]),.I3(q_reg_1[30:30]),.I4(q_reg_2[30:30]),.I5(q_reg_3[30:30]),.O(ram_buffer_0_2[30:30]));
defparam desc2799.INIT=64'hFEDCBA9876543210;
  LUT6 desc2800(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[31:31]),.I3(q_reg_1[31:31]),.I4(q_reg_2[31:31]),.I5(q_reg_3[31:31]),.O(ram_buffer_1_1[31:31]));
defparam desc2800.INIT=64'hFEDCBA9876543210;
  LUT6 desc2801(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[31:31]),.I3(q_reg_1[31:31]),.I4(q_reg_2[31:31]),.I5(q_reg_3[31:31]),.O(ram_buffer_0_2[31:31]));
defparam desc2801.INIT=64'hFEDCBA9876543210;
  LUT6 desc2802(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[32:32]),.I3(q_reg_1[32:32]),.I4(q_reg_2[32:32]),.I5(q_reg_3[32:32]),.O(ram_buffer_1_1[32:32]));
defparam desc2802.INIT=64'hFEDCBA9876543210;
  LUT6 desc2803(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[32:32]),.I3(q_reg_1[32:32]),.I4(q_reg_2[32:32]),.I5(q_reg_3[32:32]),.O(ram_buffer_0_2[32:32]));
defparam desc2803.INIT=64'hFEDCBA9876543210;
  LUT6 desc2804(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[33:33]),.I3(q_reg_1[33:33]),.I4(q_reg_2[33:33]),.I5(q_reg_3[33:33]),.O(ram_buffer_1_1[33:33]));
defparam desc2804.INIT=64'hFEDCBA9876543210;
  LUT6 desc2805(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[33:33]),.I3(q_reg_1[33:33]),.I4(q_reg_2[33:33]),.I5(q_reg_3[33:33]),.O(ram_buffer_0_2[33:33]));
defparam desc2805.INIT=64'hFEDCBA9876543210;
  LUT6 desc2806(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[34:34]),.I3(q_reg_1[34:34]),.I4(q_reg_2[34:34]),.I5(q_reg_3[34:34]),.O(ram_buffer_1_1[34:34]));
defparam desc2806.INIT=64'hFEDCBA9876543210;
  LUT6 desc2807(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[34:34]),.I3(q_reg_1[34:34]),.I4(q_reg_2[34:34]),.I5(q_reg_3[34:34]),.O(ram_buffer_0_2[34:34]));
defparam desc2807.INIT=64'hFEDCBA9876543210;
  LUT6 desc2808(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[35:35]),.I3(q_reg_1[35:35]),.I4(q_reg_2[35:35]),.I5(q_reg_3[35:35]),.O(ram_buffer_1_1[35:35]));
defparam desc2808.INIT=64'hFEDCBA9876543210;
  LUT6 desc2809(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[35:35]),.I3(q_reg_1[35:35]),.I4(q_reg_2[35:35]),.I5(q_reg_3[35:35]),.O(ram_buffer_0_2[35:35]));
defparam desc2809.INIT=64'hFEDCBA9876543210;
  LUT6 desc2810(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[36:36]),.I3(q_reg_1[36:36]),.I4(q_reg_2[36:36]),.I5(q_reg_3[36:36]),.O(ram_buffer_1_1[36:36]));
defparam desc2810.INIT=64'hFEDCBA9876543210;
  LUT6 desc2811(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[36:36]),.I3(q_reg_1[36:36]),.I4(q_reg_2[36:36]),.I5(q_reg_3[36:36]),.O(ram_buffer_0_2[36:36]));
defparam desc2811.INIT=64'hFEDCBA9876543210;
  LUT6 desc2812(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[37:37]),.I3(q_reg_1[37:37]),.I4(q_reg_2[37:37]),.I5(q_reg_3[37:37]),.O(ram_buffer_1_1[37:37]));
defparam desc2812.INIT=64'hFEDCBA9876543210;
  LUT6 desc2813(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[37:37]),.I3(q_reg_1[37:37]),.I4(q_reg_2[37:37]),.I5(q_reg_3[37:37]),.O(ram_buffer_0_2[37:37]));
defparam desc2813.INIT=64'hFEDCBA9876543210;
  LUT6 desc2814(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[38:38]),.I3(q_reg_1[38:38]),.I4(q_reg_2[38:38]),.I5(q_reg_3[38:38]),.O(ram_buffer_1_1[38:38]));
defparam desc2814.INIT=64'hFEDCBA9876543210;
  LUT6 desc2815(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[38:38]),.I3(q_reg_1[38:38]),.I4(q_reg_2[38:38]),.I5(q_reg_3[38:38]),.O(ram_buffer_0_2[38:38]));
defparam desc2815.INIT=64'hFEDCBA9876543210;
  LUT6 desc2816(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[39:39]),.I3(q_reg_1[39:39]),.I4(q_reg_2[39:39]),.I5(q_reg_3[39:39]),.O(ram_buffer_1_1[39:39]));
defparam desc2816.INIT=64'hFEDCBA9876543210;
  LUT6 desc2817(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[39:39]),.I3(q_reg_1[39:39]),.I4(q_reg_2[39:39]),.I5(q_reg_3[39:39]),.O(ram_buffer_0_2[39:39]));
defparam desc2817.INIT=64'hFEDCBA9876543210;
  LUT6 desc2818(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[40:40]),.I3(q_reg_1[40:40]),.I4(q_reg_2[40:40]),.I5(q_reg_3[40:40]),.O(ram_buffer_1_1[40:40]));
defparam desc2818.INIT=64'hFEDCBA9876543210;
  LUT6 desc2819(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[40:40]),.I3(q_reg_1[40:40]),.I4(q_reg_2[40:40]),.I5(q_reg_3[40:40]),.O(ram_buffer_0_2[40:40]));
defparam desc2819.INIT=64'hFEDCBA9876543210;
  LUT6 desc2820(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[41:41]),.I3(q_reg_1[41:41]),.I4(q_reg_2[41:41]),.I5(q_reg_3[41:41]),.O(ram_buffer_1_1[41:41]));
defparam desc2820.INIT=64'hFEDCBA9876543210;
  LUT6 desc2821(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[41:41]),.I3(q_reg_1[41:41]),.I4(q_reg_2[41:41]),.I5(q_reg_3[41:41]),.O(ram_buffer_0_2[41:41]));
defparam desc2821.INIT=64'hFEDCBA9876543210;
  LUT6 desc2822(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[42:42]),.I3(q_reg_1[42:42]),.I4(q_reg_2[42:42]),.I5(q_reg_3[42:42]),.O(ram_buffer_1_1[42:42]));
defparam desc2822.INIT=64'hFEDCBA9876543210;
  LUT6 desc2823(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[42:42]),.I3(q_reg_1[42:42]),.I4(q_reg_2[42:42]),.I5(q_reg_3[42:42]),.O(ram_buffer_0_2[42:42]));
defparam desc2823.INIT=64'hFEDCBA9876543210;
  LUT6 desc2824(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[43:43]),.I3(q_reg_1[43:43]),.I4(q_reg_2[43:43]),.I5(q_reg_3[43:43]),.O(ram_buffer_1_1[43:43]));
defparam desc2824.INIT=64'hFEDCBA9876543210;
  LUT6 desc2825(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[43:43]),.I3(q_reg_1[43:43]),.I4(q_reg_2[43:43]),.I5(q_reg_3[43:43]),.O(ram_buffer_0_2[43:43]));
defparam desc2825.INIT=64'hFEDCBA9876543210;
  LUT6 desc2826(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[44:44]),.I3(q_reg_1[44:44]),.I4(q_reg_2[44:44]),.I5(q_reg_3[44:44]),.O(ram_buffer_1_1[44:44]));
defparam desc2826.INIT=64'hFEDCBA9876543210;
  LUT6 desc2827(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[44:44]),.I3(q_reg_1[44:44]),.I4(q_reg_2[44:44]),.I5(q_reg_3[44:44]),.O(ram_buffer_0_2[44:44]));
defparam desc2827.INIT=64'hFEDCBA9876543210;
  LUT6 desc2828(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[45:45]),.I3(q_reg_1[45:45]),.I4(q_reg_2[45:45]),.I5(q_reg_3[45:45]),.O(ram_buffer_1_1[45:45]));
defparam desc2828.INIT=64'hFEDCBA9876543210;
  LUT6 desc2829(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[45:45]),.I3(q_reg_1[45:45]),.I4(q_reg_2[45:45]),.I5(q_reg_3[45:45]),.O(ram_buffer_0_2[45:45]));
defparam desc2829.INIT=64'hFEDCBA9876543210;
  LUT6 desc2830(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[46:46]),.I3(q_reg_1[46:46]),.I4(q_reg_2[46:46]),.I5(q_reg_3[46:46]),.O(ram_buffer_1_1[46:46]));
defparam desc2830.INIT=64'hFEDCBA9876543210;
  LUT6 desc2831(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[46:46]),.I3(q_reg_1[46:46]),.I4(q_reg_2[46:46]),.I5(q_reg_3[46:46]),.O(ram_buffer_0_2[46:46]));
defparam desc2831.INIT=64'hFEDCBA9876543210;
  LUT6 desc2832(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[47:47]),.I3(q_reg_1[47:47]),.I4(q_reg_2[47:47]),.I5(q_reg_3[47:47]),.O(ram_buffer_1_1[47:47]));
defparam desc2832.INIT=64'hFEDCBA9876543210;
  LUT6 desc2833(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[47:47]),.I3(q_reg_1[47:47]),.I4(q_reg_2[47:47]),.I5(q_reg_3[47:47]),.O(ram_buffer_0_2[47:47]));
defparam desc2833.INIT=64'hFEDCBA9876543210;
  LUT6 desc2834(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[48:48]),.I3(q_reg_1[48:48]),.I4(q_reg_2[48:48]),.I5(q_reg_3[48:48]),.O(ram_buffer_1_1[48:48]));
defparam desc2834.INIT=64'hFEDCBA9876543210;
  LUT6 desc2835(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[48:48]),.I3(q_reg_1[48:48]),.I4(q_reg_2[48:48]),.I5(q_reg_3[48:48]),.O(ram_buffer_0_2[48:48]));
defparam desc2835.INIT=64'hFEDCBA9876543210;
  LUT6 desc2836(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[49:49]),.I3(q_reg_1[49:49]),.I4(q_reg_2[49:49]),.I5(q_reg_3[49:49]),.O(ram_buffer_1_1[49:49]));
defparam desc2836.INIT=64'hFEDCBA9876543210;
  LUT6 desc2837(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[49:49]),.I3(q_reg_1[49:49]),.I4(q_reg_2[49:49]),.I5(q_reg_3[49:49]),.O(ram_buffer_0_2[49:49]));
defparam desc2837.INIT=64'hFEDCBA9876543210;
  LUT6 desc2838(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[50:50]),.I3(q_reg_1[50:50]),.I4(q_reg_2[50:50]),.I5(q_reg_3[50:50]),.O(ram_buffer_1_1[50:50]));
defparam desc2838.INIT=64'hFEDCBA9876543210;
  LUT6 desc2839(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[50:50]),.I3(q_reg_1[50:50]),.I4(q_reg_2[50:50]),.I5(q_reg_3[50:50]),.O(ram_buffer_0_2[50:50]));
defparam desc2839.INIT=64'hFEDCBA9876543210;
  LUT6 desc2840(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[51:51]),.I3(q_reg_1[51:51]),.I4(q_reg_2[51:51]),.I5(q_reg_3[51:51]),.O(ram_buffer_1_1[51:51]));
defparam desc2840.INIT=64'hFEDCBA9876543210;
  LUT6 desc2841(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[51:51]),.I3(q_reg_1[51:51]),.I4(q_reg_2[51:51]),.I5(q_reg_3[51:51]),.O(ram_buffer_0_2[51:51]));
defparam desc2841.INIT=64'hFEDCBA9876543210;
  LUT6 desc2842(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[52:52]),.I3(q_reg_1[52:52]),.I4(q_reg_2[52:52]),.I5(q_reg_3[52:52]),.O(ram_buffer_1_1[52:52]));
defparam desc2842.INIT=64'hFEDCBA9876543210;
  LUT6 desc2843(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[52:52]),.I3(q_reg_1[52:52]),.I4(q_reg_2[52:52]),.I5(q_reg_3[52:52]),.O(ram_buffer_0_2[52:52]));
defparam desc2843.INIT=64'hFEDCBA9876543210;
  LUT6 desc2844(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[53:53]),.I3(q_reg_1[53:53]),.I4(q_reg_2[53:53]),.I5(q_reg_3[53:53]),.O(ram_buffer_1_1[53:53]));
defparam desc2844.INIT=64'hFEDCBA9876543210;
  LUT6 desc2845(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[53:53]),.I3(q_reg_1[53:53]),.I4(q_reg_2[53:53]),.I5(q_reg_3[53:53]),.O(ram_buffer_0_2[53:53]));
defparam desc2845.INIT=64'hFEDCBA9876543210;
  LUT6 desc2846(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[54:54]),.I3(q_reg_1[54:54]),.I4(q_reg_2[54:54]),.I5(q_reg_3[54:54]),.O(ram_buffer_1_1[54:54]));
defparam desc2846.INIT=64'hFEDCBA9876543210;
  LUT6 desc2847(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[54:54]),.I3(q_reg_1[54:54]),.I4(q_reg_2[54:54]),.I5(q_reg_3[54:54]),.O(ram_buffer_0_2[54:54]));
defparam desc2847.INIT=64'hFEDCBA9876543210;
  LUT6 desc2848(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[55:55]),.I3(q_reg_1[55:55]),.I4(q_reg_2[55:55]),.I5(q_reg_3[55:55]),.O(ram_buffer_1_1[55:55]));
defparam desc2848.INIT=64'hFEDCBA9876543210;
  LUT6 desc2849(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[55:55]),.I3(q_reg_1[55:55]),.I4(q_reg_2[55:55]),.I5(q_reg_3[55:55]),.O(ram_buffer_0_2[55:55]));
defparam desc2849.INIT=64'hFEDCBA9876543210;
  LUT6 desc2850(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[56:56]),.I3(q_reg_1[56:56]),.I4(q_reg_2[56:56]),.I5(q_reg_3[56:56]),.O(ram_buffer_1_1[56:56]));
defparam desc2850.INIT=64'hFEDCBA9876543210;
  LUT6 desc2851(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[56:56]),.I3(q_reg_1[56:56]),.I4(q_reg_2[56:56]),.I5(q_reg_3[56:56]),.O(ram_buffer_0_2[56:56]));
defparam desc2851.INIT=64'hFEDCBA9876543210;
  LUT6 desc2852(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[57:57]),.I3(q_reg_1[57:57]),.I4(q_reg_2[57:57]),.I5(q_reg_3[57:57]),.O(ram_buffer_1_1[57:57]));
defparam desc2852.INIT=64'hFEDCBA9876543210;
  LUT6 desc2853(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[57:57]),.I3(q_reg_1[57:57]),.I4(q_reg_2[57:57]),.I5(q_reg_3[57:57]),.O(ram_buffer_0_2[57:57]));
defparam desc2853.INIT=64'hFEDCBA9876543210;
  LUT6 desc2854(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[58:58]),.I3(q_reg_1[58:58]),.I4(q_reg_2[58:58]),.I5(q_reg_3[58:58]),.O(ram_buffer_1_1[58:58]));
defparam desc2854.INIT=64'hFEDCBA9876543210;
  LUT6 desc2855(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[58:58]),.I3(q_reg_1[58:58]),.I4(q_reg_2[58:58]),.I5(q_reg_3[58:58]),.O(ram_buffer_0_2[58:58]));
defparam desc2855.INIT=64'hFEDCBA9876543210;
  LUT6 desc2856(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[59:59]),.I3(q_reg_1[59:59]),.I4(q_reg_2[59:59]),.I5(q_reg_3[59:59]),.O(ram_buffer_1_1[59:59]));
defparam desc2856.INIT=64'hFEDCBA9876543210;
  LUT6 desc2857(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[59:59]),.I3(q_reg_1[59:59]),.I4(q_reg_2[59:59]),.I5(q_reg_3[59:59]),.O(ram_buffer_0_2[59:59]));
defparam desc2857.INIT=64'hFEDCBA9876543210;
  LUT6 desc2858(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[60:60]),.I3(q_reg_1[60:60]),.I4(q_reg_2[60:60]),.I5(q_reg_3[60:60]),.O(ram_buffer_1_1[60:60]));
defparam desc2858.INIT=64'hFEDCBA9876543210;
  LUT6 desc2859(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[60:60]),.I3(q_reg_1[60:60]),.I4(q_reg_2[60:60]),.I5(q_reg_3[60:60]),.O(ram_buffer_0_2[60:60]));
defparam desc2859.INIT=64'hFEDCBA9876543210;
  LUT6 desc2860(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[61:61]),.I3(q_reg_1[61:61]),.I4(q_reg_2[61:61]),.I5(q_reg_3[61:61]),.O(ram_buffer_1_1[61:61]));
defparam desc2860.INIT=64'hFEDCBA9876543210;
  LUT6 desc2861(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[61:61]),.I3(q_reg_1[61:61]),.I4(q_reg_2[61:61]),.I5(q_reg_3[61:61]),.O(ram_buffer_0_2[61:61]));
defparam desc2861.INIT=64'hFEDCBA9876543210;
  LUT6 desc2862(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[62:62]),.I3(q_reg_1[62:62]),.I4(q_reg_2[62:62]),.I5(q_reg_3[62:62]),.O(ram_buffer_1_1[62:62]));
defparam desc2862.INIT=64'hFEDCBA9876543210;
  LUT6 desc2863(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[62:62]),.I3(q_reg_1[62:62]),.I4(q_reg_2[62:62]),.I5(q_reg_3[62:62]),.O(ram_buffer_0_2[62:62]));
defparam desc2863.INIT=64'hFEDCBA9876543210;
  LUT6 desc2864(.I0(read_ram_ptr_d_1[0:0]),.I1(read_ram_ptr_d_1[1:1]),.I2(q_reg_0[63:63]),.I3(q_reg_1[63:63]),.I4(q_reg_2[63:63]),.I5(q_reg_3[63:63]),.O(ram_buffer_1_1[63:63]));
defparam desc2864.INIT=64'hFEDCBA9876543210;
  LUT6 desc2865(.I0(read_ram_ptr_d_0[0:0]),.I1(read_ram_ptr_d_0[1:1]),.I2(q_reg_0[63:63]),.I3(q_reg_1[63:63]),.I4(q_reg_2[63:63]),.I5(q_reg_3[63:63]),.O(ram_buffer_0_2[63:63]));
defparam desc2865.INIT=64'hFEDCBA9876543210;
  LUT3 desc2866(.I0(write_window_complete),.I1(write_last_window_complete),.I2(next_traceback),.O(N_41_mux));
defparam desc2866.INIT=8'h0E;
  LUT6 read_addr_ptr_1_1_sqmuxa_3_cZ(.I0(reorder_tvalid_fast[1:1]),.I1(ram_tvalid[1:1]),.I2(read_ram_fsm_1_0_rep1),.I3(traceback_tvalid[1:1]),.I4(read_ram_fsm_1[1:1]),.I5(un64_m_axis_output_tready),.O(read_addr_ptr_1_1_sqmuxa_3));
defparam read_addr_ptr_1_1_sqmuxa_3_cZ.INIT=64'h2000000070F00000;
  LUT5_L desc2867(.I0(aresetn),.I1(ram_tvalid[1:1]),.I2(traceback_tvalid[1:1]),.I3(reorder_tvalid_1_rep1),.I4(ram_buffer_full[1:1]),.LO(ram_buffer_full_nss[1:1]));
defparam desc2867.INIT=32'hA2228000;
  LUT6 read_ram_fsm_0_2_sqmuxa_0_cZ(.I0(read_ram_fsm_0_0_rep1),.I1(read_addr_ptr_0[0:0]),.I2(read_addr_ptr_0[1:1]),.I3(read_addr_ptr_0[2:2]),.I4(read_ram_fsm_0_1_rep1),.I5(un6_m_axis_output_tready_3),.O(read_ram_fsm_0_2_sqmuxa_0));
defparam read_ram_fsm_0_2_sqmuxa_0_cZ.INIT=64'h0000AAA80000AAAA;
  LUT6 desc2868(.I0(read_ram_ptr_1[1:1]),.I1(read_ram_ptr_1[0:0]),.I2(read_ram_fsm_0_0_rep1),.I3(read_ram_fsm_0_1_rep1),.I4(read_ram_ptr_0[1:1]),.I5(read_ram_ptr_0[0:0]),.O(un44_m_axis_output_tready));
defparam desc2868.INIT=64'h0010002000800040;
  LUT6 desc2869(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_1[2:2]),.I2(read_addr_ptr_1[0:0]),.I3(un21_m_axis_output_tready_axb_0),.I4(un21_m_axis_output_tready_s_1),.I5(un21_m_axis_output_tready_s_2),.O(un57_m_axis_output_tready_0_N_11));
defparam desc2869.INIT=64'h8008400420021001;
  LUT6 desc2870(.I0(read_addr_ptr_0[0:0]),.I1(read_addr_ptr_0[1:1]),.I2(read_addr_ptr_0[2:2]),.I3(un21_m_axis_output_tready_axb_0),.I4(un21_m_axis_output_tready_s_1),.I5(un21_m_axis_output_tready_s_2),.O(un23_m_axis_output_tready_0_N_11));
defparam desc2870.INIT=64'h8040201008040201;
  LUT5 desc2871(.I0(read_addr_ptr_0[1:1]),.I1(read_addr_ptr_0[2:2]),.I2(un30_m_axis_output_tready_0_N_14),.I3(un18_m_axis_output_tready[1:1]),.I4(un18_m_axis_output_tready[2:2]),.O(un30_m_axis_output_tready_0_N_11));
defparam desc2871.INIT=32'h08040201;
  LUT6 desc2872(.I0(window_length[1:1]),.I1(window_length[2:2]),.I2(window_length[0:0]),.I3(write_addr_ptr[1:1]),.I4(write_addr_ptr[2:2]),.I5(write_addr_ptr[0:0]),.O(un9_s_axis_input_tvalid_0_N_11));
defparam desc2872.INIT=64'h0108040280402010;
  LUT6_L desc2873(.I0(ram_window_tuser[0:0]),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(un13_write_last_window_complete),.I4(N_99),.I5(un23_m_axis_output_tready),.LO(m_axis_output_window_tuser_int_RNO[0:0]));
defparam desc2873.INIT=64'hABA8BBB8ABA8ABA8;
  LUT6 desc2874(.I0(s_axis_ctrl_tvalid),.I1(write_ram_fsm_fast[4:4]),.I2(read_ram_fsm_0_0_rep1),.I3(read_ram_fsm_0_1_rep1),.I4(read_ram_fsm_1_1_rep1),.I5(read_ram_fsm_1_0_rep1),.O(N_1754));
defparam desc2874.INIT=64'h0000000000000008;
  LUT5 read_ram_fsm_1_1_sqmuxa_2_0_a2(.I0(reorder_tvalid_fast[1:1]),.I1(read_ram_fsm_1_1_rep1),.I2(read_ram_fsm_1_0_rep1),.I3(traceback_tvalid[1:1]),.I4(N_743),.O(N_745));
defparam read_ram_fsm_1_1_sqmuxa_2_0_a2.INIT=32'h10300000;
  LUT6 read_ram_fsm_0_0_sqmuxa_cZ(.I0(reorder_tvalid_fast[0:0]),.I1(read_addr_ptr_0[0:0]),.I2(read_addr_ptr_0[1:1]),.I3(read_addr_ptr_0[2:2]),.I4(traceback_tvalid[0:0]),.I5(un6_m_axis_output_tready_3),.O(read_ram_fsm_0_0_sqmuxa));
defparam read_ram_fsm_0_0_sqmuxa_cZ.INIT=64'h0001000300000000;
  LUT6 un1_read_addr_ptr_1_1_sqmuxa_0_cZ(.I0(write_window_complete),.I1(write_last_window_complete),.I2(next_traceback),.I3(N_720),.I4(N_1733),.I5(N_743),.O(un1_read_addr_ptr_1_1_sqmuxa_0));
defparam un1_read_addr_ptr_1_1_sqmuxa_0_cZ.INIT=64'h0000202000FF20FF;
  LUT6_L desc2875(.I0(read_addr_ptr_0[6:6]),.I1(read_addr_ptr_0[1:1]),.I2(un30_m_axis_output_tready_0_N_14),.I3(N_99),.I4(un18_m_axis_output_tready[1:1]),.I5(un18_m_axis_output_tready[6:6]),.LO(m33_2));
defparam desc2875.INIT=64'h0008000200040001;
  LUT5 desc2876(.I0(window_length[3:3]),.I1(write_addr_ptr[3:3]),.I2(write_addr_ptr[1:1]),.I3(write_addr_ptr[2:2]),.I4(write_addr_ptr[0:0]),.O(N_2339));
defparam desc2876.INIT=32'h69999999;
  LUT4 un27_s_axis_input_tready_int_c(.I0(write_ram_fsm_fast[0:0]),.I1(write_ram_fsm_fast[4:4]),.I2(write_ram_fsm_1),.I3(N_1756_1),.O(un27_s_axis_input_tready_int));
defparam un27_s_axis_input_tready_int_c.INIT=16'hFEFF;
  LUT6 desc2877(.I0(read_addr_ptr_1[3:3]),.I1(read_addr_ptr_1[4:4]),.I2(un18_m_axis_output_tready[3:3]),.I3(un18_m_axis_output_tready[4:4]),.I4(m33_0_2),.I5(m33_0),.O(N_54_mux_0));
defparam desc2877.INIT=64'h8421000000000000;
  LUT6_L desc2878(.I0(traceback_tvalid[1:1]),.I1(reorder_tvalid_1_rep1),.I2(read_ram_fsm_1[0:0]),.I3(read_ram_fsm_1[1:1]),.I4(un1_m_axis_output_window_tuser_int_0_sqmuxa_set_0),.I5(un57_m_axis_output_tready),.LO(m_axis_output_window_tuser_int_RNO[1:1]));
defparam desc2878.INIT=64'hFFFF0070FFFF0000;
  LUT4_L desc2879(.I0(write_window_complete),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(next_traceback),.LO(m_axis_output_tvalid_int_RNO));
defparam desc2879.INIT=16'hF0F2;
  LUT6 wen_ram_0_sqmuxa_3_cZ(.I0(aresetn),.I1(s_axis_ctrl_tvalid),.I2(read_ram_fsm_1_1_rep1),.I3(read_ram_fsm_1_0_rep1),.I4(write_ram_fsm_4_rep1),.I5(read_ram_fsm_0_d_i_0[3:3]),.O(wen_ram_0_sqmuxa_3));
defparam wen_ram_0_sqmuxa_3_cZ.INIT=64'h0000000000080000;
  LUT6_L desc2880(.I0(ram_last_tuser[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep1),.I3(read_ram_fsm_1[0:0]),.I4(read_ram_fsm_1[1:1]),.I5(un64_m_axis_output_tready),.LO(m_axis_output_last_tuser_int[1:1]));
defparam desc2880.INIT=64'hBFAA0000AAAA0000;
  LUT6 desc2881(.I0(read_addr_ptr_0[4:4]),.I1(read_addr_ptr_0[5:5]),.I2(un18_m_axis_output_tready[4:4]),.I3(un18_m_axis_output_tready[5:5]),.I4(m33_1),.I5(m33_2),.O(N_54_mux));
defparam desc2881.INIT=64'h8421000000000000;
  LUT4 desc2882(.I0(write_addr_ptr[3:3]),.I1(write_addr_ptr[1:1]),.I2(write_addr_ptr[2:2]),.I3(write_addr_ptr[0:0]),.O(un9_s_axis_input_tvalid_a_4_c4));
defparam desc2882.INIT=16'h7FFF;
  LUT5 desc2883(.I0(write_addr_ptr[6:6]),.I1(read_addr_ptr_0[6:6]),.I2(read_addr_ptr_1[6:6]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[6:6]));
defparam desc2883.INIT=32'hAACCAAF0;
  LUT5 desc2884(.I0(read_addr_ptr_0[5:5]),.I1(read_addr_ptr_1[5:5]),.I2(write_addr_ptr[5:5]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[5:5]));
defparam desc2884.INIT=32'hF0AAF0CC;
  LUT5 desc2885(.I0(read_addr_ptr_0[4:4]),.I1(read_addr_ptr_1[4:4]),.I2(write_addr_ptr[4:4]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[4:4]));
defparam desc2885.INIT=32'hF0AAF0CC;
  LUT5 desc2886(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_1[3:3]),.I2(write_addr_ptr[3:3]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[3:3]));
defparam desc2886.INIT=32'hF0AAF0CC;
  LUT5 desc2887(.I0(read_addr_ptr_1[2:2]),.I1(read_addr_ptr_0[2:2]),.I2(write_addr_ptr[2:2]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[2:2]));
defparam desc2887.INIT=32'hF0CCF0AA;
  LUT5 desc2888(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_0[1:1]),.I2(write_addr_ptr[1:1]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[1:1]));
defparam desc2888.INIT=32'hF0CCF0AA;
  LUT5 desc2889(.I0(read_addr_ptr_0[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(write_addr_ptr[0:0]),.I3(un42_addr),.I4(un55_addr),.O(addr_1[0:0]));
defparam desc2889.INIT=32'hF0AAF0CC;
  LUT5 desc2890(.I0(read_addr_ptr_0[5:5]),.I1(read_addr_ptr_1[5:5]),.I2(write_addr_ptr[5:5]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[5:5]));
defparam desc2890.INIT=32'hF0AAF0CC;
  LUT5 desc2891(.I0(read_addr_ptr_1[2:2]),.I1(read_addr_ptr_0[2:2]),.I2(write_addr_ptr[2:2]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[2:2]));
defparam desc2891.INIT=32'hF0CCF0AA;
  LUT5 desc2892(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_0[1:1]),.I2(write_addr_ptr[1:1]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[1:1]));
defparam desc2892.INIT=32'hF0CCF0AA;
  LUT5 desc2893(.I0(read_addr_ptr_0[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(write_addr_ptr[0:0]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[0:0]));
defparam desc2893.INIT=32'hF0AAF0CC;
  LUT5 desc2894(.I0(read_addr_ptr_0[5:5]),.I1(read_addr_ptr_1[5:5]),.I2(write_addr_ptr[5:5]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[5:5]));
defparam desc2894.INIT=32'hF0AAF0CC;
  LUT5 desc2895(.I0(read_addr_ptr_1[2:2]),.I1(read_addr_ptr_0[2:2]),.I2(write_addr_ptr[2:2]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[2:2]));
defparam desc2895.INIT=32'hF0CCF0AA;
  LUT5 desc2896(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_0[1:1]),.I2(write_addr_ptr[1:1]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[1:1]));
defparam desc2896.INIT=32'hF0CCF0AA;
  LUT5 desc2897(.I0(read_addr_ptr_0[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(write_addr_ptr[0:0]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[0:0]));
defparam desc2897.INIT=32'hF0AAF0CC;
  LUT5 desc2898(.I0(read_addr_ptr_0[4:4]),.I1(read_addr_ptr_1[4:4]),.I2(write_addr_ptr[4:4]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[4:4]));
defparam desc2898.INIT=32'hF0AAF0CC;
  LUT5 desc2899(.I0(read_addr_ptr_0[4:4]),.I1(read_addr_ptr_1[4:4]),.I2(write_addr_ptr[4:4]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[4:4]));
defparam desc2899.INIT=32'hF0AAF0CC;
  LUT5 desc2900(.I0(write_addr_ptr[6:6]),.I1(read_addr_ptr_0[6:6]),.I2(read_addr_ptr_1[6:6]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[6:6]));
defparam desc2900.INIT=32'hAACCAAF0;
  LUT5 desc2901(.I0(read_addr_ptr_0[5:5]),.I1(read_addr_ptr_1[5:5]),.I2(write_addr_ptr[5:5]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[5:5]));
defparam desc2901.INIT=32'hF0AAF0CC;
  LUT5 desc2902(.I0(read_addr_ptr_0[4:4]),.I1(read_addr_ptr_1[4:4]),.I2(write_addr_ptr[4:4]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[4:4]));
defparam desc2902.INIT=32'hF0AAF0CC;
  LUT5 desc2903(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_1[3:3]),.I2(write_addr_ptr[3:3]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[3:3]));
defparam desc2903.INIT=32'hF0AAF0CC;
  LUT5 desc2904(.I0(read_addr_ptr_1[2:2]),.I1(read_addr_ptr_0[2:2]),.I2(write_addr_ptr[2:2]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[2:2]));
defparam desc2904.INIT=32'hF0CCF0AA;
  LUT5 desc2905(.I0(read_addr_ptr_1[1:1]),.I1(read_addr_ptr_0[1:1]),.I2(write_addr_ptr[1:1]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[1:1]));
defparam desc2905.INIT=32'hF0CCF0AA;
  LUT5 desc2906(.I0(read_addr_ptr_0[0:0]),.I1(read_addr_ptr_1[0:0]),.I2(write_addr_ptr[0:0]),.I3(un74_addr),.I4(un87_addr),.O(addr_2[0:0]));
defparam desc2906.INIT=32'hF0AAF0CC;
  LUT5 desc2907(.I0(write_addr_ptr[6:6]),.I1(read_addr_ptr_0[6:6]),.I2(read_addr_ptr_1[6:6]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[6:6]));
defparam desc2907.INIT=32'hAACCAAF0;
  LUT5 desc2908(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_1[3:3]),.I2(write_addr_ptr[3:3]),.I3(un3_addr),.I4(un16_addr),.O(addr_0[3:3]));
defparam desc2908.INIT=32'hF0AAF0CC;
  LUT5 desc2909(.I0(write_addr_ptr[6:6]),.I1(read_addr_ptr_0[6:6]),.I2(read_addr_ptr_1[6:6]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[6:6]));
defparam desc2909.INIT=32'hAACCAAF0;
  LUT5 desc2910(.I0(read_addr_ptr_0[3:3]),.I1(read_addr_ptr_1[3:3]),.I2(write_addr_ptr[3:3]),.I3(un106_addr),.I4(un119_addr),.O(addr_3[3:3]));
defparam desc2910.INIT=32'hF0AAF0CC;
  LUT5 un1_read_ram_ptr_0_1_sqmuxa_1_cZ(.I0(read_ram_fsm_0_0_rep1),.I1(read_ram_fsm_0_1_rep1),.I2(N_41_mux),.I3(un10_m_axis_output_tready),.I4(read_ram_fsm_0_0_sqmuxa),.O(un1_read_ram_ptr_0_1_sqmuxa_1));
defparam un1_read_ram_ptr_0_1_sqmuxa_1_cZ.INIT=32'h01670145;
  LUT5 desc2911(.I0(aresetn),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(un10_m_axis_output_tready),.I4(read_ram_fsm_0_0_sqmuxa),.O(un1_read_addr_ptr_0_1_sqmuxa_2_f0_0[6:6]));
defparam desc2911.INIT=32'h8AAAAAAA;
  LUT6 un1_read_addr_ptr_1_1_sqmuxa_1_1_cZ(.I0(reorder_tvalid_fast[1:1]),.I1(ram_tvalid[1:1]),.I2(read_ram_fsm_1_1_rep1),.I3(read_ram_fsm_1_0_rep1),.I4(traceback_tvalid[1:1]),.I5(un44_m_axis_output_tready),.O(un1_read_addr_ptr_1_1_sqmuxa_1_1));
defparam un1_read_addr_ptr_1_1_sqmuxa_1_1_cZ.INIT=64'h8AF000F08A000000;
  LUT5 desc2912(.I0(write_ram_fsm[2:2]),.I1(acs_tvalid),.I2(write_ram_fsm_1),.I3(N_1731),.I4(N_1756_1),.O(write_ram_fsm_ns_0_0[2:2]));
defparam desc2912.INIT=32'hF222FAAA;
  LUT5 desc2913(.I0(write_window_complete),.I1(acs_tvalid),.I2(write_ram_fsm_0),.I3(N_1731),.I4(N_1756_1),.O(write_ram_fsm_ns_i_0[4:4]));
defparam desc2913.INIT=32'h57035F0F;
  LUT4 write_ram_ptr_0_sqmuxa_1_cZ(.I0(acs_tlast),.I1(write_ram_fsm[2:2]),.I2(acs_tvalid),.I3(un27_s_axis_input_tready_int),.O(write_ram_ptr_0_sqmuxa_1));
defparam write_ram_ptr_0_sqmuxa_1_cZ.INIT=16'h0080;
  LUT5 desc2914(.I0(aresetn),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(un44_m_axis_output_tready),.I4(N_745),.O(un2_write_ram_ptr_2_1[1:1]));
defparam desc2914.INIT=32'h00AA0020;
  LUT5 desc2915(.I0(aresetn),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(un10_m_axis_output_tready),.I4(read_ram_fsm_0_0_sqmuxa),.O(un2_write_ram_ptr_3_1[1:1]));
defparam desc2915.INIT=32'h00280008;
  LUT5_L desc2916(.I0(ram_tlast[1:1]),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(m_axis_output_tlast_int_0_sqmuxa_1_1),.I4(un64_m_axis_output_tready),.LO(m_axis_output_tlast_int[1:1]));
defparam desc2916.INIT=32'hE0A0A0A0;
  LUT6_L desc2917(.I0(ram_tlast[0:0]),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(m_axis_output_tlast_int_0_sqmuxa_0),.I4(N_99),.I5(un30_m_axis_output_tready),.LO(m_axis_output_tlast_int[0:0]));
defparam desc2917.INIT=64'h8888C88888888888;
  LUT6 un1_write_addr_ptr_0_s_6_RNO(.I0(aresetn),.I1(s_axis_ctrl_tdata_6),.I2(s_axis_ctrl_tdata_22),.I3(write_addr_ptr[6:6]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_0_axb_6));
defparam un1_write_addr_ptr_0_s_6_RNO.INIT=64'hFF00FF00D782FF00;
  LUT6 un1_write_addr_ptr_s_6_RNO(.I0(aresetn),.I1(s_axis_ctrl_tdata_6),.I2(s_axis_ctrl_tdata_22),.I3(write_addr_ptr[6:6]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_6));
defparam un1_write_addr_ptr_s_6_RNO.INIT=64'hFF00FF00D782FF00;
  LUT6 desc2918(.I0(aresetn),.I1(s_axis_ctrl_tdata_5),.I2(s_axis_ctrl_tdata_21),.I3(write_addr_ptr[5:5]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_5));
defparam desc2918.INIT=64'hFF00FF00D782FF00;
  LUT6 desc2919(.I0(aresetn),.I1(s_axis_ctrl_tdata_4),.I2(s_axis_ctrl_tdata_20),.I3(write_addr_ptr[4:4]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_4));
defparam desc2919.INIT=64'hFF00FF00D782FF00;
  LUT6 desc2920(.I0(aresetn),.I1(s_axis_ctrl_tdata_3),.I2(s_axis_ctrl_tdata_19),.I3(write_addr_ptr[3:3]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_3));
defparam desc2920.INIT=64'hFF00FF00D782FF00;
  LUT6 desc2921(.I0(aresetn),.I1(s_axis_ctrl_tdata_2),.I2(s_axis_ctrl_tdata_18),.I3(write_addr_ptr[2:2]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_2));
defparam desc2921.INIT=64'hFF00FF00D782FF00;
  LUT6 desc2922(.I0(aresetn),.I1(s_axis_ctrl_tdata_1),.I2(s_axis_ctrl_tdata_17),.I3(write_addr_ptr[1:1]),.I4(write_ram_fsm_4_rep1),.I5(N_1743),.O(un1_write_addr_ptr_axb_1));
defparam desc2922.INIT=64'hFF00FF00D782FF00;
  LUT6_L write_window_complete_e(.I0(write_ram_fsm[3:3]),.I1(write_window_complete),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1_sqmuxa),.I4(un9_s_axis_input_tvalid),.I5(un1_s_axis_input_tvalid),.LO(write_window_complete_0));
defparam write_window_complete_e.INIT=64'hCCCDCCC8CCC8CCC8;
  LUT6_L write_last_window_complete_e(.I0(write_ram_fsm[3:3]),.I1(write_last_window_complete),.I2(write_ram_fsm_0),.I3(write_ram_fsm_1),.I4(N_1731),.I5(write_ram_ptr_0_sqmuxa_1),.LO(write_last_window_complete_0));
defparam write_last_window_complete_e.INIT=64'hCCDDCCCDCC88CCC8;
  LUT6 read_addr_ptr_0_2_sqmuxa_1_cZ(.I0(aresetn),.I1(read_ram_fsm_0_0_rep1),.I2(read_ram_fsm_0[1:1]),.I3(N_99),.I4(un1_read_ram_ptr_0_1_sqmuxa_1),.I5(un30_m_axis_output_tready),.O(read_addr_ptr_0_2_sqmuxa_1));
defparam read_addr_ptr_0_2_sqmuxa_1_cZ.INIT=64'hAAAA0080AAAA0000;
  LUT6 desc2923(.I0(aresetn),.I1(read_ram_ptr_0[1:1]),.I2(write_ram_ptr[1:1]),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(N_41_mux),.I5(un2_write_ram_ptr_3_1[1:1]),.O(SUM1_3_0));
defparam desc2923.INIT=64'h7755775F880A88A0;
  LUT6 desc2924(.I0(aresetn),.I1(read_ram_ptr_1[1:1]),.I2(write_ram_ptr[1:1]),.I3(N_1733),.I4(N_709),.I5(un2_write_ram_ptr_2_1[1:1]),.O(SUM1_4_0));
defparam desc2924.INIT=64'h775F775588A0880A;
  LUT6_L desc2925(.I0(aresetn),.I1(write_ram_fsm[3:3]),.I2(acs_tvalid),.I3(N_1754),.I4(N_1756_1),.I5(un9_s_axis_input_tvalid),.LO(write_ram_fsm_nss[1:1]));
defparam desc2925.INIT=64'hAA08AA88AA88AA88;
  LUT4 un1_ram_buffer_05_4_cZ(.I0(aresetn),.I1(un1_read_addr_ptr_1_1_sqmuxa_1_1),.I2(un1_read_addr_ptr_1_1_sqmuxa_0),.I3(read_addr_ptr_1_1_sqmuxa_3),.O(un1_ram_buffer_05_4));
defparam un1_ram_buffer_05_4_cZ.INIT=16'hAAA8;
  LUT6_L desc2926(.I0(aresetn),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(un44_m_axis_output_tready),.I4(N_13),.I5(N_54_mux_0),.LO(read_ram_fsm_1_nss[0:0]));
defparam desc2926.INIT=64'h00200A2A80A08AAA;
  LUT5 read_addr_ptr_1_2_sqmuxa_1_cZ(.I0(aresetn),.I1(un44_m_axis_output_tready),.I2(un1_read_ram_ptr_1_1_sqmuxa_0),.I3(N_745),.I4(read_ram_fsm_1_0_sqmuxa_1),.O(read_addr_ptr_1_2_sqmuxa_1));
defparam read_addr_ptr_1_2_sqmuxa_1_cZ.INIT=32'hAAAAA2A0;
  LUT5_L desc2927(.I0(aresetn),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(N_745),.I4(N_54_mux_0),.LO(read_ram_fsm_1_nss[1:1]));
defparam desc2927.INIT=32'h2820A8A0;
  LUT6 desc2928(.I0(aresetn),.I1(read_ram_ptr_0[0:0]),.I2(write_ram_ptr[0:0]),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(N_41_mux),.I5(un2_write_ram_ptr_3_1[1:1]),.O(CO0_3));
defparam desc2928.INIT=64'h88AA88A000A00000;
  LUT6 desc2929(.I0(aresetn),.I1(read_ram_ptr_1[0:0]),.I2(write_ram_ptr[0:0]),.I3(N_1733),.I4(N_709),.I5(un2_write_ram_ptr_2_1[1:1]),.O(CO0_4));
defparam desc2929.INIT=64'h88A088AA000000A0;
  LUT6_L desc2930(.I0(aresetn),.I1(read_ram_ptr_0[0:0]),.I2(write_ram_ptr[0:0]),.I3(read_ram_fsm_0_d_i_0[3:3]),.I4(N_41_mux),.I5(un2_write_ram_ptr_3_1[1:1]),.LO(read_ram_ptr_0_RNO));
defparam desc2930.INIT=64'h7755775F880A88A0;
  LUT6_L desc2931(.I0(aresetn),.I1(read_ram_ptr_1[0:0]),.I2(write_ram_ptr[0:0]),.I3(N_1733),.I4(N_709),.I5(un2_write_ram_ptr_2_1[1:1]),.LO(read_ram_ptr_1_RNO));
defparam desc2931.INIT=64'h775F775588A0880A;
  LUT5_L desc2932(.I0(wen_ram[0:0]),.I1(write_ram_ptr[1:1]),.I2(write_ram_ptr[0:0]),.I3(un9_s_axis_input_tvalid),.I4(un1_write_ram_ptr_0_sqmuxa),.LO(N_1872));
defparam desc2932.INIT=32'hE8ABABAB;
  LUT5_L desc2933(.I0(wen_ram[1:1]),.I1(write_ram_ptr[1:1]),.I2(write_ram_ptr[0:0]),.I3(un9_s_axis_input_tvalid),.I4(un1_write_ram_ptr_0_sqmuxa),.LO(N_1873));
defparam desc2933.INIT=32'h8BBABABA;
  LUT5_L desc2934(.I0(wen_ram[2:2]),.I1(write_ram_ptr[1:1]),.I2(write_ram_ptr[0:0]),.I3(un9_s_axis_input_tvalid),.I4(un1_write_ram_ptr_0_sqmuxa),.LO(N_1874));
defparam desc2934.INIT=32'hB2AEAEAE;
  LUT5_L desc2935(.I0(wen_ram[3:3]),.I1(write_ram_ptr[1:1]),.I2(write_ram_ptr[0:0]),.I3(un9_s_axis_input_tvalid),.I4(un1_write_ram_ptr_0_sqmuxa),.LO(N_1875));
defparam desc2935.INIT=32'h2EEAEAEA;
  LUT6 desc2936(.I0(window_length[4:4]),.I1(window_length[5:5]),.I2(write_addr_ptr[4:4]),.I3(write_addr_ptr[5:5]),.I4(N_2339),.I5(un9_s_axis_input_tvalid_a_4_c4),.O(un9_s_axis_input_tvalid_0_N_4));
defparam desc2936.INIT=64'h8421000018420000;
  LUT4 desc2937(.I0(aresetn),.I1(un9_s_axis_input_tvalid),.I2(un1_s_axis_input_tvalid),.I3(un1_write_ram_ptr_0_sqmuxa),.O(un9_s_axis_input_tvalid_0_I_19_RNIUQCT));
defparam desc2937.INIT=16'hD5F5;
  LUT3 desc2938(.I0(un1_read_addr_ptr_1_1_sqmuxa_0),.I1(read_addr_ptr_1_2_sqmuxa_1),.I2(read_addr_ptr_1_1_sqmuxa_3),.O(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]));
defparam desc2938.INIT=8'hFE;
  LUT6_L desc2939(.I0(aresetn),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(un10_m_axis_output_tready),.I4(N_13_0),.I5(N_54_mux),.LO(read_ram_fsm_0_nss[0:0]));
defparam desc2939.INIT=64'h0008222A8088A2AA;
  LUT6 read_ram_fsm_1_0_sqmuxa_1_RNIIUMB1(.I0(aresetn),.I1(window_length[5:5]),.I2(un44_m_axis_output_tready),.I3(un1_read_ram_ptr_1_1_sqmuxa_0),.I4(N_745),.I5(read_ram_fsm_1_0_sqmuxa_1),.O(window_length_m_0[5:5]));
defparam read_ram_fsm_1_0_sqmuxa_1_RNIIUMB1.INIT=64'h8888888888088800;
  LUT5 un1_read_addr_ptr_1_1_sqmuxa_1_1_RNIOBCO(.I0(aresetn),.I1(read_addr_ptr_1[5:5]),.I2(un1_read_addr_ptr_1_1_sqmuxa_1_1),.I3(un1_read_addr_ptr_1_1_sqmuxa_0),.I4(read_addr_ptr_1_1_sqmuxa_3),.O(read_addr_ptr_1_m[5:5]));
defparam un1_read_addr_ptr_1_1_sqmuxa_1_1_RNIOBCO.INIT=32'h88888880;
  LUT6_L desc2940(.I0(aresetn),.I1(N_1739),.I2(write_ram_fsm_ns_0_a4_0_0[2:2]),.I3(write_ram_fsm_ns_0_0[2:2]),.I4(N_1747),.I5(N_1740),.LO(write_ram_fsm_nss[2:2]));
defparam desc2940.INIT=64'hAA22AA00AAA2AAA0;
  LUT5_L desc2941(.I0(aresetn),.I1(read_ram_fsm_0[1:1]),.I2(read_ram_fsm_0[0:0]),.I3(read_ram_fsm_0_0_sqmuxa),.I4(N_54_mux),.LO(read_ram_fsm_0_nss[1:1]));
defparam desc2941.INIT=32'h2808A888;
  LUT6_L desc2942(.I0(aresetn),.I1(N_1754),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(un1_write_addr_ptr_11[6:6]),.I4(un1_write_addr_ptr_10[6:6]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1791));
defparam desc2942.INIT=64'hFFFF0000FFFD0200;
  LUT6_L desc2943(.I0(aresetn),.I1(N_1754),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(un1_write_addr_ptr_11[5:5]),.I4(un1_write_addr_ptr_10[5:5]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1790));
defparam desc2943.INIT=64'hFFFF0000FFFD0200;
  LUT6_L desc2944(.I0(aresetn),.I1(N_1754),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(un1_write_addr_ptr_11[4:4]),.I4(un1_write_addr_ptr_10[4:4]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1789));
defparam desc2944.INIT=64'hFFFF0000FFFD0200;
  LUT6_L desc2945(.I0(aresetn),.I1(N_1754),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(un1_write_addr_ptr_11[3:3]),.I4(un1_write_addr_ptr_10[3:3]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1788));
defparam desc2945.INIT=64'hFFFF0000FFFD0200;
  LUT6_L desc2946(.I0(aresetn),.I1(N_1754),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(un1_write_addr_ptr_11[2:2]),.I4(un1_write_addr_ptr_10[2:2]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1787));
defparam desc2946.INIT=64'hFFFF0000FFFD0200;
  LUT6_L desc2947(.I0(aresetn),.I1(N_1754),.I2(un1_write_addr_ptr_11[1:1]),.I3(un1_write_ram_ptr_0_sqmuxa),.I4(un1_write_addr_ptr_10[1:1]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1786));
defparam desc2947.INIT=64'hFFFF0000FFFD0020;
  LUT6_L desc2948(.I0(aresetn),.I1(N_1754),.I2(un1_write_addr_ptr_11[0:0]),.I3(un1_write_ram_ptr_0_sqmuxa),.I4(un1_write_addr_ptr_10[0:0]),.I5(write_ram_ptr_0_sqmuxa_1),.LO(N_1785));
defparam desc2948.INIT=64'hFFFF0000FFFD0020;
  LUT5 desc2949(.I0(window_length[6:6]),.I1(write_addr_ptr[6:6]),.I2(write_addr_ptr[4:4]),.I3(write_addr_ptr[5:5]),.I4(un9_s_axis_input_tvalid_a_4_c4),.O(un9_s_axis_input_tvalid_0_I_19_RNO));
defparam desc2949.INIT=32'h99996999;
  LUT5 desc2950(.I0(aresetn),.I1(N_1754),.I2(un9_s_axis_input_tvalid),.I3(un1_write_ram_ptr_0_sqmuxa),.I4(write_ram_ptr_0_sqmuxa_1),.O(un1_wen_ram_1_sqmuxa_1_i));
defparam desc2950.INIT=32'hF0FFF0DD;
  LUT4 desc2951(.I0(aresetn),.I1(un9_s_axis_input_tvalid),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(write_ram_ptr_0_sqmuxa_1),.O(un9_s_axis_input_tvalid_0_I_19_RNIN8NO));
defparam desc2951.INIT=16'hDF55;
  LUT2 desc2952(.I0(acquisition_length[0:0]),.I1(window_length[0:0]),.O(un64_m_axis_output_tready_a_5_axb_0));
defparam desc2952.INIT=4'h9;
  LUT5 desc2953(.I0(aresetn),.I1(s_axis_ctrl_tdata_0),.I2(s_axis_ctrl_tdata_16),.I3(write_addr_ptr[0:0]),.I4(N_1754),.O(un1_write_addr_ptr_axb_0));
defparam desc2953.INIT=32'h82D700FF;
  LUT4 un1_write_addr_ptr_cry_0_RNO(.I0(aresetn),.I1(s_axis_ctrl_tdata_0),.I2(write_addr_ptr[0:0]),.I3(N_1754),.O(un1_write_addr_ptr_2[6:6]));
defparam un1_write_addr_ptr_cry_0_RNO.INIT=16'h72F0;
  LUT5 desc2954(.I0(aresetn),.I1(s_axis_ctrl_tdata_0),.I2(s_axis_ctrl_tdata_16),.I3(write_addr_ptr[0:0]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_0));
defparam desc2954.INIT=32'hD782FF00;
  LUT3 un1_write_addr_ptr_0_cry_0_RNO_cZ(.I0(aresetn),.I1(s_axis_ctrl_tdata_16),.I2(N_1754),.O(un1_write_addr_ptr_0_cry_0_RNO));
defparam un1_write_addr_ptr_0_cry_0_RNO_cZ.INIT=8'h80;
  LUT5 desc2955(.I0(aresetn),.I1(s_axis_ctrl_tdata_1),.I2(s_axis_ctrl_tdata_17),.I3(write_addr_ptr[1:1]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_1));
defparam desc2955.INIT=32'hD782FF00;
  LUT3 desc2956(.I0(aresetn),.I1(s_axis_ctrl_tdata_17),.I2(N_1754),.O(write_ram_fsm_ns_0_a4_0_RNI314E[1:1]));
defparam desc2956.INIT=8'h80;
  LUT5 desc2957(.I0(aresetn),.I1(s_axis_ctrl_tdata_2),.I2(s_axis_ctrl_tdata_18),.I3(write_addr_ptr[2:2]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_2));
defparam desc2957.INIT=32'hD782FF00;
  LUT3 desc2958(.I0(aresetn),.I1(s_axis_ctrl_tdata_18),.I2(N_1754),.O(write_ram_fsm_ns_0_a4_0_RNI424E[1:1]));
defparam desc2958.INIT=8'h80;
  LUT5 desc2959(.I0(aresetn),.I1(s_axis_ctrl_tdata_3),.I2(s_axis_ctrl_tdata_19),.I3(write_addr_ptr[3:3]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_3));
defparam desc2959.INIT=32'hD782FF00;
  LUT3 desc2960(.I0(aresetn),.I1(s_axis_ctrl_tdata_19),.I2(N_1754),.O(write_ram_fsm_ns_0_a4_0_RNI534E[1:1]));
defparam desc2960.INIT=8'h80;
  LUT5 desc2961(.I0(aresetn),.I1(s_axis_ctrl_tdata_4),.I2(s_axis_ctrl_tdata_20),.I3(write_addr_ptr[4:4]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_4));
defparam desc2961.INIT=32'hD782FF00;
  LUT3 desc2962(.I0(aresetn),.I1(s_axis_ctrl_tdata_20),.I2(N_1754),.O(write_ram_fsm_ns_0_a4_0_RNITR4E[1:1]));
defparam desc2962.INIT=8'h80;
  LUT5 desc2963(.I0(aresetn),.I1(s_axis_ctrl_tdata_5),.I2(s_axis_ctrl_tdata_21),.I3(write_addr_ptr[5:5]),.I4(N_1754),.O(un1_write_addr_ptr_0_axb_5));
defparam desc2963.INIT=32'hD782FF00;
  LUT3 desc2964(.I0(aresetn),.I1(s_axis_ctrl_tdata_21),.I2(N_1754),.O(write_ram_fsm_ns_0_a4_0_RNIUS4E[1:1]));
defparam desc2964.INIT=8'h80;
  LUT5_L desc2965(.I0(read_last_addr_ptr_m_0[5:5]),.I1(un1_read_addr_ptr_1_1_sqmuxa_2_f0_0[6:6]),.I2(window_length_m_0[5:5]),.I3(read_addr_ptr_1_m[5:5]),.I4(un1_read_addr_ptr_1_1_sqmuxa_2_f1[6:6]),.LO(un1_read_addr_ptr_1_2_axb_5));
defparam desc2965.INIT=32'h3336FFFA;
  FDR desc2966(.Q(ram_window_tuser[1:1]),.D(m_axis_output_window_tuser_int_RNO[1:1]),.C(aclk),.R(aresetn_i));
  FDR desc2967(.Q(ram_window_tuser[0:0]),.D(m_axis_output_window_tuser_int_RNO[0:0]),.C(aclk),.R(aresetn_i));
  FDR desc2968(.Q(ram_tvalid[1:1]),.D(write_window_complete_RNIV26T_O6),.C(aclk),.R(aresetn_i));
  FDR desc2969(.Q(ram_tvalid[0:0]),.D(m_axis_output_tvalid_int_RNO),.C(aclk),.R(aresetn_i));
  XORCY un21_m_axis_output_tready_s_6_cZ(.LI(un21_m_axis_output_tready_axb_6),.CI(un21_m_axis_output_tready_cry_5),.O(un21_m_axis_output_tready_s_6));
  XORCY un21_m_axis_output_tready_s_5_cZ(.LI(un21_m_axis_output_tready_axb_5),.CI(un21_m_axis_output_tready_cry_4),.O(un21_m_axis_output_tready_s_5));
  MUXCY_L un21_m_axis_output_tready_cry_5_cZ(.DI(window_length[5:5]),.CI(un21_m_axis_output_tready_cry_4),.S(un21_m_axis_output_tready_axb_5),.LO(un21_m_axis_output_tready_cry_5));
  XORCY un21_m_axis_output_tready_s_4_cZ(.LI(un21_m_axis_output_tready_axb_4),.CI(un21_m_axis_output_tready_cry_3),.O(un21_m_axis_output_tready_s_4));
  MUXCY_L un21_m_axis_output_tready_cry_4_cZ(.DI(window_length[4:4]),.CI(un21_m_axis_output_tready_cry_3),.S(un21_m_axis_output_tready_axb_4),.LO(un21_m_axis_output_tready_cry_4));
  XORCY un21_m_axis_output_tready_s_3_cZ(.LI(un21_m_axis_output_tready_axb_3),.CI(un21_m_axis_output_tready_cry_2),.O(un21_m_axis_output_tready_s_3));
  MUXCY_L un21_m_axis_output_tready_cry_3_cZ(.DI(window_length[3:3]),.CI(un21_m_axis_output_tready_cry_2),.S(un21_m_axis_output_tready_axb_3),.LO(un21_m_axis_output_tready_cry_3));
  XORCY un21_m_axis_output_tready_s_2_cZ(.LI(un21_m_axis_output_tready_axb_2),.CI(un21_m_axis_output_tready_cry_1),.O(un21_m_axis_output_tready_s_2));
  MUXCY_L un21_m_axis_output_tready_cry_2_cZ(.DI(window_length[2:2]),.CI(un21_m_axis_output_tready_cry_1),.S(un21_m_axis_output_tready_axb_2),.LO(un21_m_axis_output_tready_cry_2));
  XORCY un21_m_axis_output_tready_s_1_cZ(.LI(un21_m_axis_output_tready_axb_1),.CI(un21_m_axis_output_tready_cry_0),.O(un21_m_axis_output_tready_s_1));
  MUXCY_L un21_m_axis_output_tready_cry_1_cZ(.DI(window_length[1:1]),.CI(un21_m_axis_output_tready_cry_0),.S(un21_m_axis_output_tready_axb_1),.LO(un21_m_axis_output_tready_cry_1));
  MUXCY_L un21_m_axis_output_tready_cry_0_cZ(.DI(window_length[0:0]),.CI(GND),.S(un21_m_axis_output_tready_axb_0),.LO(un21_m_axis_output_tready_cry_0));
  XORCY un1_read_addr_ptr_0_2_s_6_cZ(.LI(un1_read_addr_ptr_0_2_axb_6),.CI(un1_read_addr_ptr_0_2_cry_5),.O(un1_read_addr_ptr_0_2_s_6));
  XORCY un1_read_addr_ptr_0_2_s_5_cZ(.LI(un1_read_addr_ptr_0_2_axb_5),.CI(un1_read_addr_ptr_0_2_cry_4),.O(un1_read_addr_ptr_0_2_s_5));
  MUXCY_L un1_read_addr_ptr_0_2_cry_5_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(un1_read_addr_ptr_0_2_cry_4),.S(un1_read_addr_ptr_0_2_axb_5),.LO(un1_read_addr_ptr_0_2_cry_5));
  XORCY un1_read_addr_ptr_0_2_s_4_cZ(.LI(un1_read_addr_ptr_0_2_axb_4),.CI(un1_read_addr_ptr_0_2_cry_3),.O(un1_read_addr_ptr_0_2_s_4));
  MUXCY_L un1_read_addr_ptr_0_2_cry_4_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(un1_read_addr_ptr_0_2_cry_3),.S(un1_read_addr_ptr_0_2_axb_4),.LO(un1_read_addr_ptr_0_2_cry_4));
  XORCY un1_read_addr_ptr_0_2_s_3_cZ(.LI(un1_read_addr_ptr_0_2_axb_3),.CI(un1_read_addr_ptr_0_2_cry_2),.O(un1_read_addr_ptr_0_2_s_3));
  MUXCY_L un1_read_addr_ptr_0_2_cry_3_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(un1_read_addr_ptr_0_2_cry_2),.S(un1_read_addr_ptr_0_2_axb_3),.LO(un1_read_addr_ptr_0_2_cry_3));
  XORCY un1_read_addr_ptr_0_2_s_2_cZ(.LI(un1_read_addr_ptr_0_2_axb_2),.CI(un1_read_addr_ptr_0_2_cry_1),.O(un1_read_addr_ptr_0_2_s_2));
  MUXCY_L un1_read_addr_ptr_0_2_cry_2_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(un1_read_addr_ptr_0_2_cry_1),.S(un1_read_addr_ptr_0_2_axb_2),.LO(un1_read_addr_ptr_0_2_cry_2));
  XORCY un1_read_addr_ptr_0_2_s_1_cZ(.LI(un1_read_addr_ptr_0_2_axb_1),.CI(un1_read_addr_ptr_0_2_cry_0),.O(un1_read_addr_ptr_0_2_s_1));
  MUXCY_L un1_read_addr_ptr_0_2_cry_1_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(un1_read_addr_ptr_0_2_cry_0),.S(un1_read_addr_ptr_0_2_axb_1),.LO(un1_read_addr_ptr_0_2_cry_1));
  MUXCY_L un1_read_addr_ptr_0_2_cry_0_cZ(.DI(read_addr_ptr_0_1_sqmuxa_3_RNIVHT32),.CI(GND),.S(un1_read_addr_ptr_0_2_cry_0_RNO),.LO(un1_read_addr_ptr_0_2_cry_0));
  XORCY un1_read_addr_ptr_1_2_s_6_cZ(.LI(un1_read_addr_ptr_1_2_axb_6),.CI(un1_read_addr_ptr_1_2_cry_5),.O(un1_read_addr_ptr_1_2_s_6));
  XORCY un1_read_addr_ptr_1_2_s_5_cZ(.LI(un1_read_addr_ptr_1_2_axb_5),.CI(un1_read_addr_ptr_1_2_cry_4),.O(un1_read_addr_ptr_1_2_s_5));
  MUXCY_L un1_read_addr_ptr_1_2_cry_5_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(un1_read_addr_ptr_1_2_cry_4),.S(un1_read_addr_ptr_1_2_axb_5),.LO(un1_read_addr_ptr_1_2_cry_5));
  XORCY un1_read_addr_ptr_1_2_s_4_cZ(.LI(un1_read_addr_ptr_1_2_axb_4),.CI(un1_read_addr_ptr_1_2_cry_3),.O(un1_read_addr_ptr_1_2_s_4));
  MUXCY_L un1_read_addr_ptr_1_2_cry_4_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(un1_read_addr_ptr_1_2_cry_3),.S(un1_read_addr_ptr_1_2_axb_4),.LO(un1_read_addr_ptr_1_2_cry_4));
  XORCY un1_read_addr_ptr_1_2_s_3_cZ(.LI(un1_read_addr_ptr_1_2_axb_3),.CI(un1_read_addr_ptr_1_2_cry_2),.O(un1_read_addr_ptr_1_2_s_3));
  MUXCY_L un1_read_addr_ptr_1_2_cry_3_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(un1_read_addr_ptr_1_2_cry_2),.S(un1_read_addr_ptr_1_2_axb_3),.LO(un1_read_addr_ptr_1_2_cry_3));
  XORCY un1_read_addr_ptr_1_2_s_2_cZ(.LI(un1_read_addr_ptr_1_2_axb_2),.CI(un1_read_addr_ptr_1_2_cry_1),.O(un1_read_addr_ptr_1_2_s_2));
  MUXCY_L un1_read_addr_ptr_1_2_cry_2_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(un1_read_addr_ptr_1_2_cry_1),.S(un1_read_addr_ptr_1_2_axb_2),.LO(un1_read_addr_ptr_1_2_cry_2));
  XORCY un1_read_addr_ptr_1_2_s_1_cZ(.LI(un1_read_addr_ptr_1_2_axb_1),.CI(un1_read_addr_ptr_1_2_cry_0),.O(un1_read_addr_ptr_1_2_s_1));
  MUXCY_L un1_read_addr_ptr_1_2_cry_1_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(un1_read_addr_ptr_1_2_cry_0),.S(un1_read_addr_ptr_1_2_axb_1),.LO(un1_read_addr_ptr_1_2_cry_1));
  MUXCY_L un1_read_addr_ptr_1_2_cry_0_cZ(.DI(read_addr_ptr_1_2_sqmuxa_1_RNIRVDQ),.CI(GND),.S(un1_read_addr_ptr_1_2_cry_0_RNO),.LO(un1_read_addr_ptr_1_2_cry_0));
  XORCY desc2970(.LI(un18_m_axis_output_tready_axb_6),.CI(un18_m_axis_output_tready_cry_5),.O(un18_m_axis_output_tready[6:6]));
  XORCY desc2971(.LI(un18_m_axis_output_tready_axb_5),.CI(un18_m_axis_output_tready_cry_4),.O(un18_m_axis_output_tready[5:5]));
  MUXCY_L desc2972(.DI(window_length[5:5]),.CI(un18_m_axis_output_tready_cry_4),.S(un18_m_axis_output_tready_axb_5),.LO(un18_m_axis_output_tready_cry_5));
  XORCY desc2973(.LI(un18_m_axis_output_tready_axb_4),.CI(un18_m_axis_output_tready_cry_3),.O(un18_m_axis_output_tready[4:4]));
  MUXCY_L desc2974(.DI(window_length[4:4]),.CI(un18_m_axis_output_tready_cry_3),.S(un18_m_axis_output_tready_axb_4),.LO(un18_m_axis_output_tready_cry_4));
  XORCY desc2975(.LI(un18_m_axis_output_tready_axb_3),.CI(un18_m_axis_output_tready_cry_2),.O(un18_m_axis_output_tready[3:3]));
  MUXCY_L desc2976(.DI(window_length[3:3]),.CI(un18_m_axis_output_tready_cry_2),.S(un18_m_axis_output_tready_axb_3),.LO(un18_m_axis_output_tready_cry_3));
  XORCY desc2977(.LI(un18_m_axis_output_tready_axb_2),.CI(un18_m_axis_output_tready_cry_1),.O(un18_m_axis_output_tready[2:2]));
  MUXCY_L desc2978(.DI(window_length[2:2]),.CI(un18_m_axis_output_tready_cry_1),.S(un18_m_axis_output_tready_axb_2),.LO(un18_m_axis_output_tready_cry_2));
  XORCY desc2979(.LI(un18_m_axis_output_tready_axb_1),.CI(un18_m_axis_output_tready_cry_0),.O(un18_m_axis_output_tready[1:1]));
  MUXCY_L desc2980(.DI(window_length[1:1]),.CI(un18_m_axis_output_tready_cry_0),.S(un18_m_axis_output_tready_axb_1),.LO(un18_m_axis_output_tready_cry_1));
  MUXCY_L desc2981(.DI(window_length_fast[0:0]),.CI(VCC),.S(un18_m_axis_output_tready_cry_0_RNO),.LO(un18_m_axis_output_tready_cry_0));
  XORCY un1_write_addr_ptr_0_s_6(.LI(un1_write_addr_ptr_0_axb_6),.CI(un1_write_addr_ptr_0_cry_5),.O(un1_write_addr_ptr_11[6:6]));
  XORCY un1_write_addr_ptr_0_s_5(.LI(un1_write_addr_ptr_0_axb_5),.CI(un1_write_addr_ptr_0_cry_4),.O(un1_write_addr_ptr_11[5:5]));
  MUXCY_L un1_write_addr_ptr_0_cry_5_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNIUS4E[1:1]),.CI(un1_write_addr_ptr_0_cry_4),.S(un1_write_addr_ptr_0_axb_5),.LO(un1_write_addr_ptr_0_cry_5));
  XORCY un1_write_addr_ptr_0_s_4(.LI(un1_write_addr_ptr_0_axb_4),.CI(un1_write_addr_ptr_0_cry_3),.O(un1_write_addr_ptr_11[4:4]));
  MUXCY_L un1_write_addr_ptr_0_cry_4_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNITR4E[1:1]),.CI(un1_write_addr_ptr_0_cry_3),.S(un1_write_addr_ptr_0_axb_4),.LO(un1_write_addr_ptr_0_cry_4));
  XORCY un1_write_addr_ptr_0_s_3(.LI(un1_write_addr_ptr_0_axb_3),.CI(un1_write_addr_ptr_0_cry_2),.O(un1_write_addr_ptr_11[3:3]));
  MUXCY_L un1_write_addr_ptr_0_cry_3_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI534E[1:1]),.CI(un1_write_addr_ptr_0_cry_2),.S(un1_write_addr_ptr_0_axb_3),.LO(un1_write_addr_ptr_0_cry_3));
  XORCY un1_write_addr_ptr_0_s_2(.LI(un1_write_addr_ptr_0_axb_2),.CI(un1_write_addr_ptr_0_cry_1),.O(un1_write_addr_ptr_11[2:2]));
  MUXCY_L un1_write_addr_ptr_0_cry_2_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI424E[1:1]),.CI(un1_write_addr_ptr_0_cry_1),.S(un1_write_addr_ptr_0_axb_2),.LO(un1_write_addr_ptr_0_cry_2));
  XORCY un1_write_addr_ptr_0_s_1(.LI(un1_write_addr_ptr_0_axb_1),.CI(un1_write_addr_ptr_0_cry_0),.O(un1_write_addr_ptr_11[1:1]));
  MUXCY_L un1_write_addr_ptr_0_cry_1_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI314E[1:1]),.CI(un1_write_addr_ptr_0_cry_0),.S(un1_write_addr_ptr_0_axb_1),.LO(un1_write_addr_ptr_0_cry_1));
  XORCY un1_write_addr_ptr_0_s_0(.LI(un1_write_addr_ptr_0_axb_0),.CI(un1_write_addr_ptr_0_cry_0_cy),.O(un1_write_addr_ptr_11[0:0]));
  MUXCY_L un1_write_addr_ptr_0_cry_0_cZ(.DI(un1_write_addr_ptr_0_cry_0_RNO),.CI(un1_write_addr_ptr_0_cry_0_cy),.S(un1_write_addr_ptr_0_axb_0),.LO(un1_write_addr_ptr_0_cry_0));
  XORCY un1_write_addr_ptr_s_6(.LI(un1_write_addr_ptr_axb_6),.CI(un1_write_addr_ptr_cry_5),.O(un1_write_addr_ptr_10[6:6]));
  XORCY un1_write_addr_ptr_s_5(.LI(un1_write_addr_ptr_axb_5),.CI(un1_write_addr_ptr_cry_4),.O(un1_write_addr_ptr_10[5:5]));
  MUXCY_L un1_write_addr_ptr_cry_5_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNIUS4E[1:1]),.CI(un1_write_addr_ptr_cry_4),.S(un1_write_addr_ptr_axb_5),.LO(un1_write_addr_ptr_cry_5));
  XORCY un1_write_addr_ptr_s_4(.LI(un1_write_addr_ptr_axb_4),.CI(un1_write_addr_ptr_cry_3),.O(un1_write_addr_ptr_10[4:4]));
  MUXCY_L un1_write_addr_ptr_cry_4_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNITR4E[1:1]),.CI(un1_write_addr_ptr_cry_3),.S(un1_write_addr_ptr_axb_4),.LO(un1_write_addr_ptr_cry_4));
  XORCY un1_write_addr_ptr_s_3(.LI(un1_write_addr_ptr_axb_3),.CI(un1_write_addr_ptr_cry_2),.O(un1_write_addr_ptr_10[3:3]));
  MUXCY_L un1_write_addr_ptr_cry_3_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI534E[1:1]),.CI(un1_write_addr_ptr_cry_2),.S(un1_write_addr_ptr_axb_3),.LO(un1_write_addr_ptr_cry_3));
  XORCY un1_write_addr_ptr_s_2(.LI(un1_write_addr_ptr_axb_2),.CI(un1_write_addr_ptr_cry_1),.O(un1_write_addr_ptr_10[2:2]));
  MUXCY_L un1_write_addr_ptr_cry_2_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI424E[1:1]),.CI(un1_write_addr_ptr_cry_1),.S(un1_write_addr_ptr_axb_2),.LO(un1_write_addr_ptr_cry_2));
  XORCY un1_write_addr_ptr_s_1(.LI(un1_write_addr_ptr_axb_1),.CI(un1_write_addr_ptr_cry_0),.O(un1_write_addr_ptr_10[1:1]));
  MUXCY_L un1_write_addr_ptr_cry_1_cZ(.DI(write_ram_fsm_ns_0_a4_0_RNI314E[1:1]),.CI(un1_write_addr_ptr_cry_0),.S(un1_write_addr_ptr_axb_1),.LO(un1_write_addr_ptr_cry_1));
  XORCY un1_write_addr_ptr_s_0(.LI(un1_write_addr_ptr_axb_0),.CI(un1_write_addr_ptr_cry_0_cy),.O(un1_write_addr_ptr_10[0:0]));
  MUXCY_L un1_write_addr_ptr_cry_0_cZ(.DI(un1_write_addr_ptr_2[6:6]),.CI(un1_write_addr_ptr_cry_0_cy),.S(un1_write_addr_ptr_axb_0),.LO(un1_write_addr_ptr_cry_0));
  XORCY desc2982(.LI(un64_m_axis_output_tready_a_5_axb_6),.CI(un64_m_axis_output_tready_a_5_cry_5),.O(un64_m_axis_output_tready_a_5[6:6]));
  XORCY desc2983(.LI(un64_m_axis_output_tready_a_5_axb_5),.CI(un64_m_axis_output_tready_a_5_cry_4),.O(un64_m_axis_output_tready_a_5[5:5]));
  MUXCY_L desc2984(.DI(window_length[5:5]),.CI(un64_m_axis_output_tready_a_5_cry_4),.S(un64_m_axis_output_tready_a_5_axb_5),.LO(un64_m_axis_output_tready_a_5_cry_5));
  XORCY desc2985(.LI(un64_m_axis_output_tready_a_5_axb_4),.CI(un64_m_axis_output_tready_a_5_cry_3),.O(un64_m_axis_output_tready_a_5[4:4]));
  MUXCY_L desc2986(.DI(window_length_fast[4:4]),.CI(un64_m_axis_output_tready_a_5_cry_3),.S(un64_m_axis_output_tready_a_5_axb_4),.LO(un64_m_axis_output_tready_a_5_cry_4));
  XORCY desc2987(.LI(un64_m_axis_output_tready_a_5_axb_3),.CI(un64_m_axis_output_tready_a_5_cry_2),.O(un64_m_axis_output_tready_a_5[3:3]));
  MUXCY_L desc2988(.DI(window_length_fast[3:3]),.CI(un64_m_axis_output_tready_a_5_cry_2),.S(un64_m_axis_output_tready_a_5_axb_3),.LO(un64_m_axis_output_tready_a_5_cry_3));
  XORCY desc2989(.LI(un64_m_axis_output_tready_a_5_axb_2),.CI(un64_m_axis_output_tready_a_5_cry_1),.O(un64_m_axis_output_tready_a_5[2:2]));
  MUXCY_L desc2990(.DI(window_length_fast[2:2]),.CI(un64_m_axis_output_tready_a_5_cry_1),.S(un64_m_axis_output_tready_a_5_axb_2),.LO(un64_m_axis_output_tready_a_5_cry_2));
  XORCY desc2991(.LI(un64_m_axis_output_tready_a_5_axb_1),.CI(un64_m_axis_output_tready_a_5_cry_0),.O(un64_m_axis_output_tready_a_5[1:1]));
  MUXCY_L desc2992(.DI(window_length_fast[1:1]),.CI(un64_m_axis_output_tready_a_5_cry_0),.S(un64_m_axis_output_tready_a_5_axb_1),.LO(un64_m_axis_output_tready_a_5_cry_1));
  MUXCY_L desc2993(.DI(window_length_fast[0:0]),.CI(VCC),.S(un64_m_axis_output_tready_a_5_cry_0_RNO),.LO(un64_m_axis_output_tready_a_5_cry_0));
  MUXCY_L desc2994(.DI(GND),.CI(un57_m_axis_output_tready_0_data_tmp[0:0]),.S(un57_m_axis_output_tready_0_N_4),.LO(un57_m_axis_output_tready_0_data_tmp[1:1]));
  MUXCY_L desc2995(.DI(GND),.CI(VCC),.S(un57_m_axis_output_tready_0_N_11),.LO(un57_m_axis_output_tready_0_data_tmp[0:0]));
  MUXCY_L desc2996(.DI(GND),.CI(un23_m_axis_output_tready_0_data_tmp[0:0]),.S(un23_m_axis_output_tready_0_N_4),.LO(un23_m_axis_output_tready_0_data_tmp[1:1]));
  MUXCY_L desc2997(.DI(GND),.CI(VCC),.S(un23_m_axis_output_tready_0_N_11),.LO(un23_m_axis_output_tready_0_data_tmp[0:0]));
  MUXCY_L desc2998(.DI(GND),.CI(un64_m_axis_output_tready_0_data_tmp[0:0]),.S(un64_m_axis_output_tready_0_N_4),.LO(un64_m_axis_output_tready_0_data_tmp[1:1]));
  MUXCY_L desc2999(.DI(GND),.CI(VCC),.S(un64_m_axis_output_tready_0_N_11),.LO(un64_m_axis_output_tready_0_data_tmp[0:0]));
  MUXCY_L desc3000(.DI(GND),.CI(un30_m_axis_output_tready_0_data_tmp[0:0]),.S(un30_m_axis_output_tready_0_N_4),.LO(un30_m_axis_output_tready_0_data_tmp[1:1]));
  MUXCY_L desc3001(.DI(GND),.CI(VCC),.S(un30_m_axis_output_tready_0_N_11),.LO(un30_m_axis_output_tready_0_data_tmp[0:0]));
  MUXCY_L desc3002(.DI(GND),.CI(un9_s_axis_input_tvalid_0_data_tmp[0:0]),.S(un9_s_axis_input_tvalid_0_N_4),.LO(un9_s_axis_input_tvalid_0_data_tmp[1:1]));
  MUXCY_L desc3003(.DI(GND),.CI(VCC),.S(un9_s_axis_input_tvalid_0_N_11),.LO(un9_s_axis_input_tvalid_0_data_tmp[0:0]));
  FDRE desc3004(.Q(ram_buffer_0[63:63]),.D(ram_buffer_0_2[63:63]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3005(.Q(ram_buffer_0[62:62]),.D(ram_buffer_0_2[62:62]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3006(.Q(ram_buffer_0[61:61]),.D(ram_buffer_0_2[61:61]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3007(.Q(ram_buffer_0[60:60]),.D(ram_buffer_0_2[60:60]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3008(.Q(ram_buffer_0[59:59]),.D(ram_buffer_0_2[59:59]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3009(.Q(ram_buffer_0[58:58]),.D(ram_buffer_0_2[58:58]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3010(.Q(ram_buffer_0[57:57]),.D(ram_buffer_0_2[57:57]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3011(.Q(ram_buffer_0[56:56]),.D(ram_buffer_0_2[56:56]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3012(.Q(ram_buffer_0[55:55]),.D(ram_buffer_0_2[55:55]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3013(.Q(ram_buffer_0[54:54]),.D(ram_buffer_0_2[54:54]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3014(.Q(ram_buffer_0[53:53]),.D(ram_buffer_0_2[53:53]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3015(.Q(ram_buffer_0[52:52]),.D(ram_buffer_0_2[52:52]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3016(.Q(ram_buffer_0[51:51]),.D(ram_buffer_0_2[51:51]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3017(.Q(ram_buffer_0[50:50]),.D(ram_buffer_0_2[50:50]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3018(.Q(ram_buffer_0[49:49]),.D(ram_buffer_0_2[49:49]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3019(.Q(ram_buffer_0[48:48]),.D(ram_buffer_0_2[48:48]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3020(.Q(ram_buffer_0[47:47]),.D(ram_buffer_0_2[47:47]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3021(.Q(ram_buffer_0[46:46]),.D(ram_buffer_0_2[46:46]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3022(.Q(ram_buffer_0[45:45]),.D(ram_buffer_0_2[45:45]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3023(.Q(ram_buffer_0[44:44]),.D(ram_buffer_0_2[44:44]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3024(.Q(ram_buffer_0[43:43]),.D(ram_buffer_0_2[43:43]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3025(.Q(ram_buffer_0[42:42]),.D(ram_buffer_0_2[42:42]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3026(.Q(ram_buffer_0[41:41]),.D(ram_buffer_0_2[41:41]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3027(.Q(ram_buffer_0[40:40]),.D(ram_buffer_0_2[40:40]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3028(.Q(ram_buffer_0[39:39]),.D(ram_buffer_0_2[39:39]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3029(.Q(ram_buffer_0[38:38]),.D(ram_buffer_0_2[38:38]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3030(.Q(ram_buffer_0[37:37]),.D(ram_buffer_0_2[37:37]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3031(.Q(ram_buffer_0[36:36]),.D(ram_buffer_0_2[36:36]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3032(.Q(ram_buffer_0[35:35]),.D(ram_buffer_0_2[35:35]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3033(.Q(ram_buffer_0[34:34]),.D(ram_buffer_0_2[34:34]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3034(.Q(ram_buffer_0[33:33]),.D(ram_buffer_0_2[33:33]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3035(.Q(ram_buffer_0[32:32]),.D(ram_buffer_0_2[32:32]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3036(.Q(ram_buffer_0[31:31]),.D(ram_buffer_0_2[31:31]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3037(.Q(ram_buffer_0[30:30]),.D(ram_buffer_0_2[30:30]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3038(.Q(ram_buffer_0[29:29]),.D(ram_buffer_0_2[29:29]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3039(.Q(ram_buffer_0[28:28]),.D(ram_buffer_0_2[28:28]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3040(.Q(ram_buffer_0[27:27]),.D(ram_buffer_0_2[27:27]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3041(.Q(ram_buffer_0[26:26]),.D(ram_buffer_0_2[26:26]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3042(.Q(ram_buffer_0[25:25]),.D(ram_buffer_0_2[25:25]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3043(.Q(ram_buffer_0[24:24]),.D(ram_buffer_0_2[24:24]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3044(.Q(ram_buffer_0[23:23]),.D(ram_buffer_0_2[23:23]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3045(.Q(ram_buffer_0[22:22]),.D(ram_buffer_0_2[22:22]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3046(.Q(ram_buffer_0[21:21]),.D(ram_buffer_0_2[21:21]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3047(.Q(ram_buffer_0[20:20]),.D(ram_buffer_0_2[20:20]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3048(.Q(ram_buffer_0[19:19]),.D(ram_buffer_0_2[19:19]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3049(.Q(ram_buffer_0[18:18]),.D(ram_buffer_0_2[18:18]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3050(.Q(ram_buffer_0[17:17]),.D(ram_buffer_0_2[17:17]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3051(.Q(ram_buffer_0[16:16]),.D(ram_buffer_0_2[16:16]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3052(.Q(ram_buffer_0[15:15]),.D(ram_buffer_0_2[15:15]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3053(.Q(ram_buffer_0[14:14]),.D(ram_buffer_0_2[14:14]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3054(.Q(ram_buffer_0[13:13]),.D(ram_buffer_0_2[13:13]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3055(.Q(ram_buffer_0[12:12]),.D(ram_buffer_0_2[12:12]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3056(.Q(ram_buffer_0[11:11]),.D(ram_buffer_0_2[11:11]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3057(.Q(ram_buffer_0[10:10]),.D(ram_buffer_0_2[10:10]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3058(.Q(ram_buffer_0[9:9]),.D(ram_buffer_0_2[9:9]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3059(.Q(ram_buffer_0[8:8]),.D(ram_buffer_0_2[8:8]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3060(.Q(ram_buffer_0[7:7]),.D(ram_buffer_0_2[7:7]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3061(.Q(ram_buffer_0[6:6]),.D(ram_buffer_0_2[6:6]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3062(.Q(ram_buffer_0[5:5]),.D(ram_buffer_0_2[5:5]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3063(.Q(ram_buffer_0[4:4]),.D(ram_buffer_0_2[4:4]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3064(.Q(ram_buffer_0[3:3]),.D(ram_buffer_0_2[3:3]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3065(.Q(ram_buffer_0[2:2]),.D(ram_buffer_0_2[2:2]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3066(.Q(ram_buffer_0[1:1]),.D(ram_buffer_0_2[1:1]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3067(.Q(ram_buffer_0[0:0]),.D(ram_buffer_0_2[0:0]),.C(aclk),.R(aresetn_i),.CE(un5_m_axis_output_tvalid_int));
  FDRE desc3068(.Q(ram_buffer_1[63:63]),.D(ram_buffer_1_1[63:63]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3069(.Q(ram_buffer_1[62:62]),.D(ram_buffer_1_1[62:62]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3070(.Q(ram_buffer_1[61:61]),.D(ram_buffer_1_1[61:61]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3071(.Q(ram_buffer_1[60:60]),.D(ram_buffer_1_1[60:60]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3072(.Q(ram_buffer_1[59:59]),.D(ram_buffer_1_1[59:59]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3073(.Q(ram_buffer_1[58:58]),.D(ram_buffer_1_1[58:58]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3074(.Q(ram_buffer_1[57:57]),.D(ram_buffer_1_1[57:57]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3075(.Q(ram_buffer_1[56:56]),.D(ram_buffer_1_1[56:56]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3076(.Q(ram_buffer_1[55:55]),.D(ram_buffer_1_1[55:55]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3077(.Q(ram_buffer_1[54:54]),.D(ram_buffer_1_1[54:54]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3078(.Q(ram_buffer_1[53:53]),.D(ram_buffer_1_1[53:53]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3079(.Q(ram_buffer_1[52:52]),.D(ram_buffer_1_1[52:52]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3080(.Q(ram_buffer_1[51:51]),.D(ram_buffer_1_1[51:51]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3081(.Q(ram_buffer_1[50:50]),.D(ram_buffer_1_1[50:50]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3082(.Q(ram_buffer_1[49:49]),.D(ram_buffer_1_1[49:49]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3083(.Q(ram_buffer_1[48:48]),.D(ram_buffer_1_1[48:48]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3084(.Q(ram_buffer_1[47:47]),.D(ram_buffer_1_1[47:47]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3085(.Q(ram_buffer_1[46:46]),.D(ram_buffer_1_1[46:46]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3086(.Q(ram_buffer_1[45:45]),.D(ram_buffer_1_1[45:45]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3087(.Q(ram_buffer_1[44:44]),.D(ram_buffer_1_1[44:44]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3088(.Q(ram_buffer_1[43:43]),.D(ram_buffer_1_1[43:43]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3089(.Q(ram_buffer_1[42:42]),.D(ram_buffer_1_1[42:42]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3090(.Q(ram_buffer_1[41:41]),.D(ram_buffer_1_1[41:41]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3091(.Q(ram_buffer_1[40:40]),.D(ram_buffer_1_1[40:40]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3092(.Q(ram_buffer_1[39:39]),.D(ram_buffer_1_1[39:39]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3093(.Q(ram_buffer_1[38:38]),.D(ram_buffer_1_1[38:38]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3094(.Q(ram_buffer_1[37:37]),.D(ram_buffer_1_1[37:37]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3095(.Q(ram_buffer_1[36:36]),.D(ram_buffer_1_1[36:36]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3096(.Q(ram_buffer_1[35:35]),.D(ram_buffer_1_1[35:35]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3097(.Q(ram_buffer_1[34:34]),.D(ram_buffer_1_1[34:34]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3098(.Q(ram_buffer_1[33:33]),.D(ram_buffer_1_1[33:33]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3099(.Q(ram_buffer_1[32:32]),.D(ram_buffer_1_1[32:32]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3100(.Q(ram_buffer_1[31:31]),.D(ram_buffer_1_1[31:31]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3101(.Q(ram_buffer_1[30:30]),.D(ram_buffer_1_1[30:30]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3102(.Q(ram_buffer_1[29:29]),.D(ram_buffer_1_1[29:29]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3103(.Q(ram_buffer_1[28:28]),.D(ram_buffer_1_1[28:28]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3104(.Q(ram_buffer_1[27:27]),.D(ram_buffer_1_1[27:27]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3105(.Q(ram_buffer_1[26:26]),.D(ram_buffer_1_1[26:26]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3106(.Q(ram_buffer_1[25:25]),.D(ram_buffer_1_1[25:25]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3107(.Q(ram_buffer_1[24:24]),.D(ram_buffer_1_1[24:24]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3108(.Q(ram_buffer_1[23:23]),.D(ram_buffer_1_1[23:23]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3109(.Q(ram_buffer_1[22:22]),.D(ram_buffer_1_1[22:22]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3110(.Q(ram_buffer_1[21:21]),.D(ram_buffer_1_1[21:21]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3111(.Q(ram_buffer_1[20:20]),.D(ram_buffer_1_1[20:20]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3112(.Q(ram_buffer_1[19:19]),.D(ram_buffer_1_1[19:19]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3113(.Q(ram_buffer_1[18:18]),.D(ram_buffer_1_1[18:18]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3114(.Q(ram_buffer_1[17:17]),.D(ram_buffer_1_1[17:17]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3115(.Q(ram_buffer_1[16:16]),.D(ram_buffer_1_1[16:16]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3116(.Q(ram_buffer_1[15:15]),.D(ram_buffer_1_1[15:15]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3117(.Q(ram_buffer_1[14:14]),.D(ram_buffer_1_1[14:14]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3118(.Q(ram_buffer_1[13:13]),.D(ram_buffer_1_1[13:13]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3119(.Q(ram_buffer_1[12:12]),.D(ram_buffer_1_1[12:12]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3120(.Q(ram_buffer_1[11:11]),.D(ram_buffer_1_1[11:11]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3121(.Q(ram_buffer_1[10:10]),.D(ram_buffer_1_1[10:10]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3122(.Q(ram_buffer_1[9:9]),.D(ram_buffer_1_1[9:9]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3123(.Q(ram_buffer_1[8:8]),.D(ram_buffer_1_1[8:8]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3124(.Q(ram_buffer_1[7:7]),.D(ram_buffer_1_1[7:7]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3125(.Q(ram_buffer_1[6:6]),.D(ram_buffer_1_1[6:6]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3126(.Q(ram_buffer_1[5:5]),.D(ram_buffer_1_1[5:5]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3127(.Q(ram_buffer_1[4:4]),.D(ram_buffer_1_1[4:4]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3128(.Q(ram_buffer_1[3:3]),.D(ram_buffer_1_1[3:3]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3129(.Q(ram_buffer_1[2:2]),.D(ram_buffer_1_1[2:2]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3130(.Q(ram_buffer_1[1:1]),.D(ram_buffer_1_1[1:1]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3131(.Q(ram_buffer_1[0:0]),.D(ram_buffer_1_1[0:0]),.C(aclk),.R(aresetn_i),.CE(un21_m_axis_output_tvalid_int));
  FDRE desc3132(.Q(read_last_addr_ptr[6:6]),.D(write_addr_ptr[6:6]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3133(.Q(read_last_addr_ptr[5:5]),.D(write_addr_ptr[5:5]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3134(.Q(read_last_addr_ptr[4:4]),.D(write_addr_ptr[4:4]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3135(.Q(read_last_addr_ptr[3:3]),.D(write_addr_ptr[3:3]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3136(.Q(read_last_addr_ptr[2:2]),.D(write_addr_ptr[2:2]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3137(.Q(read_last_addr_ptr[1:1]),.D(write_addr_ptr[1:1]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDRE desc3138(.Q(read_last_addr_ptr[0:0]),.D(write_addr_ptr[0:0]),.C(aclk),.R(aresetn_i),.CE(write_ram_ptr_0_sqmuxa_1));
  FDR desc3139(.Q(read_ram_ptr_d_0[1:1]),.D(read_ram_ptr_0[1:1]),.C(aclk),.R(aresetn_i));
  FDR desc3140(.Q(read_ram_ptr_d_0[0:0]),.D(read_ram_ptr_0[0:0]),.C(aclk),.R(aresetn_i));
  FDR desc3141(.Q(read_ram_ptr_d_1[1:1]),.D(read_ram_ptr_1[1:1]),.C(aclk),.R(aresetn_i));
  FDR desc3142(.Q(read_ram_ptr_d_1[0:0]),.D(read_ram_ptr_1[0:0]),.C(aclk),.R(aresetn_i));
  generic_sp_ram_inj desc3143(.q_reg_1(q_reg_1[63:0]),.addr_1(addr_1[6:0]),.acs_dec_tdata(acs_dec_tdata[63:0]),.wen_ram(wen_ram[1:1]),.aclk(aclk));
  generic_sp_ram_1_inj desc3144(.q_reg_2(q_reg_2[63:0]),.addr_2(addr_2[6:0]),.acs_dec_tdata(acs_dec_tdata[63:0]),.wen_ram(wen_ram[2:2]),.aclk(aclk));
  generic_sp_ram_2_inj desc3145(.q_reg_3(q_reg_3[63:0]),.addr_3(addr_3[6:0]),.acs_dec_tdata(acs_dec_tdata[63:0]),.wen_ram(wen_ram[3:3]),.aclk(aclk));
  generic_sp_ram_3_inj desc3146(.q_reg_0(q_reg_0[63:0]),.addr_0(addr_0[6:0]),.acs_dec_tdata(acs_dec_tdata[63:0]),.wen_ram(wen_ram[0:0]),.aclk(aclk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT5 desc3147(.I0(un1_s_axis_input_tvalid),.I1(un9_s_axis_input_tvalid),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(write_ram_ptr[1:1]),.I4(write_ram_ptr[0:0]),.O(SUM1_5));
defparam desc3147.INIT=32'h758AFF00;
  LUT4 desc3148(.I0(un1_s_axis_input_tvalid),.I1(un9_s_axis_input_tvalid),.I2(un1_write_ram_ptr_0_sqmuxa),.I3(write_ram_ptr[0:0]),.O(N_2332_i_0));
defparam desc3148.INIT=16'h758A;
  LUT4 desc3149(.I0(read_ram_fsm_0[1:1]),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(read_ram_fsm_0[0:0]),.O(N_1731));
defparam desc3149.INIT=16'h0357;
  LUT5 desc3150(.I0(read_ram_fsm_0[1:1]),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(read_ram_fsm_0[0:0]),.I4(write_ram_fsm_1),.O(write_ram_fsm_1_sqmuxa));
defparam desc3150.INIT=32'hFCA80000;
  LUT4 un1_write_ram_ptr_0_sqmuxa_sx_lut6_2_o6(.I0(write_ram_fsm_fast[0:0]),.I1(write_ram_fsm_fast[4:4]),.I2(write_ram_fsm[3:3]),.I3(acs_tlast),.O(un1_write_ram_ptr_0_sqmuxa_sx));
defparam un1_write_ram_ptr_0_sqmuxa_sx_lut6_2_o6.INIT=16'hEFEE;
  LUT2 un1_write_ram_ptr_0_sqmuxa_sx_lut6_2_o5(.I0(acs_tlast),.I1(write_ram_fsm[2:2]),.O(N_1739));
defparam un1_write_ram_ptr_0_sqmuxa_sx_lut6_2_o5.INIT=4'hB;
  LUT2 desc3151(.I0(write_last_window_complete),.I1(next_traceback),.O(un13_write_last_window_complete));
defparam desc3151.INIT=4'h2;
  LUT5 desc3152(.I0(ram_window_tuser[1:1]),.I1(write_last_window_complete),.I2(read_ram_fsm_1[0:0]),.I3(read_ram_fsm_1[1:1]),.I4(next_traceback),.O(un1_m_axis_output_window_tuser_int_0_sqmuxa_set_0));
defparam desc3152.INIT=32'hAAACAAA0;
  LUT2 desc3153(.I0(read_ram_fsm_0_0_rep1),.I1(read_ram_fsm_0_1_rep1),.O(read_ram_fsm_0_d_i_0[3:3]));
defparam desc3153.INIT=4'hE;
  LUT5 desc3154(.I0(read_ram_fsm_0_0_rep1),.I1(read_ram_fsm_0_1_rep1),.I2(write_window_complete),.I3(write_last_window_complete),.I4(next_traceback),.O(read_addr_ptr_0_1_sqmuxa_1));
defparam desc3154.INIT=32'h00000010;
  LUT2 desc3155(.I0(acs_tvalid),.I1(un9_s_axis_input_tvalid),.O(N_1740));
defparam desc3155.INIT=4'h7;
  LUT4 desc3156(.I0(un1_write_ram_ptr_0_sqmuxa),.I1(write_ram_ptr_fast[0:0]),.I2(un1_s_axis_input_tvalid),.I3(un9_s_axis_input_tvalid),.O(N_2332_i_fast_0));
defparam desc3156.INIT=16'h3C9C;
  LUT3 m_axis_output_tlast_int_0_sqmuxa_0_lut6_2_o6(.I0(last_of_block),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.O(m_axis_output_tlast_int_0_sqmuxa_0));
defparam m_axis_output_tlast_int_0_sqmuxa_0_lut6_2_o6.INIT=8'h02;
  LUT2 m_axis_output_tlast_int_0_sqmuxa_0_lut6_2_o5(.I0(last_of_block),.I1(acs_tlast),.O(last_of_block_0));
defparam m_axis_output_tlast_int_0_sqmuxa_0_lut6_2_o5.INIT=4'hE;
  LUT4 desc3157(.I0(write_ram_ptr[1:1]),.I1(write_ram_ptr[0:0]),.I2(write_ram_fsm[3:3]),.I3(write_ram_fsm[2:2]),.O(un3_addr));
defparam desc3157.INIT=16'h1110;
  LUT4 desc3158(.I0(write_ram_ptr[1:1]),.I1(write_ram_ptr[0:0]),.I2(write_ram_fsm[3:3]),.I3(write_ram_fsm[2:2]),.O(un74_addr));
defparam desc3158.INIT=16'h2220;
  LUT4 desc3159(.I0(write_ram_ptr[1:1]),.I1(write_ram_ptr[0:0]),.I2(write_ram_fsm[3:3]),.I3(write_ram_fsm[2:2]),.O(un106_addr));
defparam desc3159.INIT=16'h8880;
  LUT4 desc3160(.I0(write_ram_ptr[1:1]),.I1(write_ram_ptr[0:0]),.I2(write_ram_fsm[3:3]),.I3(write_ram_fsm[2:2]),.O(un42_addr));
defparam desc3160.INIT=16'h4440;
  LUT4 read_ram_fsm_1_2_sqmuxa_i_o3_lut6_2_o6(.I0(reorder_tvalid_fast[1:1]),.I1(read_ram_fsm_1_1_rep1),.I2(read_ram_fsm_1_0_rep1),.I3(traceback_tvalid[1:1]),.O(N_720));
defparam read_ram_fsm_1_2_sqmuxa_i_o3_lut6_2_o6.INIT=16'hEFCF;
  LUT2 read_ram_fsm_1_2_sqmuxa_i_o3_lut6_2_o5(.I0(read_ram_fsm_1_1_rep1),.I1(read_ram_fsm_1_0_rep1),.O(N_1733));
defparam read_ram_fsm_1_2_sqmuxa_i_o3_lut6_2_o5.INIT=4'hE;
  LUT4 desc3161(.I0(ram_tvalid[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep1),.I3(ram_buffer_full[1:1]),.O(un21_m_axis_output_tvalid_int));
defparam desc3161.INIT=16'h0080;
  LUT4 desc3162(.I0(ram_window_tuser[1:1]),.I1(ram_tvalid[1:1]),.I2(traceback_tvalid[1:1]),.I3(reorder_tvalid_1_rep1),.O(un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5));
defparam desc3162.INIT=16'hF888;
  LUT4 write_window_complete_RNIV26T_o6(.I0(write_window_complete),.I1(read_ram_fsm_1[0:0]),.I2(read_ram_fsm_1[1:1]),.I3(next_traceback),.O(write_window_complete_RNIV26T_O6));
defparam write_window_complete_RNIV26T_o6.INIT=16'hCECC;
  LUT3 write_window_complete_RNIV26T_o5(.I0(aresetn),.I1(write_window_complete),.I2(next_traceback),.O(N_941s));
defparam write_window_complete_RNIV26T_o5.INIT=8'h28;
  LUT2 desc3163(.I0(CO0_4),.I1(SUM1_4_0),.O(un2_write_ram_ptr_2_iv_1_RNIGNT55_O6));
defparam desc3163.INIT=4'h6;
  LUT2 desc3164(.I0(CO0_4),.I1(SUM1_4_0),.O(N_430_fast));
defparam desc3164.INIT=4'h6;
  LUT2 desc3165(.I0(CO0_3),.I1(SUM1_3_0),.O(un2_write_ram_ptr_3_iv_1_RNI880U2_O6));
defparam desc3165.INIT=4'h6;
  LUT2 desc3166(.I0(CO0_3),.I1(SUM1_3_0),.O(N_426_fast));
defparam desc3166.INIT=4'h6;
endmodule
module trellis_traceback_inj (ram_window_tuser,ram_tvalid,traceback_tvalid,traceback_tdata,buffer_cnt,ram_last_tuser,buffer_cnt_0,ram_buffer_full,ram_buffer_0,ram_buffer_0_2,traceback_last_tuser,traceback_tlast,ram_tlast,reorder_tvalid_0_rep1,reorder_tvalid_0_rep2,aclk,aresetn_i,N_129,last_window,aresetn,N_130,last_window_0,m_axis_output_tlast);
input ram_window_tuser ;
input ram_tvalid ;
output traceback_tvalid ;
output traceback_tdata ;
input [2:0] buffer_cnt ;
input ram_last_tuser ;
input [2:0] buffer_cnt_0 ;
input ram_buffer_full ;
input [63:0] ram_buffer_0 ;
input [63:0] ram_buffer_0_2 ;
output traceback_last_tuser ;
output traceback_tlast ;
input ram_tlast ;
input reorder_tvalid_0_rep1 ;
input reorder_tvalid_0_rep2 ;
input aclk ;
input aresetn_i ;
input N_129 ;
input last_window ;
input aresetn ;
input N_130 ;
input last_window_0 ;
output m_axis_output_tlast ;
wire reorder_tvalid_0_rep1 ;
wire reorder_tvalid_0_rep2 ;
wire aclk ;
wire aresetn_i ;
wire N_129 ;
wire last_window ;
wire aresetn ;
wire N_130 ;
wire last_window_0 ;
wire m_axis_output_tlast ;
wire current_node_3_7muxnet_0_0 ;
wire current_node_3_7muxnet_1_0 ;
wire [5:0] current_node ;
wire current_node_3_4 ;
wire current_node_3_5 ;
wire current_node_3_1 ;
wire current_node_3_2 ;
wire current_node_3_60muxnet_0_0 ;
wire current_node_3_60muxnet_1_0 ;
wire current_node_3_57 ;
wire current_node_3_58 ;
wire current_node_3_54 ;
wire current_node_3_55 ;
wire current_node_3_53muxnet_0_0 ;
wire current_node_3_53muxnet_1_0 ;
wire current_node_3_50 ;
wire current_node_3_51 ;
wire current_node_3_47 ;
wire current_node_3_48 ;
wire current_node_3_45muxnet_0_0 ;
wire current_node_3_45muxnet_1_0 ;
wire current_node_3_42 ;
wire current_node_3_43 ;
wire current_node_3_39 ;
wire current_node_3_40 ;
wire current_node_3_38muxnet_0_0 ;
wire current_node_3_38muxnet_1_0 ;
wire current_node_3_35 ;
wire current_node_3_36 ;
wire current_node_3_32 ;
wire current_node_3_33 ;
wire current_node_3_29muxnet_0_0 ;
wire current_node_3_29muxnet_1_0 ;
wire current_node_3_26 ;
wire current_node_3_27 ;
wire current_node_3_23 ;
wire current_node_3_24 ;
wire current_node_3_22muxnet_0_0 ;
wire current_node_3_22muxnet_1_0 ;
wire current_node_3_19 ;
wire current_node_3_20 ;
wire current_node_3_16 ;
wire current_node_3_17 ;
wire current_node_3_14muxnet_0_0 ;
wire current_node_3_14muxnet_1_0 ;
wire current_node_3_11 ;
wire current_node_3_12 ;
wire current_node_3_8 ;
wire current_node_3_9 ;
wire current_node_3 ;
wire VCC ;
wire N_89_i ;
wire m_axis_output_tvalid_int_RNIKUO21_O5 ;
wire m_axis_output_tdata ;
wire N_2396 ;
wire N_2449 ;
wire N_2442 ;
wire N_2434 ;
wire N_2427 ;
wire N_2418 ;
wire N_2411 ;
wire N_2403 ;
wire N_113 ;
wire m_axis_output_tvalid_int_RNITMA01 ;
wire N_2420 ;
wire N_2451 ;
wire GND ;
// instances
  FDR m_axis_output_tdata_Z(.Q(traceback_tdata),.D(m_axis_output_tdata),.C(aclk),.R(aresetn_i));
  MUXF8 desc3167(.I0(current_node_3_7muxnet_0_0),.I1(current_node_3_7muxnet_1_0),.S(current_node[3:3]),.O(N_2396));
  MUXF7 desc3168(.I0(current_node_3_4),.I1(current_node_3_5),.S(current_node[4:4]),.O(current_node_3_7muxnet_1_0));
  MUXF7 desc3169(.I0(current_node_3_1),.I1(current_node_3_2),.S(current_node[4:4]),.O(current_node_3_7muxnet_0_0));
  MUXF8 desc3170(.I0(current_node_3_60muxnet_0_0),.I1(current_node_3_60muxnet_1_0),.S(current_node[3:3]),.O(N_2449));
  MUXF7 desc3171(.I0(current_node_3_57),.I1(current_node_3_58),.S(current_node[4:4]),.O(current_node_3_60muxnet_1_0));
  MUXF7 desc3172(.I0(current_node_3_54),.I1(current_node_3_55),.S(current_node[4:4]),.O(current_node_3_60muxnet_0_0));
  MUXF8 desc3173(.I0(current_node_3_53muxnet_0_0),.I1(current_node_3_53muxnet_1_0),.S(current_node[3:3]),.O(N_2442));
  MUXF7 desc3174(.I0(current_node_3_50),.I1(current_node_3_51),.S(current_node[4:4]),.O(current_node_3_53muxnet_1_0));
  MUXF7 desc3175(.I0(current_node_3_47),.I1(current_node_3_48),.S(current_node[4:4]),.O(current_node_3_53muxnet_0_0));
  MUXF8 desc3176(.I0(current_node_3_45muxnet_0_0),.I1(current_node_3_45muxnet_1_0),.S(current_node[3:3]),.O(N_2434));
  MUXF7 desc3177(.I0(current_node_3_42),.I1(current_node_3_43),.S(current_node[4:4]),.O(current_node_3_45muxnet_1_0));
  MUXF7 desc3178(.I0(current_node_3_39),.I1(current_node_3_40),.S(current_node[4:4]),.O(current_node_3_45muxnet_0_0));
  MUXF8 desc3179(.I0(current_node_3_38muxnet_0_0),.I1(current_node_3_38muxnet_1_0),.S(current_node[3:3]),.O(N_2427));
  MUXF7 desc3180(.I0(current_node_3_35),.I1(current_node_3_36),.S(current_node[4:4]),.O(current_node_3_38muxnet_1_0));
  MUXF7 desc3181(.I0(current_node_3_32),.I1(current_node_3_33),.S(current_node[4:4]),.O(current_node_3_38muxnet_0_0));
  MUXF8 desc3182(.I0(current_node_3_29muxnet_0_0),.I1(current_node_3_29muxnet_1_0),.S(current_node[3:3]),.O(N_2418));
  MUXF7 desc3183(.I0(current_node_3_26),.I1(current_node_3_27),.S(current_node[4:4]),.O(current_node_3_29muxnet_1_0));
  MUXF7 desc3184(.I0(current_node_3_23),.I1(current_node_3_24),.S(current_node[4:4]),.O(current_node_3_29muxnet_0_0));
  MUXF8 desc3185(.I0(current_node_3_22muxnet_0_0),.I1(current_node_3_22muxnet_1_0),.S(current_node[3:3]),.O(N_2411));
  MUXF7 desc3186(.I0(current_node_3_19),.I1(current_node_3_20),.S(current_node[4:4]),.O(current_node_3_22muxnet_1_0));
  MUXF7 desc3187(.I0(current_node_3_16),.I1(current_node_3_17),.S(current_node[4:4]),.O(current_node_3_22muxnet_0_0));
  MUXF8 desc3188(.I0(current_node_3_14muxnet_0_0),.I1(current_node_3_14muxnet_1_0),.S(current_node[3:3]),.O(N_2403));
  MUXF7 desc3189(.I0(current_node_3_11),.I1(current_node_3_12),.S(current_node[4:4]),.O(current_node_3_14muxnet_1_0));
  MUXF7 desc3190(.I0(current_node_3_8),.I1(current_node_3_9),.S(current_node[4:4]),.O(current_node_3_14muxnet_0_0));
  LUT5 desc3191(.I0(N_129),.I1(buffer_cnt[0:0]),.I2(buffer_cnt[1:1]),.I3(buffer_cnt[2:2]),.I4(last_window),.O(N_113));
defparam desc3191.INIT=32'h20000000;
  LUT6_L m_axis_output_tdata_e(.I0(traceback_tdata),.I1(ram_window_tuser),.I2(ram_tvalid),.I3(traceback_tvalid),.I4(reorder_tvalid_0_rep1),.I5(current_node[5:5]),.LO(m_axis_output_tdata));
defparam m_axis_output_tdata_e.INIT=64'hAAEAEAEAAA2A2A2A;
  LUT5 m_axis_output_tvalid_int_RNITMA01_cZ(.I0(aresetn),.I1(ram_last_tuser),.I2(ram_tvalid),.I3(traceback_tvalid),.I4(reorder_tvalid_0_rep1),.O(m_axis_output_tvalid_int_RNITMA01));
defparam m_axis_output_tvalid_int_RNITMA01_cZ.INIT=32'h55D5D5D5;
  MUXF7 desc3192(.I0(N_2420),.I1(N_2451),.S(current_node[0:0]),.O(current_node_3));
  LUT6 desc3193(.I0(N_113),.I1(N_130),.I2(buffer_cnt_0[0:0]),.I3(buffer_cnt_0[1:1]),.I4(buffer_cnt_0[2:2]),.I5(last_window_0),.O(m_axis_output_tlast));
defparam desc3193.INIT=64'hAEAAAAAAAAAAAAAA;
  LUT6 desc3194(.I0(ram_buffer_0[10:10]),.I1(ram_buffer_0[42:42]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[10:10]),.I5(ram_buffer_0_2[42:42]),.O(current_node_3_19));
defparam desc3194.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3195(.I0(ram_buffer_0[18:18]),.I1(ram_buffer_0[50:50]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[18:18]),.I5(ram_buffer_0_2[50:50]),.O(current_node_3_17));
defparam desc3195.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3196(.I0(ram_buffer_0[2:2]),.I1(ram_buffer_0[34:34]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[2:2]),.I5(ram_buffer_0_2[34:34]),.O(current_node_3_16));
defparam desc3196.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3197(.I0(ram_buffer_0[28:28]),.I1(ram_buffer_0[60:60]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[28:28]),.I5(ram_buffer_0_2[60:60]),.O(current_node_3_12));
defparam desc3197.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3198(.I0(ram_buffer_0[12:12]),.I1(ram_buffer_0[44:44]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[12:12]),.I5(ram_buffer_0_2[44:44]),.O(current_node_3_11));
defparam desc3198.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3199(.I0(ram_buffer_0[20:20]),.I1(ram_buffer_0[52:52]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[20:20]),.I5(ram_buffer_0_2[52:52]),.O(current_node_3_9));
defparam desc3199.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3200(.I0(ram_buffer_0[4:4]),.I1(ram_buffer_0[36:36]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[4:4]),.I5(ram_buffer_0_2[36:36]),.O(current_node_3_8));
defparam desc3200.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3201(.I0(ram_buffer_0[17:17]),.I1(ram_buffer_0[49:49]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[17:17]),.I5(ram_buffer_0_2[49:49]),.O(current_node_3_33));
defparam desc3201.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3202(.I0(ram_buffer_0[1:1]),.I1(ram_buffer_0[33:33]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[1:1]),.I5(ram_buffer_0_2[33:33]),.O(current_node_3_32));
defparam desc3202.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3203(.I0(ram_buffer_0[30:30]),.I1(ram_buffer_0[62:62]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[30:30]),.I5(ram_buffer_0_2[62:62]),.O(current_node_3_27));
defparam desc3203.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3204(.I0(ram_buffer_0[14:14]),.I1(ram_buffer_0[46:46]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[14:14]),.I5(ram_buffer_0_2[46:46]),.O(current_node_3_26));
defparam desc3204.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3205(.I0(ram_buffer_0[22:22]),.I1(ram_buffer_0[54:54]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[22:22]),.I5(ram_buffer_0_2[54:54]),.O(current_node_3_24));
defparam desc3205.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3206(.I0(ram_buffer_0[6:6]),.I1(ram_buffer_0[38:38]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[6:6]),.I5(ram_buffer_0_2[38:38]),.O(current_node_3_23));
defparam desc3206.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3207(.I0(ram_buffer_0[26:26]),.I1(ram_buffer_0[58:58]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[26:26]),.I5(ram_buffer_0_2[58:58]),.O(current_node_3_20));
defparam desc3207.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3208(.I0(ram_buffer_0[3:3]),.I1(ram_buffer_0[35:35]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[3:3]),.I5(ram_buffer_0_2[35:35]),.O(current_node_3_47));
defparam desc3208.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3209(.I0(ram_buffer_0[29:29]),.I1(ram_buffer_0[61:61]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[29:29]),.I5(ram_buffer_0_2[61:61]),.O(current_node_3_43));
defparam desc3209.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3210(.I0(ram_buffer_0[13:13]),.I1(ram_buffer_0[45:45]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[13:13]),.I5(ram_buffer_0_2[45:45]),.O(current_node_3_42));
defparam desc3210.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3211(.I0(ram_buffer_0[21:21]),.I1(ram_buffer_0[53:53]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[21:21]),.I5(ram_buffer_0_2[53:53]),.O(current_node_3_40));
defparam desc3211.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3212(.I0(ram_buffer_0[5:5]),.I1(ram_buffer_0[37:37]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[5:5]),.I5(ram_buffer_0_2[37:37]),.O(current_node_3_39));
defparam desc3212.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3213(.I0(ram_buffer_0[25:25]),.I1(ram_buffer_0[57:57]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[25:25]),.I5(ram_buffer_0_2[57:57]),.O(current_node_3_36));
defparam desc3213.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3214(.I0(ram_buffer_0[9:9]),.I1(ram_buffer_0[41:41]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[9:9]),.I5(ram_buffer_0_2[41:41]),.O(current_node_3_35));
defparam desc3214.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3215(.I0(ram_buffer_0[31:31]),.I1(ram_buffer_0[63:63]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[31:31]),.I5(ram_buffer_0_2[63:63]),.O(current_node_3_58));
defparam desc3215.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3216(.I0(ram_buffer_0[15:15]),.I1(ram_buffer_0[47:47]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[15:15]),.I5(ram_buffer_0_2[47:47]),.O(current_node_3_57));
defparam desc3216.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3217(.I0(ram_buffer_0[23:23]),.I1(ram_buffer_0[55:55]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[23:23]),.I5(ram_buffer_0_2[55:55]),.O(current_node_3_55));
defparam desc3217.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3218(.I0(ram_buffer_0[7:7]),.I1(ram_buffer_0[39:39]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[7:7]),.I5(ram_buffer_0_2[39:39]),.O(current_node_3_54));
defparam desc3218.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3219(.I0(ram_buffer_0[27:27]),.I1(ram_buffer_0[59:59]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[27:27]),.I5(ram_buffer_0_2[59:59]),.O(current_node_3_51));
defparam desc3219.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3220(.I0(ram_buffer_0[11:11]),.I1(ram_buffer_0[43:43]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[11:11]),.I5(ram_buffer_0_2[43:43]),.O(current_node_3_50));
defparam desc3220.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3221(.I0(ram_buffer_0[19:19]),.I1(ram_buffer_0[51:51]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[19:19]),.I5(ram_buffer_0_2[51:51]),.O(current_node_3_48));
defparam desc3221.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3222(.I0(ram_buffer_0[24:24]),.I1(ram_buffer_0[56:56]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[24:24]),.I5(ram_buffer_0_2[56:56]),.O(current_node_3_5));
defparam desc3222.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3223(.I0(ram_buffer_0[8:8]),.I1(ram_buffer_0[40:40]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[8:8]),.I5(ram_buffer_0_2[40:40]),.O(current_node_3_4));
defparam desc3223.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3224(.I0(ram_buffer_0[16:16]),.I1(ram_buffer_0[48:48]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[16:16]),.I5(ram_buffer_0_2[48:48]),.O(current_node_3_2));
defparam desc3224.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3225(.I0(ram_buffer_0[0:0]),.I1(ram_buffer_0[32:32]),.I2(current_node[5:5]),.I3(ram_buffer_full),.I4(ram_buffer_0_2[0:0]),.I5(ram_buffer_0_2[32:32]),.O(current_node_3_1));
defparam desc3225.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3226(.I0(current_node[1:1]),.I1(current_node[2:2]),.I2(N_2427),.I3(N_2434),.I4(N_2442),.I5(N_2449),.O(N_2451));
defparam desc3226.INIT=64'hFEBADC9876325410;
  LUT6 desc3227(.I0(current_node[1:1]),.I1(current_node[2:2]),.I2(N_2396),.I3(N_2403),.I4(N_2411),.I5(N_2418),.O(N_2420));
defparam desc3227.INIT=64'hFEBADC9876325410;
  FDR m_axis_output_tvalid_int_Z(.Q(traceback_tvalid),.D(m_axis_output_tvalid_int_RNIKUO21_O5),.C(aclk),.R(aresetn_i));
  FDRE desc3228(.Q(current_node[5:5]),.D(current_node[4:4]),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE desc3229(.Q(current_node[4:4]),.D(current_node[3:3]),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE desc3230(.Q(current_node[3:3]),.D(current_node[2:2]),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE desc3231(.Q(current_node[2:2]),.D(current_node[1:1]),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE desc3232(.Q(current_node[1:1]),.D(current_node[0:0]),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE desc3233(.Q(current_node[0:0]),.D(current_node_3),.C(aclk),.R(m_axis_output_tvalid_int_RNITMA01),.CE(N_89_i));
  FDRE m_axis_output_last_tuser_Z(.Q(traceback_last_tuser),.D(ram_last_tuser),.C(aclk),.R(aresetn_i),.CE(N_89_i));
  FDRE m_axis_output_tlast_Z(.Q(traceback_tlast),.D(ram_tlast),.C(aclk),.R(aresetn_i),.CE(N_89_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 m_axis_output_tvalid_int_RNIKUO21_o6(.I0(ram_tvalid),.I1(traceback_tvalid),.I2(reorder_tvalid_0_rep1),.O(N_89_i));
defparam m_axis_output_tvalid_int_RNIKUO21_o6.INIT=8'h2A;
  LUT4 m_axis_output_tvalid_int_RNIKUO21_o5(.I0(ram_window_tuser),.I1(ram_tvalid),.I2(traceback_tvalid),.I3(reorder_tvalid_0_rep2),.O(m_axis_output_tvalid_int_RNIKUO21_O5));
defparam m_axis_output_tvalid_int_RNIKUO21_o5.INIT=16'hF888;
endmodule
module trellis_traceback_1_inj (traceback_last_tuser,ram_tvalid,traceback_tvalid,traceback_tdata,ram_last_tuser,ram_window_tuser,ram_buffer_full,ram_buffer_1,ram_buffer_1_1,traceback_tlast,ram_tlast,reorder_tvalid_1_rep1,N_104,send_output_rep1,aclk,aresetn_i,aresetn,un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5);
output [1:1] traceback_last_tuser ;
input [1:1] ram_tvalid ;
output [1:1] traceback_tvalid ;
output [1:1] traceback_tdata ;
input [1:1] ram_last_tuser ;
input [1:1] ram_window_tuser ;
input [1:1] ram_buffer_full ;
input [63:0] ram_buffer_1 ;
input [63:0] ram_buffer_1_1 ;
output [1:1] traceback_tlast ;
input [1:1] ram_tlast ;
input reorder_tvalid_1_rep1 ;
input N_104 ;
output send_output_rep1 ;
input aclk ;
input aresetn_i ;
input aresetn ;
input un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ;
wire reorder_tvalid_1_rep1 ;
wire N_104 ;
wire send_output_rep1 ;
wire aclk ;
wire aresetn_i ;
wire aresetn ;
wire un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ;
wire current_node_3_60muxnet_0_0 ;
wire current_node_3_60muxnet_1_0 ;
wire [5:0] current_node ;
wire current_node_3_57_0 ;
wire current_node_3_58_0 ;
wire current_node_3_54_0 ;
wire current_node_3_55_0 ;
wire current_node_3_53muxnet_0_0 ;
wire current_node_3_53muxnet_1_0 ;
wire current_node_3_50_0 ;
wire current_node_3_51_0 ;
wire current_node_3_47_0 ;
wire current_node_3_48_0 ;
wire current_node_3_45muxnet_0_0 ;
wire current_node_3_45muxnet_1_0 ;
wire current_node_3_42_0 ;
wire current_node_3_43_0 ;
wire current_node_3_39_0 ;
wire current_node_3_40_0 ;
wire current_node_3_38muxnet_0_0 ;
wire current_node_3_38muxnet_1_0 ;
wire current_node_3_35_0 ;
wire current_node_3_36_0 ;
wire current_node_3_32_0 ;
wire current_node_3_33_0 ;
wire current_node_3_29muxnet_0_0 ;
wire current_node_3_29muxnet_1_0 ;
wire current_node_3_26_0 ;
wire current_node_3_27_0 ;
wire current_node_3_23_0 ;
wire current_node_3_24_0 ;
wire current_node_3_7muxnet_0_0 ;
wire current_node_3_7muxnet_1_0 ;
wire current_node_3_4_0 ;
wire current_node_3_5_0 ;
wire current_node_3_1_0 ;
wire current_node_3_2_0 ;
wire current_node_3_22muxnet_0_0 ;
wire current_node_3_22muxnet_1_0 ;
wire current_node_3_19_0 ;
wire current_node_3_20_0 ;
wire current_node_3_16_0 ;
wire current_node_3_17_0 ;
wire current_node_3_14muxnet_0_0 ;
wire current_node_3_14muxnet_1_0 ;
wire current_node_3_11_0 ;
wire current_node_3_12_0 ;
wire current_node_3_8_0 ;
wire current_node_3_9_0 ;
wire current_node_3 ;
wire VCC ;
wire N_90_i ;
wire m_axis_output_tdata ;
wire N_2512 ;
wire N_2505 ;
wire N_2497 ;
wire N_2490 ;
wire N_2481 ;
wire N_2459 ;
wire N_2474 ;
wire N_2466 ;
wire N_2483 ;
wire N_2514 ;
wire m_axis_output_tvalid_int_RNI3R871 ;
wire GND ;
// instances
  FDR m_axis_output_tdata_Z(.Q(traceback_tdata[1:1]),.D(m_axis_output_tdata),.C(aclk),.R(aresetn_i));
  MUXF8 desc3234(.I0(current_node_3_60muxnet_0_0),.I1(current_node_3_60muxnet_1_0),.S(current_node[3:3]),.O(N_2512));
  MUXF7 desc3235(.I0(current_node_3_57_0),.I1(current_node_3_58_0),.S(current_node[4:4]),.O(current_node_3_60muxnet_1_0));
  MUXF7 desc3236(.I0(current_node_3_54_0),.I1(current_node_3_55_0),.S(current_node[4:4]),.O(current_node_3_60muxnet_0_0));
  MUXF8 desc3237(.I0(current_node_3_53muxnet_0_0),.I1(current_node_3_53muxnet_1_0),.S(current_node[3:3]),.O(N_2505));
  MUXF7 desc3238(.I0(current_node_3_50_0),.I1(current_node_3_51_0),.S(current_node[4:4]),.O(current_node_3_53muxnet_1_0));
  MUXF7 desc3239(.I0(current_node_3_47_0),.I1(current_node_3_48_0),.S(current_node[4:4]),.O(current_node_3_53muxnet_0_0));
  MUXF8 desc3240(.I0(current_node_3_45muxnet_0_0),.I1(current_node_3_45muxnet_1_0),.S(current_node[3:3]),.O(N_2497));
  MUXF7 desc3241(.I0(current_node_3_42_0),.I1(current_node_3_43_0),.S(current_node[4:4]),.O(current_node_3_45muxnet_1_0));
  MUXF7 desc3242(.I0(current_node_3_39_0),.I1(current_node_3_40_0),.S(current_node[4:4]),.O(current_node_3_45muxnet_0_0));
  MUXF8 desc3243(.I0(current_node_3_38muxnet_0_0),.I1(current_node_3_38muxnet_1_0),.S(current_node[3:3]),.O(N_2490));
  MUXF7 desc3244(.I0(current_node_3_35_0),.I1(current_node_3_36_0),.S(current_node[4:4]),.O(current_node_3_38muxnet_1_0));
  MUXF7 desc3245(.I0(current_node_3_32_0),.I1(current_node_3_33_0),.S(current_node[4:4]),.O(current_node_3_38muxnet_0_0));
  MUXF8 desc3246(.I0(current_node_3_29muxnet_0_0),.I1(current_node_3_29muxnet_1_0),.S(current_node[3:3]),.O(N_2481));
  MUXF7 desc3247(.I0(current_node_3_26_0),.I1(current_node_3_27_0),.S(current_node[4:4]),.O(current_node_3_29muxnet_1_0));
  MUXF7 desc3248(.I0(current_node_3_23_0),.I1(current_node_3_24_0),.S(current_node[4:4]),.O(current_node_3_29muxnet_0_0));
  MUXF8 desc3249(.I0(current_node_3_7muxnet_0_0),.I1(current_node_3_7muxnet_1_0),.S(current_node[3:3]),.O(N_2459));
  MUXF7 desc3250(.I0(current_node_3_4_0),.I1(current_node_3_5_0),.S(current_node[4:4]),.O(current_node_3_7muxnet_1_0));
  MUXF7 desc3251(.I0(current_node_3_1_0),.I1(current_node_3_2_0),.S(current_node[4:4]),.O(current_node_3_7muxnet_0_0));
  MUXF8 desc3252(.I0(current_node_3_22muxnet_0_0),.I1(current_node_3_22muxnet_1_0),.S(current_node[3:3]),.O(N_2474));
  MUXF7 desc3253(.I0(current_node_3_19_0),.I1(current_node_3_20_0),.S(current_node[4:4]),.O(current_node_3_22muxnet_1_0));
  MUXF7 desc3254(.I0(current_node_3_16_0),.I1(current_node_3_17_0),.S(current_node[4:4]),.O(current_node_3_22muxnet_0_0));
  MUXF8 desc3255(.I0(current_node_3_14muxnet_0_0),.I1(current_node_3_14muxnet_1_0),.S(current_node[3:3]),.O(N_2466));
  MUXF7 desc3256(.I0(current_node_3_11_0),.I1(current_node_3_12_0),.S(current_node[4:4]),.O(current_node_3_14muxnet_1_0));
  MUXF7 desc3257(.I0(current_node_3_8_0),.I1(current_node_3_9_0),.S(current_node[4:4]),.O(current_node_3_14muxnet_0_0));
  MUXF7 desc3258(.I0(N_2483),.I1(N_2514),.S(current_node[0:0]),.O(current_node_3));
  LUT5 m_axis_output_tvalid_int_RNI3R871_cZ(.I0(aresetn),.I1(ram_last_tuser[1:1]),.I2(ram_tvalid[1:1]),.I3(traceback_tvalid[1:1]),.I4(reorder_tvalid_1_rep1),.O(m_axis_output_tvalid_int_RNI3R871));
defparam m_axis_output_tvalid_int_RNI3R871_cZ.INIT=32'h55D5D5D5;
  LUT6_L m_axis_output_tdata_e(.I0(traceback_tdata[1:1]),.I1(ram_window_tuser[1:1]),.I2(ram_tvalid[1:1]),.I3(traceback_tvalid[1:1]),.I4(reorder_tvalid_1_rep1),.I5(current_node[5:5]),.LO(m_axis_output_tdata));
defparam m_axis_output_tdata_e.INIT=64'hAAEAEAEAAA2A2A2A;
  LUT6 desc3259(.I0(ram_buffer_1[1:1]),.I1(ram_buffer_1[33:33]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[1:1]),.I5(ram_buffer_1_1[33:33]),.O(current_node_3_32_0));
defparam desc3259.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3260(.I0(ram_buffer_1[4:4]),.I1(ram_buffer_1[36:36]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[4:4]),.I5(ram_buffer_1_1[36:36]),.O(current_node_3_8_0));
defparam desc3260.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3261(.I0(ram_buffer_1[10:10]),.I1(ram_buffer_1[42:42]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[10:10]),.I5(ram_buffer_1_1[42:42]),.O(current_node_3_19_0));
defparam desc3261.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3262(.I0(ram_buffer_1[18:18]),.I1(ram_buffer_1[50:50]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[18:18]),.I5(ram_buffer_1_1[50:50]),.O(current_node_3_17_0));
defparam desc3262.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3263(.I0(ram_buffer_1[2:2]),.I1(ram_buffer_1[34:34]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[2:2]),.I5(ram_buffer_1_1[34:34]),.O(current_node_3_16_0));
defparam desc3263.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3264(.I0(ram_buffer_1[28:28]),.I1(ram_buffer_1[60:60]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[28:28]),.I5(ram_buffer_1_1[60:60]),.O(current_node_3_12_0));
defparam desc3264.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3265(.I0(ram_buffer_1[12:12]),.I1(ram_buffer_1[44:44]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[12:12]),.I5(ram_buffer_1_1[44:44]),.O(current_node_3_11_0));
defparam desc3265.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3266(.I0(ram_buffer_1[20:20]),.I1(ram_buffer_1[52:52]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[20:20]),.I5(ram_buffer_1_1[52:52]),.O(current_node_3_9_0));
defparam desc3266.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3267(.I0(ram_buffer_1[17:17]),.I1(ram_buffer_1[49:49]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[17:17]),.I5(ram_buffer_1_1[49:49]),.O(current_node_3_33_0));
defparam desc3267.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3268(.I0(ram_buffer_1[30:30]),.I1(ram_buffer_1[62:62]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[30:30]),.I5(ram_buffer_1_1[62:62]),.O(current_node_3_27_0));
defparam desc3268.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3269(.I0(ram_buffer_1[14:14]),.I1(ram_buffer_1[46:46]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[14:14]),.I5(ram_buffer_1_1[46:46]),.O(current_node_3_26_0));
defparam desc3269.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3270(.I0(ram_buffer_1[22:22]),.I1(ram_buffer_1[54:54]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[22:22]),.I5(ram_buffer_1_1[54:54]),.O(current_node_3_24_0));
defparam desc3270.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3271(.I0(ram_buffer_1[6:6]),.I1(ram_buffer_1[38:38]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[6:6]),.I5(ram_buffer_1_1[38:38]),.O(current_node_3_23_0));
defparam desc3271.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3272(.I0(ram_buffer_1[26:26]),.I1(ram_buffer_1[58:58]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[26:26]),.I5(ram_buffer_1_1[58:58]),.O(current_node_3_20_0));
defparam desc3272.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3273(.I0(ram_buffer_1[3:3]),.I1(ram_buffer_1[35:35]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[3:3]),.I5(ram_buffer_1_1[35:35]),.O(current_node_3_47_0));
defparam desc3273.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3274(.I0(ram_buffer_1[29:29]),.I1(ram_buffer_1[61:61]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[29:29]),.I5(ram_buffer_1_1[61:61]),.O(current_node_3_43_0));
defparam desc3274.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3275(.I0(ram_buffer_1[13:13]),.I1(ram_buffer_1[45:45]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[13:13]),.I5(ram_buffer_1_1[45:45]),.O(current_node_3_42_0));
defparam desc3275.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3276(.I0(ram_buffer_1[21:21]),.I1(ram_buffer_1[53:53]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[21:21]),.I5(ram_buffer_1_1[53:53]),.O(current_node_3_40_0));
defparam desc3276.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3277(.I0(ram_buffer_1[5:5]),.I1(ram_buffer_1[37:37]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[5:5]),.I5(ram_buffer_1_1[37:37]),.O(current_node_3_39_0));
defparam desc3277.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3278(.I0(ram_buffer_1[25:25]),.I1(ram_buffer_1[57:57]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[25:25]),.I5(ram_buffer_1_1[57:57]),.O(current_node_3_36_0));
defparam desc3278.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3279(.I0(ram_buffer_1[9:9]),.I1(ram_buffer_1[41:41]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[9:9]),.I5(ram_buffer_1_1[41:41]),.O(current_node_3_35_0));
defparam desc3279.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3280(.I0(ram_buffer_1[31:31]),.I1(ram_buffer_1[63:63]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[31:31]),.I5(ram_buffer_1_1[63:63]),.O(current_node_3_58_0));
defparam desc3280.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3281(.I0(ram_buffer_1[15:15]),.I1(ram_buffer_1[47:47]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[15:15]),.I5(ram_buffer_1_1[47:47]),.O(current_node_3_57_0));
defparam desc3281.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3282(.I0(ram_buffer_1[23:23]),.I1(ram_buffer_1[55:55]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[23:23]),.I5(ram_buffer_1_1[55:55]),.O(current_node_3_55_0));
defparam desc3282.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3283(.I0(ram_buffer_1[7:7]),.I1(ram_buffer_1[39:39]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[7:7]),.I5(ram_buffer_1_1[39:39]),.O(current_node_3_54_0));
defparam desc3283.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3284(.I0(ram_buffer_1[27:27]),.I1(ram_buffer_1[59:59]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[27:27]),.I5(ram_buffer_1_1[59:59]),.O(current_node_3_51_0));
defparam desc3284.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3285(.I0(ram_buffer_1[11:11]),.I1(ram_buffer_1[43:43]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[11:11]),.I5(ram_buffer_1_1[43:43]),.O(current_node_3_50_0));
defparam desc3285.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3286(.I0(ram_buffer_1[19:19]),.I1(ram_buffer_1[51:51]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[19:19]),.I5(ram_buffer_1_1[51:51]),.O(current_node_3_48_0));
defparam desc3286.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3287(.I0(ram_buffer_1[24:24]),.I1(ram_buffer_1[56:56]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[24:24]),.I5(ram_buffer_1_1[56:56]),.O(current_node_3_5_0));
defparam desc3287.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3288(.I0(ram_buffer_1[8:8]),.I1(ram_buffer_1[40:40]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[8:8]),.I5(ram_buffer_1_1[40:40]),.O(current_node_3_4_0));
defparam desc3288.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3289(.I0(ram_buffer_1[16:16]),.I1(ram_buffer_1[48:48]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[16:16]),.I5(ram_buffer_1_1[48:48]),.O(current_node_3_2_0));
defparam desc3289.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3290(.I0(ram_buffer_1[0:0]),.I1(ram_buffer_1[32:32]),.I2(current_node[5:5]),.I3(ram_buffer_full[1:1]),.I4(ram_buffer_1_1[0:0]),.I5(ram_buffer_1_1[32:32]),.O(current_node_3_1_0));
defparam desc3290.INIT=64'hCAFFCAF0CA0FCA00;
  LUT6 desc3291(.I0(current_node[1:1]),.I1(current_node[2:2]),.I2(N_2490),.I3(N_2497),.I4(N_2505),.I5(N_2512),.O(N_2514));
defparam desc3291.INIT=64'hFEBADC9876325410;
  LUT6 desc3292(.I0(current_node[1:1]),.I1(current_node[2:2]),.I2(N_2459),.I3(N_2466),.I4(N_2474),.I5(N_2481),.O(N_2483));
defparam desc3292.INIT=64'hFEBADC9876325410;
  FDR m_axis_output_tvalid_int_Z(.Q(traceback_tvalid[1:1]),.D(un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5),.C(aclk),.R(aresetn_i));
  FDRE desc3293(.Q(current_node[5:5]),.D(current_node[4:4]),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE desc3294(.Q(current_node[4:4]),.D(current_node[3:3]),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE desc3295(.Q(current_node[3:3]),.D(current_node[2:2]),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE desc3296(.Q(current_node[2:2]),.D(current_node[1:1]),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE desc3297(.Q(current_node[1:1]),.D(current_node[0:0]),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE desc3298(.Q(current_node[0:0]),.D(current_node_3),.C(aclk),.R(m_axis_output_tvalid_int_RNI3R871),.CE(N_90_i));
  FDRE m_axis_output_last_tuser_Z(.Q(traceback_last_tuser[1:1]),.D(ram_last_tuser[1:1]),.C(aclk),.R(aresetn_i),.CE(N_90_i));
  FDRE m_axis_output_tlast_Z(.Q(traceback_tlast[1:1]),.D(ram_tlast[1:1]),.C(aclk),.R(aresetn_i),.CE(N_90_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 m_axis_output_last_tuser_RNIVMJF1_o6(.I0(ram_tvalid[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep1),.O(N_90_i));
defparam m_axis_output_last_tuser_RNIVMJF1_o6.INIT=8'h2A;
  LUT4 m_axis_output_last_tuser_RNIVMJF1_o5(.I0(traceback_last_tuser[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep1),.I3(N_104),.O(send_output_rep1));
defparam m_axis_output_last_tuser_RNIVMJF1_o5.INIT=16'h08F8;
endmodule
module reorder_inj (traceback_last_tuser,traceback_tvalid,reorder_tvalid_fast,reorder_tvalid_0,traceback_tlast,current_active,reorder_last_tuser,buffer_cnt_1,buffer_cnt_2,buffer_cnt_0,reorder_tdata_0,traceback_tdata,N_104,m_axis_output_tvalid,aresetn,reorder_tvalid_1_rep1,m_axis_output_tready,aclk,aresetn_i,last_window,send_output_rep1,m_axis_output_tdata,N_130);
input [1:1] traceback_last_tuser ;
input [1:1] traceback_tvalid ;
output [1:1] reorder_tvalid_fast ;
input reorder_tvalid_0 ;
input [1:1] traceback_tlast ;
input current_active ;
output [1:1] reorder_last_tuser ;
output buffer_cnt_1 ;
output buffer_cnt_2 ;
output buffer_cnt_0 ;
input reorder_tdata_0 ;
input [1:1] traceback_tdata ;
output N_104 ;
output m_axis_output_tvalid ;
input aresetn ;
output reorder_tvalid_1_rep1 ;
input m_axis_output_tready ;
input aclk ;
input aresetn_i ;
output last_window ;
input send_output_rep1 ;
output m_axis_output_tdata ;
output N_130 ;
wire reorder_tvalid_0 ;
wire buffer_cnt_1 ;
wire buffer_cnt_2 ;
wire buffer_cnt_0 ;
wire reorder_tdata_0 ;
wire N_104 ;
wire m_axis_output_tvalid ;
wire aresetn ;
wire reorder_tvalid_1_rep1 ;
wire m_axis_output_tready ;
wire aclk ;
wire aresetn_i ;
wire last_window ;
wire send_output_rep1 ;
wire m_axis_output_tdata ;
wire N_130 ;
wire [1:1] reorder_tvalid ;
wire [95:1] buffer_sreg ;
wire [95:0] buffer_sreg_7 ;
wire [1:1] reorder_tdata ;
wire [2:2] buffer_end ;
wire [1:1] buffer_end_0_0 ;
wire [6:3] buffer_cnt ;
wire reorder_tvalid_1_rep2 ;
wire VCC ;
wire send_output ;
wire send_output_rep2 ;
wire un1_buffer_cnt_1_axb_0 ;
wire un1_buffer_cnt_1_s_2 ;
wire GND ;
wire N_35_i ;
wire N_31_i ;
wire un1_buffer_cnt_1_s_1 ;
wire un1_buffer_cnt_1_s_3 ;
wire N_33_i ;
wire N_37_i ;
wire un1_buffer_cnt_1_s_4 ;
wire un1_buffer_cnt_1_s_6 ;
wire N_39_i ;
wire N_43_i ;
wire un1_buffer_cnt_1_s_5 ;
wire N_41_i ;
wire send_output_fast ;
wire un1_buffer_cnt_1_axb_1 ;
wire un1_buffer_cnt_1_axb_2 ;
wire un1_buffer_cnt_1_axb_3 ;
wire un1_buffer_cnt_1_axb_4 ;
wire un1_buffer_cnt_1_axb_5 ;
wire m_axis_output_last_tuser ;
wire last_window_0 ;
wire N_21 ;
wire un1_buffer_cnt_1_axb_6 ;
wire N_15_i ;
wire N_105 ;
wire un1_buffer_cnt_1_cry_5 ;
wire un1_buffer_cnt_1_cry_4 ;
wire un1_buffer_cnt_1_cry_3 ;
wire un1_buffer_cnt_1_cry_2 ;
wire un1_buffer_cnt_1_cry_1 ;
wire un1_buffer_cnt_1_cry_0 ;
// instances
  LUT6 desc3299(.I0(N_104),.I1(aresetn),.I2(buffer_end[2:2]),.I3(reorder_tvalid_1_rep1),.I4(traceback_tlast[1:1]),.I5(traceback_tvalid[1:1]),.O(buffer_end_0_0[1:1]));
defparam desc3299.INIT=64'h4044404040404040;
  LUT4 un1_buffer_cnt_1_axb_1_cZ(.I0(current_active),.I1(buffer_cnt_1),.I2(m_axis_output_tready),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_1));
defparam un1_buffer_cnt_1_axb_1_cZ.INIT=16'h6CCC;
  LUT4 un1_buffer_cnt_1_axb_2_cZ(.I0(current_active),.I1(buffer_cnt_2),.I2(m_axis_output_tready),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_2));
defparam un1_buffer_cnt_1_axb_2_cZ.INIT=16'h6CCC;
  LUT4 un1_buffer_cnt_1_axb_3_cZ(.I0(current_active),.I1(buffer_cnt[3:3]),.I2(m_axis_output_tready),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_3));
defparam un1_buffer_cnt_1_axb_3_cZ.INIT=16'h6CCC;
  LUT4 un1_buffer_cnt_1_axb_4_cZ(.I0(current_active),.I1(buffer_cnt[4:4]),.I2(m_axis_output_tready),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_4));
defparam un1_buffer_cnt_1_axb_4_cZ.INIT=16'h6CCC;
  LUT4 desc3300(.I0(current_active),.I1(buffer_cnt[5:5]),.I2(m_axis_output_tready),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_5));
defparam desc3300.INIT=16'h6CCC;
  FDR send_output_Z(.Q(reorder_tvalid[1:1]),.D(send_output),.C(aclk),.R(aresetn_i));
  FDR m_axis_output_last_tuser_Z(.Q(reorder_last_tuser[1:1]),.D(m_axis_output_last_tuser),.C(aclk),.R(aresetn_i));
  FDR last_window_Z(.Q(last_window),.D(last_window_0),.C(aclk),.R(aresetn_i));
  FDR send_output_fast_Z(.Q(reorder_tvalid_fast[1:1]),.D(send_output_fast),.C(aclk),.R(aresetn_i));
  FDR send_output_rep1_Z(.Q(reorder_tvalid_1_rep1),.D(send_output_rep1),.C(aclk),.R(aresetn_i));
  FDR send_output_rep2_Z(.Q(reorder_tvalid_1_rep2),.D(send_output_rep2),.C(aclk),.R(aresetn_i));
  LUT5_L last_window_e(.I0(last_window),.I1(traceback_tlast[1:1]),.I2(traceback_tvalid[1:1]),.I3(reorder_tvalid_1_rep1),.I4(N_104),.LO(last_window_0));
defparam last_window_e.INIT=32'h00C0AAEA;
  LUT4 buffer_sreg_1_sqmuxa_i_0(.I0(m_axis_output_tready),.I1(current_active),.I2(traceback_tvalid[1:1]),.I3(reorder_tvalid_1_rep1),.O(N_21));
defparam buffer_sreg_1_sqmuxa_i_0.INIT=16'h88F0;
  LUT4 un1_buffer_cnt_1_axb_6_cZ(.I0(m_axis_output_tready),.I1(buffer_cnt[6:6]),.I2(current_active),.I3(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_6));
defparam un1_buffer_cnt_1_axb_6_cZ.INIT=16'h6CCC;
  LUT6 un1_buffer_cnt_1_axb_0_cZ(.I0(m_axis_output_tready),.I1(traceback_last_tuser[1:1]),.I2(buffer_cnt_0),.I3(current_active),.I4(traceback_tvalid[1:1]),.I5(reorder_tvalid_1_rep1),.O(un1_buffer_cnt_1_axb_0));
defparam un1_buffer_cnt_1_axb_0_cZ.INIT=64'h5AF05AF0C3C3F0F0;
  LUT3 send_output_rep1_RNI47FT(.I0(m_axis_output_tready),.I1(current_active),.I2(reorder_tvalid_1_rep1),.O(N_15_i));
defparam send_output_rep1_RNI47FT.INIT=8'h80;
  FD desc3301(.Q(buffer_end[2:2]),.D(buffer_end_0_0[1:1]),.C(aclk));
  LUT3_L m_axis_output_last_tuser_e(.I0(reorder_last_tuser[1:1]),.I1(buffer_cnt_0),.I2(N_105),.LO(m_axis_output_last_tuser));
defparam m_axis_output_last_tuser_e.INIT=8'hCA;
  LUT3 m_axis_output_tdata_i_m2(.I0(current_active),.I1(reorder_tdata_0),.I2(reorder_tdata[1:1]),.O(m_axis_output_tdata));
defparam m_axis_output_tdata_i_m2.INIT=8'hE4;
  LUT3_L desc3302(.I0(buffer_sreg[1:1]),.I1(traceback_tdata[1:1]),.I2(reorder_tvalid_1_rep1),.LO(buffer_sreg_7[0:0]));
defparam desc3302.INIT=8'hAC;
  LUT4 desc3303(.I0(buffer_cnt[3:3]),.I1(buffer_cnt[4:4]),.I2(buffer_cnt[5:5]),.I3(buffer_cnt[6:6]),.O(N_130));
defparam desc3303.INIT=16'h0001;
  LUT6_L un1_m_axis_output_tready_1_i_a2(.I0(buffer_end[2:2]),.I1(buffer_cnt_1),.I2(buffer_cnt_2),.I3(buffer_cnt_0),.I4(N_130),.I5(N_15_i),.LO(N_105));
defparam un1_m_axis_output_tready_1_i_a2.INIT=64'h0381000000000000;
  LUT6 un1_rst_0_a2(.I0(buffer_end[2:2]),.I1(buffer_cnt_1),.I2(buffer_cnt_2),.I3(buffer_cnt_0),.I4(N_130),.I5(N_15_i),.O(N_104));
defparam un1_rst_0_a2.INIT=64'h0081000000000000;
  XORCY un1_buffer_cnt_1_s_6_cZ(.LI(un1_buffer_cnt_1_axb_6),.CI(un1_buffer_cnt_1_cry_5),.O(un1_buffer_cnt_1_s_6));
  XORCY un1_buffer_cnt_1_s_5_cZ(.LI(un1_buffer_cnt_1_axb_5),.CI(un1_buffer_cnt_1_cry_4),.O(un1_buffer_cnt_1_s_5));
  MUXCY_L un1_buffer_cnt_1_cry_5_cZ(.DI(N_15_i),.CI(un1_buffer_cnt_1_cry_4),.S(un1_buffer_cnt_1_axb_5),.LO(un1_buffer_cnt_1_cry_5));
  XORCY un1_buffer_cnt_1_s_4_cZ(.LI(un1_buffer_cnt_1_axb_4),.CI(un1_buffer_cnt_1_cry_3),.O(un1_buffer_cnt_1_s_4));
  MUXCY_L un1_buffer_cnt_1_cry_4_cZ(.DI(N_15_i),.CI(un1_buffer_cnt_1_cry_3),.S(un1_buffer_cnt_1_axb_4),.LO(un1_buffer_cnt_1_cry_4));
  XORCY un1_buffer_cnt_1_s_3_cZ(.LI(un1_buffer_cnt_1_axb_3),.CI(un1_buffer_cnt_1_cry_2),.O(un1_buffer_cnt_1_s_3));
  MUXCY_L un1_buffer_cnt_1_cry_3_cZ(.DI(N_15_i),.CI(un1_buffer_cnt_1_cry_2),.S(un1_buffer_cnt_1_axb_3),.LO(un1_buffer_cnt_1_cry_3));
  XORCY un1_buffer_cnt_1_s_2_cZ(.LI(un1_buffer_cnt_1_axb_2),.CI(un1_buffer_cnt_1_cry_1),.O(un1_buffer_cnt_1_s_2));
  MUXCY_L un1_buffer_cnt_1_cry_2_cZ(.DI(N_15_i),.CI(un1_buffer_cnt_1_cry_1),.S(un1_buffer_cnt_1_axb_2),.LO(un1_buffer_cnt_1_cry_2));
  XORCY un1_buffer_cnt_1_s_1_cZ(.LI(un1_buffer_cnt_1_axb_1),.CI(un1_buffer_cnt_1_cry_0),.O(un1_buffer_cnt_1_s_1));
  MUXCY_L un1_buffer_cnt_1_cry_1_cZ(.DI(N_15_i),.CI(un1_buffer_cnt_1_cry_0),.S(un1_buffer_cnt_1_axb_1),.LO(un1_buffer_cnt_1_cry_1));
  MUXCY_L un1_buffer_cnt_1_cry_0_cZ(.DI(buffer_cnt_0),.CI(GND),.S(un1_buffer_cnt_1_axb_0),.LO(un1_buffer_cnt_1_cry_0));
  FDRE desc3304(.Q(buffer_sreg[95:95]),.D(buffer_sreg_7[95:95]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3305(.Q(buffer_sreg[94:94]),.D(buffer_sreg_7[94:94]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3306(.Q(buffer_sreg[93:93]),.D(buffer_sreg_7[93:93]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3307(.Q(buffer_sreg[92:92]),.D(buffer_sreg_7[92:92]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3308(.Q(buffer_sreg[91:91]),.D(buffer_sreg_7[91:91]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3309(.Q(buffer_sreg[90:90]),.D(buffer_sreg_7[90:90]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3310(.Q(buffer_sreg[89:89]),.D(buffer_sreg_7[89:89]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3311(.Q(buffer_sreg[88:88]),.D(buffer_sreg_7[88:88]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3312(.Q(buffer_sreg[87:87]),.D(buffer_sreg_7[87:87]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3313(.Q(buffer_sreg[86:86]),.D(buffer_sreg_7[86:86]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3314(.Q(buffer_sreg[85:85]),.D(buffer_sreg_7[85:85]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3315(.Q(buffer_sreg[84:84]),.D(buffer_sreg_7[84:84]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3316(.Q(buffer_sreg[83:83]),.D(buffer_sreg_7[83:83]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3317(.Q(buffer_sreg[82:82]),.D(buffer_sreg_7[82:82]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3318(.Q(buffer_sreg[81:81]),.D(buffer_sreg_7[81:81]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3319(.Q(buffer_sreg[80:80]),.D(buffer_sreg_7[80:80]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3320(.Q(buffer_sreg[79:79]),.D(buffer_sreg_7[79:79]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3321(.Q(buffer_sreg[78:78]),.D(buffer_sreg_7[78:78]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3322(.Q(buffer_sreg[77:77]),.D(buffer_sreg_7[77:77]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3323(.Q(buffer_sreg[76:76]),.D(buffer_sreg_7[76:76]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3324(.Q(buffer_sreg[75:75]),.D(buffer_sreg_7[75:75]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3325(.Q(buffer_sreg[74:74]),.D(buffer_sreg_7[74:74]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3326(.Q(buffer_sreg[73:73]),.D(buffer_sreg_7[73:73]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3327(.Q(buffer_sreg[72:72]),.D(buffer_sreg_7[72:72]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3328(.Q(buffer_sreg[71:71]),.D(buffer_sreg_7[71:71]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3329(.Q(buffer_sreg[70:70]),.D(buffer_sreg_7[70:70]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3330(.Q(buffer_sreg[69:69]),.D(buffer_sreg_7[69:69]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3331(.Q(buffer_sreg[68:68]),.D(buffer_sreg_7[68:68]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3332(.Q(buffer_sreg[67:67]),.D(buffer_sreg_7[67:67]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3333(.Q(buffer_sreg[66:66]),.D(buffer_sreg_7[66:66]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3334(.Q(buffer_sreg[65:65]),.D(buffer_sreg_7[65:65]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3335(.Q(buffer_sreg[64:64]),.D(buffer_sreg_7[64:64]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3336(.Q(buffer_sreg[63:63]),.D(buffer_sreg_7[63:63]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3337(.Q(buffer_sreg[62:62]),.D(buffer_sreg_7[62:62]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3338(.Q(buffer_sreg[61:61]),.D(buffer_sreg_7[61:61]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3339(.Q(buffer_sreg[60:60]),.D(buffer_sreg_7[60:60]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3340(.Q(buffer_sreg[59:59]),.D(buffer_sreg_7[59:59]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3341(.Q(buffer_sreg[58:58]),.D(buffer_sreg_7[58:58]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3342(.Q(buffer_sreg[57:57]),.D(buffer_sreg_7[57:57]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3343(.Q(buffer_sreg[56:56]),.D(buffer_sreg_7[56:56]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3344(.Q(buffer_sreg[55:55]),.D(buffer_sreg_7[55:55]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3345(.Q(buffer_sreg[54:54]),.D(buffer_sreg_7[54:54]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3346(.Q(buffer_sreg[53:53]),.D(buffer_sreg_7[53:53]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3347(.Q(buffer_sreg[52:52]),.D(buffer_sreg_7[52:52]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3348(.Q(buffer_sreg[51:51]),.D(buffer_sreg_7[51:51]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3349(.Q(buffer_sreg[50:50]),.D(buffer_sreg_7[50:50]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3350(.Q(buffer_sreg[49:49]),.D(buffer_sreg_7[49:49]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3351(.Q(buffer_sreg[48:48]),.D(buffer_sreg_7[48:48]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3352(.Q(buffer_sreg[47:47]),.D(buffer_sreg_7[47:47]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3353(.Q(buffer_sreg[46:46]),.D(buffer_sreg_7[46:46]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3354(.Q(buffer_sreg[45:45]),.D(buffer_sreg_7[45:45]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3355(.Q(buffer_sreg[44:44]),.D(buffer_sreg_7[44:44]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3356(.Q(buffer_sreg[43:43]),.D(buffer_sreg_7[43:43]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3357(.Q(buffer_sreg[42:42]),.D(buffer_sreg_7[42:42]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3358(.Q(buffer_sreg[41:41]),.D(buffer_sreg_7[41:41]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3359(.Q(buffer_sreg[40:40]),.D(buffer_sreg_7[40:40]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3360(.Q(buffer_sreg[39:39]),.D(buffer_sreg_7[39:39]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3361(.Q(buffer_sreg[38:38]),.D(buffer_sreg_7[38:38]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3362(.Q(buffer_sreg[37:37]),.D(buffer_sreg_7[37:37]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3363(.Q(buffer_sreg[36:36]),.D(buffer_sreg_7[36:36]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3364(.Q(buffer_sreg[35:35]),.D(buffer_sreg_7[35:35]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3365(.Q(buffer_sreg[34:34]),.D(buffer_sreg_7[34:34]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3366(.Q(buffer_sreg[33:33]),.D(buffer_sreg_7[33:33]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3367(.Q(buffer_sreg[32:32]),.D(buffer_sreg_7[32:32]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3368(.Q(buffer_sreg[31:31]),.D(buffer_sreg_7[31:31]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3369(.Q(buffer_sreg[30:30]),.D(buffer_sreg_7[30:30]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3370(.Q(buffer_sreg[29:29]),.D(buffer_sreg_7[29:29]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3371(.Q(buffer_sreg[28:28]),.D(buffer_sreg_7[28:28]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3372(.Q(buffer_sreg[27:27]),.D(buffer_sreg_7[27:27]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3373(.Q(buffer_sreg[26:26]),.D(buffer_sreg_7[26:26]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3374(.Q(buffer_sreg[25:25]),.D(buffer_sreg_7[25:25]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3375(.Q(buffer_sreg[24:24]),.D(buffer_sreg_7[24:24]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3376(.Q(buffer_sreg[23:23]),.D(buffer_sreg_7[23:23]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3377(.Q(buffer_sreg[22:22]),.D(buffer_sreg_7[22:22]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3378(.Q(buffer_sreg[21:21]),.D(buffer_sreg_7[21:21]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3379(.Q(buffer_sreg[20:20]),.D(buffer_sreg_7[20:20]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3380(.Q(buffer_sreg[19:19]),.D(buffer_sreg_7[19:19]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3381(.Q(buffer_sreg[18:18]),.D(buffer_sreg_7[18:18]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3382(.Q(buffer_sreg[17:17]),.D(buffer_sreg_7[17:17]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3383(.Q(buffer_sreg[16:16]),.D(buffer_sreg_7[16:16]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3384(.Q(buffer_sreg[15:15]),.D(buffer_sreg_7[15:15]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3385(.Q(buffer_sreg[14:14]),.D(buffer_sreg_7[14:14]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3386(.Q(buffer_sreg[13:13]),.D(buffer_sreg_7[13:13]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3387(.Q(buffer_sreg[12:12]),.D(buffer_sreg_7[12:12]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3388(.Q(buffer_sreg[11:11]),.D(buffer_sreg_7[11:11]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3389(.Q(buffer_sreg[10:10]),.D(buffer_sreg_7[10:10]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3390(.Q(buffer_sreg[9:9]),.D(buffer_sreg_7[9:9]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3391(.Q(buffer_sreg[8:8]),.D(buffer_sreg_7[8:8]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3392(.Q(buffer_sreg[7:7]),.D(buffer_sreg_7[7:7]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3393(.Q(buffer_sreg[6:6]),.D(buffer_sreg_7[6:6]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3394(.Q(buffer_sreg[5:5]),.D(buffer_sreg_7[5:5]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3395(.Q(buffer_sreg[4:4]),.D(buffer_sreg_7[4:4]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3396(.Q(buffer_sreg[3:3]),.D(buffer_sreg_7[3:3]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3397(.Q(buffer_sreg[2:2]),.D(buffer_sreg_7[2:2]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3398(.Q(buffer_sreg[1:1]),.D(buffer_sreg_7[1:1]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDRE desc3399(.Q(reorder_tdata[1:1]),.D(buffer_sreg_7[0:0]),.C(aclk),.R(aresetn_i),.CE(N_21));
  FDR desc3400(.Q(buffer_cnt[6:6]),.D(N_43_i),.C(aclk),.R(aresetn_i));
  FDR desc3401(.Q(buffer_cnt[5:5]),.D(N_41_i),.C(aclk),.R(aresetn_i));
  FDR desc3402(.Q(buffer_cnt[4:4]),.D(N_39_i),.C(aclk),.R(aresetn_i));
  FDR desc3403(.Q(buffer_cnt[3:3]),.D(N_37_i),.C(aclk),.R(aresetn_i));
  FDR desc3404(.Q(buffer_cnt_2),.D(N_35_i),.C(aclk),.R(aresetn_i));
  FDR desc3405(.Q(buffer_cnt_1),.D(N_33_i),.C(aclk),.R(aresetn_i));
  FDR desc3406(.Q(buffer_cnt_0),.D(N_31_i),.C(aclk),.R(aresetn_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT2 desc3407(.I0(reorder_tvalid_0),.I1(reorder_tvalid[1:1]),.O(m_axis_output_tvalid));
defparam desc3407.INIT=4'hE;
  LUT3 desc3408(.I0(buffer_sreg[52:52]),.I1(buffer_sreg[54:54]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[53:53]));
defparam desc3408.INIT=8'hCA;
  LUT3 desc3409(.I0(buffer_sreg[43:43]),.I1(buffer_sreg[45:45]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[44:44]));
defparam desc3409.INIT=8'hCA;
  LUT3 desc3410(.I0(buffer_sreg[44:44]),.I1(buffer_sreg[46:46]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[45:45]));
defparam desc3410.INIT=8'hCA;
  LUT3 desc3411(.I0(buffer_sreg[41:41]),.I1(buffer_sreg[43:43]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[42:42]));
defparam desc3411.INIT=8'hCA;
  LUT3 desc3412(.I0(buffer_sreg[42:42]),.I1(buffer_sreg[44:44]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[43:43]));
defparam desc3412.INIT=8'hCA;
  LUT3 desc3413(.I0(buffer_sreg[38:38]),.I1(buffer_sreg[40:40]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[39:39]));
defparam desc3413.INIT=8'hCA;
  LUT3 desc3414(.I0(buffer_sreg[39:39]),.I1(buffer_sreg[41:41]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[40:40]));
defparam desc3414.INIT=8'hCA;
  LUT3 desc3415(.I0(buffer_sreg[35:35]),.I1(buffer_sreg[37:37]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[36:36]));
defparam desc3415.INIT=8'hCA;
  LUT3 desc3416(.I0(buffer_sreg[36:36]),.I1(buffer_sreg[38:38]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[37:37]));
defparam desc3416.INIT=8'hCA;
  LUT3 desc3417(.I0(buffer_sreg[33:33]),.I1(buffer_sreg[35:35]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[34:34]));
defparam desc3417.INIT=8'hCA;
  LUT3 desc3418(.I0(buffer_sreg[34:34]),.I1(buffer_sreg[36:36]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[35:35]));
defparam desc3418.INIT=8'hCA;
  LUT3 desc3419(.I0(buffer_sreg[31:31]),.I1(buffer_sreg[33:33]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[32:32]));
defparam desc3419.INIT=8'hCA;
  LUT3 desc3420(.I0(buffer_sreg[32:32]),.I1(buffer_sreg[34:34]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[33:33]));
defparam desc3420.INIT=8'hCA;
  LUT3 desc3421(.I0(buffer_sreg[29:29]),.I1(buffer_sreg[31:31]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[30:30]));
defparam desc3421.INIT=8'hCA;
  LUT3 desc3422(.I0(buffer_sreg[30:30]),.I1(buffer_sreg[32:32]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[31:31]));
defparam desc3422.INIT=8'hCA;
  LUT3 desc3423(.I0(buffer_sreg[27:27]),.I1(buffer_sreg[29:29]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[28:28]));
defparam desc3423.INIT=8'hCA;
  LUT3 desc3424(.I0(buffer_sreg[28:28]),.I1(buffer_sreg[30:30]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[29:29]));
defparam desc3424.INIT=8'hCA;
  LUT3 desc3425(.I0(buffer_sreg[25:25]),.I1(buffer_sreg[27:27]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[26:26]));
defparam desc3425.INIT=8'hCA;
  LUT3 desc3426(.I0(buffer_sreg[26:26]),.I1(buffer_sreg[28:28]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[27:27]));
defparam desc3426.INIT=8'hCA;
  LUT3 desc3427(.I0(buffer_sreg[23:23]),.I1(buffer_sreg[25:25]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[24:24]));
defparam desc3427.INIT=8'hCA;
  LUT3 desc3428(.I0(buffer_sreg[24:24]),.I1(buffer_sreg[26:26]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[25:25]));
defparam desc3428.INIT=8'hCA;
  LUT3 desc3429(.I0(buffer_sreg[21:21]),.I1(buffer_sreg[23:23]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[22:22]));
defparam desc3429.INIT=8'hCA;
  LUT3 desc3430(.I0(buffer_sreg[22:22]),.I1(buffer_sreg[24:24]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[23:23]));
defparam desc3430.INIT=8'hCA;
  LUT3 desc3431(.I0(buffer_sreg[19:19]),.I1(buffer_sreg[21:21]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[20:20]));
defparam desc3431.INIT=8'hCA;
  LUT3 desc3432(.I0(buffer_sreg[20:20]),.I1(buffer_sreg[22:22]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[21:21]));
defparam desc3432.INIT=8'hCA;
  LUT3 desc3433(.I0(buffer_sreg[17:17]),.I1(buffer_sreg[19:19]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[18:18]));
defparam desc3433.INIT=8'hCA;
  LUT3 desc3434(.I0(buffer_sreg[18:18]),.I1(buffer_sreg[20:20]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[19:19]));
defparam desc3434.INIT=8'hCA;
  LUT3 desc3435(.I0(buffer_sreg[15:15]),.I1(buffer_sreg[17:17]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[16:16]));
defparam desc3435.INIT=8'hCA;
  LUT3 desc3436(.I0(buffer_sreg[16:16]),.I1(buffer_sreg[18:18]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[17:17]));
defparam desc3436.INIT=8'hCA;
  LUT3 desc3437(.I0(buffer_sreg[13:13]),.I1(buffer_sreg[15:15]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[14:14]));
defparam desc3437.INIT=8'hCA;
  LUT3 desc3438(.I0(buffer_sreg[14:14]),.I1(buffer_sreg[16:16]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[15:15]));
defparam desc3438.INIT=8'hCA;
  LUT3 desc3439(.I0(buffer_sreg[10:10]),.I1(buffer_sreg[12:12]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[11:11]));
defparam desc3439.INIT=8'hCA;
  LUT3 desc3440(.I0(buffer_sreg[11:11]),.I1(buffer_sreg[13:13]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[12:12]));
defparam desc3440.INIT=8'hCA;
  LUT3 desc3441(.I0(buffer_sreg[9:9]),.I1(buffer_sreg[11:11]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[10:10]));
defparam desc3441.INIT=8'hCA;
  LUT3 desc3442(.I0(buffer_sreg[37:37]),.I1(buffer_sreg[39:39]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[38:38]));
defparam desc3442.INIT=8'hCA;
  LUT3 desc3443(.I0(buffer_sreg[7:7]),.I1(buffer_sreg[9:9]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[8:8]));
defparam desc3443.INIT=8'hCA;
  LUT3 desc3444(.I0(buffer_sreg[8:8]),.I1(buffer_sreg[10:10]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[9:9]));
defparam desc3444.INIT=8'hCA;
  LUT3 desc3445(.I0(buffer_sreg[5:5]),.I1(buffer_sreg[7:7]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[6:6]));
defparam desc3445.INIT=8'hCA;
  LUT3 desc3446(.I0(buffer_sreg[6:6]),.I1(buffer_sreg[8:8]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[7:7]));
defparam desc3446.INIT=8'hCA;
  LUT3 desc3447(.I0(buffer_sreg[4:4]),.I1(buffer_sreg[6:6]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[5:5]));
defparam desc3447.INIT=8'hCA;
  LUT3 desc3448(.I0(buffer_sreg[40:40]),.I1(buffer_sreg[42:42]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[41:41]));
defparam desc3448.INIT=8'hCA;
  LUT3 desc3449(.I0(buffer_sreg[2:2]),.I1(buffer_sreg[4:4]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[3:3]));
defparam desc3449.INIT=8'hCA;
  LUT3 desc3450(.I0(buffer_sreg[3:3]),.I1(buffer_sreg[5:5]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[4:4]));
defparam desc3450.INIT=8'hCA;
  LUT3 desc3451(.I0(buffer_sreg[2:2]),.I1(reorder_tdata[1:1]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[1:1]));
defparam desc3451.INIT=8'hAC;
  LUT3 desc3452(.I0(buffer_sreg[1:1]),.I1(buffer_sreg[3:3]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[2:2]));
defparam desc3452.INIT=8'hCA;
  LUT3 desc3453(.I0(buffer_sreg[95:95]),.I1(buffer_sreg[93:93]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[94:94]));
defparam desc3453.INIT=8'hAC;
  LUT2 desc3454(.I0(buffer_sreg[94:94]),.I1(reorder_tvalid[1:1]),.O(buffer_sreg_7[95:95]));
defparam desc3454.INIT=4'h2;
  LUT3 desc3455(.I0(buffer_sreg[91:91]),.I1(buffer_sreg[93:93]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[92:92]));
defparam desc3455.INIT=8'hCA;
  LUT3 desc3456(.I0(buffer_sreg[92:92]),.I1(buffer_sreg[94:94]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[93:93]));
defparam desc3456.INIT=8'hCA;
  LUT3 desc3457(.I0(buffer_sreg[89:89]),.I1(buffer_sreg[91:91]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[90:90]));
defparam desc3457.INIT=8'hCA;
  LUT3 desc3458(.I0(buffer_sreg[90:90]),.I1(buffer_sreg[92:92]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[91:91]));
defparam desc3458.INIT=8'hCA;
  LUT3 desc3459(.I0(buffer_sreg[87:87]),.I1(buffer_sreg[89:89]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[88:88]));
defparam desc3459.INIT=8'hCA;
  LUT3 desc3460(.I0(buffer_sreg[88:88]),.I1(buffer_sreg[90:90]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[89:89]));
defparam desc3460.INIT=8'hCA;
  LUT3 desc3461(.I0(buffer_sreg[85:85]),.I1(buffer_sreg[87:87]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[86:86]));
defparam desc3461.INIT=8'hCA;
  LUT3 desc3462(.I0(buffer_sreg[86:86]),.I1(buffer_sreg[88:88]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[87:87]));
defparam desc3462.INIT=8'hCA;
  LUT3 desc3463(.I0(buffer_sreg[83:83]),.I1(buffer_sreg[85:85]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[84:84]));
defparam desc3463.INIT=8'hCA;
  LUT3 desc3464(.I0(buffer_sreg[84:84]),.I1(buffer_sreg[86:86]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[85:85]));
defparam desc3464.INIT=8'hCA;
  LUT3 desc3465(.I0(buffer_sreg[81:81]),.I1(buffer_sreg[83:83]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[82:82]));
defparam desc3465.INIT=8'hCA;
  LUT3 desc3466(.I0(buffer_sreg[82:82]),.I1(buffer_sreg[84:84]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[83:83]));
defparam desc3466.INIT=8'hCA;
  LUT3 desc3467(.I0(buffer_sreg[79:79]),.I1(buffer_sreg[81:81]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[80:80]));
defparam desc3467.INIT=8'hCA;
  LUT3 desc3468(.I0(buffer_sreg[80:80]),.I1(buffer_sreg[82:82]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[81:81]));
defparam desc3468.INIT=8'hCA;
  LUT3 desc3469(.I0(buffer_sreg[77:77]),.I1(buffer_sreg[79:79]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[78:78]));
defparam desc3469.INIT=8'hCA;
  LUT3 desc3470(.I0(buffer_sreg[78:78]),.I1(buffer_sreg[80:80]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[79:79]));
defparam desc3470.INIT=8'hCA;
  LUT3 desc3471(.I0(buffer_sreg[75:75]),.I1(buffer_sreg[77:77]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[76:76]));
defparam desc3471.INIT=8'hCA;
  LUT3 desc3472(.I0(buffer_sreg[76:76]),.I1(buffer_sreg[78:78]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[77:77]));
defparam desc3472.INIT=8'hCA;
  LUT3 desc3473(.I0(buffer_sreg[73:73]),.I1(buffer_sreg[75:75]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[74:74]));
defparam desc3473.INIT=8'hCA;
  LUT3 desc3474(.I0(buffer_sreg[74:74]),.I1(buffer_sreg[76:76]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[75:75]));
defparam desc3474.INIT=8'hCA;
  LUT3 desc3475(.I0(buffer_sreg[71:71]),.I1(buffer_sreg[73:73]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[72:72]));
defparam desc3475.INIT=8'hCA;
  LUT3 desc3476(.I0(buffer_sreg[72:72]),.I1(buffer_sreg[74:74]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[73:73]));
defparam desc3476.INIT=8'hCA;
  LUT3 desc3477(.I0(buffer_sreg[69:69]),.I1(buffer_sreg[71:71]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[70:70]));
defparam desc3477.INIT=8'hCA;
  LUT3 desc3478(.I0(buffer_sreg[70:70]),.I1(buffer_sreg[72:72]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[71:71]));
defparam desc3478.INIT=8'hCA;
  LUT3 desc3479(.I0(buffer_sreg[67:67]),.I1(buffer_sreg[69:69]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[68:68]));
defparam desc3479.INIT=8'hCA;
  LUT3 desc3480(.I0(buffer_sreg[68:68]),.I1(buffer_sreg[70:70]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[69:69]));
defparam desc3480.INIT=8'hCA;
  LUT3 desc3481(.I0(buffer_sreg[65:65]),.I1(buffer_sreg[67:67]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[66:66]));
defparam desc3481.INIT=8'hCA;
  LUT3 desc3482(.I0(buffer_sreg[66:66]),.I1(buffer_sreg[68:68]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[67:67]));
defparam desc3482.INIT=8'hCA;
  LUT3 desc3483(.I0(buffer_sreg[63:63]),.I1(buffer_sreg[65:65]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[64:64]));
defparam desc3483.INIT=8'hCA;
  LUT3 desc3484(.I0(buffer_sreg[64:64]),.I1(buffer_sreg[66:66]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[65:65]));
defparam desc3484.INIT=8'hCA;
  LUT3 desc3485(.I0(buffer_sreg[61:61]),.I1(buffer_sreg[63:63]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[62:62]));
defparam desc3485.INIT=8'hCA;
  LUT3 desc3486(.I0(buffer_sreg[62:62]),.I1(buffer_sreg[64:64]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[63:63]));
defparam desc3486.INIT=8'hCA;
  LUT3 desc3487(.I0(buffer_sreg[59:59]),.I1(buffer_sreg[61:61]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[60:60]));
defparam desc3487.INIT=8'hCA;
  LUT3 desc3488(.I0(buffer_sreg[60:60]),.I1(buffer_sreg[62:62]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[61:61]));
defparam desc3488.INIT=8'hCA;
  LUT3 desc3489(.I0(buffer_sreg[57:57]),.I1(buffer_sreg[59:59]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[58:58]));
defparam desc3489.INIT=8'hCA;
  LUT3 desc3490(.I0(buffer_sreg[58:58]),.I1(buffer_sreg[60:60]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[59:59]));
defparam desc3490.INIT=8'hCA;
  LUT3 desc3491(.I0(buffer_sreg[55:55]),.I1(buffer_sreg[57:57]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[56:56]));
defparam desc3491.INIT=8'hCA;
  LUT3 desc3492(.I0(buffer_sreg[56:56]),.I1(buffer_sreg[58:58]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[57:57]));
defparam desc3492.INIT=8'hCA;
  LUT3 desc3493(.I0(buffer_sreg[53:53]),.I1(buffer_sreg[55:55]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[54:54]));
defparam desc3493.INIT=8'hCA;
  LUT3 desc3494(.I0(buffer_sreg[54:54]),.I1(buffer_sreg[56:56]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[55:55]));
defparam desc3494.INIT=8'hCA;
  LUT3 desc3495(.I0(buffer_sreg[51:51]),.I1(buffer_sreg[53:53]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[52:52]));
defparam desc3495.INIT=8'hCA;
  LUT3 desc3496(.I0(buffer_sreg[50:50]),.I1(buffer_sreg[52:52]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[51:51]));
defparam desc3496.INIT=8'hCA;
  LUT3 desc3497(.I0(buffer_sreg[49:49]),.I1(buffer_sreg[51:51]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[50:50]));
defparam desc3497.INIT=8'hCA;
  LUT3 desc3498(.I0(buffer_sreg[48:48]),.I1(buffer_sreg[50:50]),.I2(reorder_tvalid[1:1]),.O(buffer_sreg_7[49:49]));
defparam desc3498.INIT=8'hCA;
  LUT3 desc3499(.I0(buffer_sreg[47:47]),.I1(buffer_sreg[49:49]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[48:48]));
defparam desc3499.INIT=8'hCA;
  LUT3 desc3500(.I0(buffer_sreg[12:12]),.I1(buffer_sreg[14:14]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[13:13]));
defparam desc3500.INIT=8'hCA;
  LUT3 desc3501(.I0(buffer_sreg[45:45]),.I1(buffer_sreg[47:47]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[46:46]));
defparam desc3501.INIT=8'hCA;
  LUT3 desc3502(.I0(buffer_sreg[46:46]),.I1(buffer_sreg[48:48]),.I2(reorder_tvalid_1_rep2),.O(buffer_sreg_7[47:47]));
defparam desc3502.INIT=8'hCA;
  LUT2 un1_buffer_cnt_1_s_5_RNIVESF1_o6(.I0(N_104),.I1(un1_buffer_cnt_1_s_5),.O(N_41_i));
defparam un1_buffer_cnt_1_s_5_RNIVESF1_o6.INIT=4'h4;
  LUT4 un1_buffer_cnt_1_s_5_RNIVESF1_o5(.I0(traceback_last_tuser[1:1]),.I1(reorder_tvalid_fast[1:1]),.I2(traceback_tvalid[1:1]),.I3(N_104),.O(send_output_fast));
defparam un1_buffer_cnt_1_s_5_RNIVESF1_o5.INIT=16'h20EC;
  LUT2 un1_buffer_cnt_1_s_4_RNINDMT_o6(.I0(N_104),.I1(un1_buffer_cnt_1_s_4),.O(N_39_i));
defparam un1_buffer_cnt_1_s_4_RNINDMT_o6.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_4_RNINDMT_o5(.I0(N_104),.I1(un1_buffer_cnt_1_s_6),.O(N_43_i));
defparam un1_buffer_cnt_1_s_4_RNINDMT_o5.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_1_RNIHDMT_o6(.I0(N_104),.I1(un1_buffer_cnt_1_s_1),.O(N_33_i));
defparam un1_buffer_cnt_1_s_1_RNIHDMT_o6.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_1_RNIHDMT_o5(.I0(N_104),.I1(un1_buffer_cnt_1_s_3),.O(N_37_i));
defparam un1_buffer_cnt_1_s_1_RNIHDMT_o5.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_2_RNIN5341_o6(.I0(N_104),.I1(un1_buffer_cnt_1_s_2),.O(N_35_i));
defparam un1_buffer_cnt_1_s_2_RNIN5341_o6.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_2_RNIN5341_o5(.I0(un1_buffer_cnt_1_axb_0),.I1(N_104),.O(N_31_i));
defparam un1_buffer_cnt_1_s_2_RNIN5341_o5.INIT=4'h2;
  LUT4 send_output_e_lut6_2_o6(.I0(traceback_last_tuser[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid[1:1]),.I3(N_104),.O(send_output));
defparam send_output_e_lut6_2_o6.INIT=16'h08F8;
  LUT4 send_output_e_lut6_2_o5(.I0(traceback_last_tuser[1:1]),.I1(traceback_tvalid[1:1]),.I2(reorder_tvalid_1_rep2),.I3(N_104),.O(send_output_rep2));
defparam send_output_e_lut6_2_o5.INIT=16'h08F8;
endmodule
module reorder_1_inj (traceback_last_tuser,traceback_tvalid,reorder_tvalid_fast,reorder_tvalid,reorder_tdata,current_active,traceback_tlast,reorder_last_tuser,buffer_cnt_1,buffer_cnt_2,buffer_cnt_0,traceback_tdata,reorder_tvalid_0_rep1,reorder_tvalid_0_rep2,m_axis_output_tready,N_99,aresetn,aclk,aresetn_i,last_window,N_129);
input traceback_last_tuser ;
input traceback_tvalid ;
output reorder_tvalid_fast ;
output reorder_tvalid ;
output reorder_tdata ;
input current_active ;
input traceback_tlast ;
output reorder_last_tuser ;
output buffer_cnt_1 ;
output buffer_cnt_2 ;
output buffer_cnt_0 ;
input traceback_tdata ;
output reorder_tvalid_0_rep1 ;
output reorder_tvalid_0_rep2 ;
input m_axis_output_tready ;
output N_99 ;
input aresetn ;
input aclk ;
input aresetn_i ;
output last_window ;
output N_129 ;
wire buffer_cnt_1 ;
wire buffer_cnt_2 ;
wire buffer_cnt_0 ;
wire reorder_tvalid_0_rep1 ;
wire reorder_tvalid_0_rep2 ;
wire m_axis_output_tready ;
wire N_99 ;
wire aresetn ;
wire aclk ;
wire aresetn_i ;
wire last_window ;
wire N_129 ;
wire [95:1] buffer_sreg ;
wire [95:95] buffer_sreg_7 ;
wire [2:2] buffer_end ;
wire [1:1] buffer_end_0_0 ;
wire [6:3] buffer_cnt ;
wire un1_buffer_cnt_1_axb_0 ;
wire N_357 ;
wire un1_buffer_cnt_1_s_2_0 ;
wire GND ;
wire VCC ;
wire N_63_i ;
wire N_59_i ;
wire un1_buffer_cnt_1_s_1_0 ;
wire un1_buffer_cnt_1_s_3_0 ;
wire N_61_i ;
wire N_65_i ;
wire un1_buffer_cnt_1_s_4_0 ;
wire N_67_i ;
wire send_output_rep1 ;
wire un1_buffer_cnt_1_s_5_0 ;
wire N_69_i ;
wire send_output_fast ;
wire un1_buffer_cnt_1_s_6_0 ;
wire N_71_i ;
wire send_output_rep2 ;
wire N_252 ;
wire N_331 ;
wire N_253 ;
wire N_328 ;
wire N_254 ;
wire N_329 ;
wire N_255 ;
wire N_330 ;
wire N_256 ;
wire N_332 ;
wire N_257 ;
wire N_333 ;
wire N_258 ;
wire N_334 ;
wire N_259 ;
wire N_335 ;
wire N_260 ;
wire N_336 ;
wire N_262 ;
wire N_337 ;
wire N_263 ;
wire N_338 ;
wire N_264 ;
wire N_339 ;
wire N_265 ;
wire N_341 ;
wire N_266 ;
wire N_270 ;
wire N_267 ;
wire N_342 ;
wire N_268 ;
wire N_343 ;
wire N_269 ;
wire N_345 ;
wire N_271 ;
wire N_346 ;
wire N_273 ;
wire N_274 ;
wire N_275 ;
wire N_276 ;
wire N_277 ;
wire N_303 ;
wire N_278 ;
wire N_279 ;
wire N_280 ;
wire N_314 ;
wire N_281 ;
wire N_282 ;
wire N_283 ;
wire N_284 ;
wire N_285 ;
wire N_286 ;
wire N_287 ;
wire N_288 ;
wire N_289 ;
wire N_290 ;
wire N_291 ;
wire N_292 ;
wire N_293 ;
wire N_294 ;
wire N_295 ;
wire N_296 ;
wire N_297 ;
wire N_298 ;
wire N_299 ;
wire N_300 ;
wire N_301 ;
wire N_302 ;
wire N_304 ;
wire N_305 ;
wire N_306 ;
wire N_307 ;
wire N_308 ;
wire N_309 ;
wire N_310 ;
wire N_311 ;
wire N_312 ;
wire N_313 ;
wire N_315 ;
wire N_316 ;
wire N_317 ;
wire N_318 ;
wire N_319 ;
wire N_320 ;
wire N_321 ;
wire N_340 ;
wire N_322 ;
wire N_323 ;
wire N_324 ;
wire N_325 ;
wire N_326 ;
wire N_327 ;
wire N_344 ;
wire N_49 ;
wire un1_buffer_cnt_1_axb_1 ;
wire un1_buffer_cnt_1_axb_2 ;
wire un1_buffer_cnt_1_axb_3 ;
wire un1_buffer_cnt_1_axb_4 ;
wire un1_buffer_cnt_1_axb_5 ;
wire send_output ;
wire m_axis_output_last_tuser ;
wire last_window_0 ;
wire N_79 ;
wire m_axis_output_tready_0 ;
wire N_272 ;
wire N_261 ;
wire un1_buffer_cnt_1_axb_6 ;
wire un1_buffer_cnt_1_cry_5 ;
wire un1_buffer_cnt_1_cry_4 ;
wire un1_buffer_cnt_1_cry_3 ;
wire un1_buffer_cnt_1_cry_2 ;
wire un1_buffer_cnt_1_cry_1 ;
wire un1_buffer_cnt_1_cry_0 ;
// instances
  LUT6 desc3503(.I0(N_357),.I1(aresetn),.I2(buffer_end[2:2]),.I3(reorder_tvalid_0_rep1),.I4(traceback_tlast),.I5(traceback_tvalid),.O(buffer_end_0_0[1:1]));
defparam desc3503.INIT=64'h4044404040404040;
  LUT4 un1_buffer_cnt_1_axb_1_cZ(.I0(current_active),.I1(buffer_cnt_1),.I2(m_axis_output_tready),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_1));
defparam un1_buffer_cnt_1_axb_1_cZ.INIT=16'h9CCC;
  LUT4 un1_buffer_cnt_1_axb_2_cZ(.I0(current_active),.I1(buffer_cnt_2),.I2(m_axis_output_tready),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_2));
defparam un1_buffer_cnt_1_axb_2_cZ.INIT=16'h9CCC;
  LUT4 un1_buffer_cnt_1_axb_3_cZ(.I0(current_active),.I1(buffer_cnt[3:3]),.I2(m_axis_output_tready),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_3));
defparam un1_buffer_cnt_1_axb_3_cZ.INIT=16'h9CCC;
  LUT4 un1_buffer_cnt_1_axb_4_cZ(.I0(current_active),.I1(buffer_cnt[4:4]),.I2(m_axis_output_tready),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_4));
defparam un1_buffer_cnt_1_axb_4_cZ.INIT=16'h9CCC;
  LUT4 desc3504(.I0(current_active),.I1(buffer_cnt[5:5]),.I2(m_axis_output_tready),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_5));
defparam desc3504.INIT=16'h9CCC;
  FDR send_output_Z(.Q(reorder_tvalid),.D(send_output),.C(aclk),.R(aresetn_i));
  FDR m_axis_output_last_tuser_Z(.Q(reorder_last_tuser),.D(m_axis_output_last_tuser),.C(aclk),.R(aresetn_i));
  FDR last_window_Z(.Q(last_window),.D(last_window_0),.C(aclk),.R(aresetn_i));
  FDR send_output_fast_Z(.Q(reorder_tvalid_fast),.D(send_output_fast),.C(aclk),.R(aresetn_i));
  FDR send_output_rep1_Z(.Q(reorder_tvalid_0_rep1),.D(send_output_rep1),.C(aclk),.R(aresetn_i));
  FDR send_output_rep2_Z(.Q(reorder_tvalid_0_rep2),.D(send_output_rep2),.C(aclk),.R(aresetn_i));
  LUT5_L last_window_e(.I0(last_window),.I1(traceback_tlast),.I2(traceback_tvalid),.I3(reorder_tvalid_0_rep1),.I4(N_357),.LO(last_window_0));
defparam last_window_e.INIT=32'h00C0AAEA;
  LUT6 un1_buffer_cnt_1_axb_0_cZ(.I0(m_axis_output_tready),.I1(traceback_last_tuser),.I2(buffer_cnt_0),.I3(current_active),.I4(traceback_tvalid),.I5(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_0));
defparam un1_buffer_cnt_1_axb_0_cZ.INIT=64'hF05AF05AC3C3F0F0;
  LUT4 un1_m_axis_output_tready_1_i_o2(.I0(buffer_end[2:2]),.I1(buffer_cnt_1),.I2(buffer_cnt_2),.I3(buffer_cnt_0),.O(N_79));
defparam un1_m_axis_output_tready_1_i_o2.INIT=16'h0381;
  FD desc3505(.Q(buffer_end[2:2]),.D(buffer_end_0_0[1:1]),.C(aclk));
  LUT5_L m_axis_output_last_tuser_e(.I0(reorder_last_tuser),.I1(buffer_cnt_0),.I2(N_79),.I3(N_129),.I4(m_axis_output_tready_0),.LO(m_axis_output_last_tuser));
defparam m_axis_output_last_tuser_e.INIT=32'hCAAAAAAA;
  LUT3_L desc3506(.I0(buffer_sreg[1:1]),.I1(traceback_tdata),.I2(reorder_tvalid_0_rep2),.LO(N_272));
defparam desc3506.INIT=8'hAC;
  LUT3_L desc3507(.I0(buffer_sreg[73:73]),.I1(buffer_sreg[75:75]),.I2(reorder_tvalid),.LO(N_261));
defparam desc3507.INIT=8'hCA;
  LUT4 desc3508(.I0(buffer_cnt[3:3]),.I1(buffer_cnt[4:4]),.I2(buffer_cnt[5:5]),.I3(buffer_cnt[6:6]),.O(N_129));
defparam desc3508.INIT=16'h0001;
  LUT4 un1_buffer_cnt_1_axb_6_cZ(.I0(m_axis_output_tready),.I1(buffer_cnt[6:6]),.I2(current_active),.I3(reorder_tvalid_0_rep1),.O(un1_buffer_cnt_1_axb_6));
defparam un1_buffer_cnt_1_axb_6_cZ.INIT=16'hC6CC;
  LUT6 un1_rst_0_0_a2(.I0(buffer_end[2:2]),.I1(buffer_cnt_1),.I2(buffer_cnt_2),.I3(buffer_cnt_0),.I4(N_129),.I5(m_axis_output_tready_0),.O(N_357));
defparam un1_rst_0_0_a2.INIT=64'h0081000000000000;
  LUT4_L send_output_e(.I0(traceback_last_tuser),.I1(traceback_tvalid),.I2(reorder_tvalid),.I3(N_357),.LO(send_output));
defparam send_output_e.INIT=16'h08F8;
  LUT3 send_output_rep1_RNI39RJ(.I0(m_axis_output_tready),.I1(current_active),.I2(reorder_tvalid_0_rep1),.O(m_axis_output_tready_0));
defparam send_output_rep1_RNI39RJ.INIT=8'h20;
  XORCY un1_buffer_cnt_1_s_6(.LI(un1_buffer_cnt_1_axb_6),.CI(un1_buffer_cnt_1_cry_5),.O(un1_buffer_cnt_1_s_6_0));
  XORCY un1_buffer_cnt_1_s_5(.LI(un1_buffer_cnt_1_axb_5),.CI(un1_buffer_cnt_1_cry_4),.O(un1_buffer_cnt_1_s_5_0));
  MUXCY_L un1_buffer_cnt_1_cry_5_cZ(.DI(m_axis_output_tready_0),.CI(un1_buffer_cnt_1_cry_4),.S(un1_buffer_cnt_1_axb_5),.LO(un1_buffer_cnt_1_cry_5));
  XORCY un1_buffer_cnt_1_s_4(.LI(un1_buffer_cnt_1_axb_4),.CI(un1_buffer_cnt_1_cry_3),.O(un1_buffer_cnt_1_s_4_0));
  MUXCY_L un1_buffer_cnt_1_cry_4_cZ(.DI(m_axis_output_tready_0),.CI(un1_buffer_cnt_1_cry_3),.S(un1_buffer_cnt_1_axb_4),.LO(un1_buffer_cnt_1_cry_4));
  XORCY un1_buffer_cnt_1_s_3(.LI(un1_buffer_cnt_1_axb_3),.CI(un1_buffer_cnt_1_cry_2),.O(un1_buffer_cnt_1_s_3_0));
  MUXCY_L un1_buffer_cnt_1_cry_3_cZ(.DI(m_axis_output_tready_0),.CI(un1_buffer_cnt_1_cry_2),.S(un1_buffer_cnt_1_axb_3),.LO(un1_buffer_cnt_1_cry_3));
  XORCY un1_buffer_cnt_1_s_2(.LI(un1_buffer_cnt_1_axb_2),.CI(un1_buffer_cnt_1_cry_1),.O(un1_buffer_cnt_1_s_2_0));
  MUXCY_L un1_buffer_cnt_1_cry_2_cZ(.DI(m_axis_output_tready_0),.CI(un1_buffer_cnt_1_cry_1),.S(un1_buffer_cnt_1_axb_2),.LO(un1_buffer_cnt_1_cry_2));
  XORCY un1_buffer_cnt_1_s_1(.LI(un1_buffer_cnt_1_axb_1),.CI(un1_buffer_cnt_1_cry_0),.O(un1_buffer_cnt_1_s_1_0));
  MUXCY_L un1_buffer_cnt_1_cry_1_cZ(.DI(m_axis_output_tready_0),.CI(un1_buffer_cnt_1_cry_0),.S(un1_buffer_cnt_1_axb_1),.LO(un1_buffer_cnt_1_cry_1));
  MUXCY_L un1_buffer_cnt_1_cry_0_cZ(.DI(buffer_cnt_0),.CI(GND),.S(un1_buffer_cnt_1_axb_0),.LO(un1_buffer_cnt_1_cry_0));
  FDRE desc3509(.Q(buffer_sreg[95:95]),.D(buffer_sreg_7[95:95]),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3510(.Q(buffer_sreg[94:94]),.D(N_271),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3511(.Q(buffer_sreg[93:93]),.D(N_346),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3512(.Q(buffer_sreg[92:92]),.D(N_270),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3513(.Q(buffer_sreg[91:91]),.D(N_345),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3514(.Q(buffer_sreg[90:90]),.D(N_269),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3515(.Q(buffer_sreg[89:89]),.D(N_344),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3516(.Q(buffer_sreg[88:88]),.D(N_268),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3517(.Q(buffer_sreg[87:87]),.D(N_343),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3518(.Q(buffer_sreg[86:86]),.D(N_267),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3519(.Q(buffer_sreg[85:85]),.D(N_342),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3520(.Q(buffer_sreg[84:84]),.D(N_266),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3521(.Q(buffer_sreg[83:83]),.D(N_341),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3522(.Q(buffer_sreg[82:82]),.D(N_265),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3523(.Q(buffer_sreg[81:81]),.D(N_340),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3524(.Q(buffer_sreg[80:80]),.D(N_264),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3525(.Q(buffer_sreg[79:79]),.D(N_339),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3526(.Q(buffer_sreg[78:78]),.D(N_263),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3527(.Q(buffer_sreg[77:77]),.D(N_338),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3528(.Q(buffer_sreg[76:76]),.D(N_262),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3529(.Q(buffer_sreg[75:75]),.D(N_337),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3530(.Q(buffer_sreg[74:74]),.D(N_261),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3531(.Q(buffer_sreg[73:73]),.D(N_336),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3532(.Q(buffer_sreg[72:72]),.D(N_260),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3533(.Q(buffer_sreg[71:71]),.D(N_335),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3534(.Q(buffer_sreg[70:70]),.D(N_259),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3535(.Q(buffer_sreg[69:69]),.D(N_334),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3536(.Q(buffer_sreg[68:68]),.D(N_258),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3537(.Q(buffer_sreg[67:67]),.D(N_333),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3538(.Q(buffer_sreg[66:66]),.D(N_257),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3539(.Q(buffer_sreg[65:65]),.D(N_332),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3540(.Q(buffer_sreg[64:64]),.D(N_256),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3541(.Q(buffer_sreg[63:63]),.D(N_331),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3542(.Q(buffer_sreg[62:62]),.D(N_255),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3543(.Q(buffer_sreg[61:61]),.D(N_330),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3544(.Q(buffer_sreg[60:60]),.D(N_254),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3545(.Q(buffer_sreg[59:59]),.D(N_329),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3546(.Q(buffer_sreg[58:58]),.D(N_253),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3547(.Q(buffer_sreg[57:57]),.D(N_328),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3548(.Q(buffer_sreg[56:56]),.D(N_252),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3549(.Q(buffer_sreg[55:55]),.D(N_327),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3550(.Q(buffer_sreg[54:54]),.D(N_326),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3551(.Q(buffer_sreg[53:53]),.D(N_325),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3552(.Q(buffer_sreg[52:52]),.D(N_324),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3553(.Q(buffer_sreg[51:51]),.D(N_323),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3554(.Q(buffer_sreg[50:50]),.D(N_322),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3555(.Q(buffer_sreg[49:49]),.D(N_321),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3556(.Q(buffer_sreg[48:48]),.D(N_320),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3557(.Q(buffer_sreg[47:47]),.D(N_319),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3558(.Q(buffer_sreg[46:46]),.D(N_318),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3559(.Q(buffer_sreg[45:45]),.D(N_317),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3560(.Q(buffer_sreg[44:44]),.D(N_316),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3561(.Q(buffer_sreg[43:43]),.D(N_315),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3562(.Q(buffer_sreg[42:42]),.D(N_314),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3563(.Q(buffer_sreg[41:41]),.D(N_313),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3564(.Q(buffer_sreg[40:40]),.D(N_312),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3565(.Q(buffer_sreg[39:39]),.D(N_311),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3566(.Q(buffer_sreg[38:38]),.D(N_310),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3567(.Q(buffer_sreg[37:37]),.D(N_309),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3568(.Q(buffer_sreg[36:36]),.D(N_308),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3569(.Q(buffer_sreg[35:35]),.D(N_307),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3570(.Q(buffer_sreg[34:34]),.D(N_306),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3571(.Q(buffer_sreg[33:33]),.D(N_305),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3572(.Q(buffer_sreg[32:32]),.D(N_304),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3573(.Q(buffer_sreg[31:31]),.D(N_303),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3574(.Q(buffer_sreg[30:30]),.D(N_302),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3575(.Q(buffer_sreg[29:29]),.D(N_301),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3576(.Q(buffer_sreg[28:28]),.D(N_300),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3577(.Q(buffer_sreg[27:27]),.D(N_299),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3578(.Q(buffer_sreg[26:26]),.D(N_298),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3579(.Q(buffer_sreg[25:25]),.D(N_297),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3580(.Q(buffer_sreg[24:24]),.D(N_296),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3581(.Q(buffer_sreg[23:23]),.D(N_295),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3582(.Q(buffer_sreg[22:22]),.D(N_294),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3583(.Q(buffer_sreg[21:21]),.D(N_293),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3584(.Q(buffer_sreg[20:20]),.D(N_292),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3585(.Q(buffer_sreg[19:19]),.D(N_291),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3586(.Q(buffer_sreg[18:18]),.D(N_290),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3587(.Q(buffer_sreg[17:17]),.D(N_289),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3588(.Q(buffer_sreg[16:16]),.D(N_288),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3589(.Q(buffer_sreg[15:15]),.D(N_287),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3590(.Q(buffer_sreg[14:14]),.D(N_286),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3591(.Q(buffer_sreg[13:13]),.D(N_285),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3592(.Q(buffer_sreg[12:12]),.D(N_284),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3593(.Q(buffer_sreg[11:11]),.D(N_283),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3594(.Q(buffer_sreg[10:10]),.D(N_282),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3595(.Q(buffer_sreg[9:9]),.D(N_281),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3596(.Q(buffer_sreg[8:8]),.D(N_280),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3597(.Q(buffer_sreg[7:7]),.D(N_279),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3598(.Q(buffer_sreg[6:6]),.D(N_278),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3599(.Q(buffer_sreg[5:5]),.D(N_277),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3600(.Q(buffer_sreg[4:4]),.D(N_276),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3601(.Q(buffer_sreg[3:3]),.D(N_275),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3602(.Q(buffer_sreg[2:2]),.D(N_274),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3603(.Q(buffer_sreg[1:1]),.D(N_273),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDRE desc3604(.Q(reorder_tdata),.D(N_272),.C(aclk),.R(aresetn_i),.CE(N_49));
  FDR desc3605(.Q(buffer_cnt[6:6]),.D(N_71_i),.C(aclk),.R(aresetn_i));
  FDR desc3606(.Q(buffer_cnt[5:5]),.D(N_69_i),.C(aclk),.R(aresetn_i));
  FDR desc3607(.Q(buffer_cnt[4:4]),.D(N_67_i),.C(aclk),.R(aresetn_i));
  FDR desc3608(.Q(buffer_cnt[3:3]),.D(N_65_i),.C(aclk),.R(aresetn_i));
  FDR desc3609(.Q(buffer_cnt_2),.D(N_63_i),.C(aclk),.R(aresetn_i));
  FDR desc3610(.Q(buffer_cnt_1),.D(N_61_i),.C(aclk),.R(aresetn_i));
  FDR desc3611(.Q(buffer_cnt_0),.D(N_59_i),.C(aclk),.R(aresetn_i));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT2 send_output_fast_RNI41TV_o6(.I0(reorder_tvalid_fast),.I1(traceback_tvalid),.O(N_99));
defparam send_output_fast_RNI41TV_o6.INIT=4'h8;
  LUT4 send_output_fast_RNI41TV_o5(.I0(m_axis_output_tready),.I1(traceback_tvalid),.I2(current_active),.I3(reorder_tvalid_0_rep1),.O(N_49));
defparam send_output_fast_RNI41TV_o5.INIT=16'h0ACC;
  LUT3 desc3612(.I0(buffer_sreg[88:88]),.I1(buffer_sreg[90:90]),.I2(reorder_tvalid),.O(N_344));
defparam desc3612.INIT=8'hCA;
  LUT2 desc3613(.I0(buffer_sreg[94:94]),.I1(reorder_tvalid),.O(buffer_sreg_7[95:95]));
defparam desc3613.INIT=4'h2;
  LUT3 desc3614(.I0(buffer_sreg[53:53]),.I1(buffer_sreg[55:55]),.I2(reorder_tvalid),.O(N_326));
defparam desc3614.INIT=8'hCA;
  LUT3 desc3615(.I0(buffer_sreg[54:54]),.I1(buffer_sreg[56:56]),.I2(reorder_tvalid),.O(N_327));
defparam desc3615.INIT=8'hCA;
  LUT3 desc3616(.I0(buffer_sreg[51:51]),.I1(buffer_sreg[53:53]),.I2(reorder_tvalid),.O(N_324));
defparam desc3616.INIT=8'hCA;
  LUT3 desc3617(.I0(buffer_sreg[52:52]),.I1(buffer_sreg[54:54]),.I2(reorder_tvalid),.O(N_325));
defparam desc3617.INIT=8'hCA;
  LUT3 desc3618(.I0(buffer_sreg[49:49]),.I1(buffer_sreg[51:51]),.I2(reorder_tvalid),.O(N_322));
defparam desc3618.INIT=8'hCA;
  LUT3 desc3619(.I0(buffer_sreg[50:50]),.I1(buffer_sreg[52:52]),.I2(reorder_tvalid),.O(N_323));
defparam desc3619.INIT=8'hCA;
  LUT3 desc3620(.I0(buffer_sreg[48:48]),.I1(buffer_sreg[50:50]),.I2(reorder_tvalid),.O(N_321));
defparam desc3620.INIT=8'hCA;
  LUT3 desc3621(.I0(buffer_sreg[80:80]),.I1(buffer_sreg[82:82]),.I2(reorder_tvalid),.O(N_340));
defparam desc3621.INIT=8'hCA;
  LUT3 desc3622(.I0(buffer_sreg[46:46]),.I1(buffer_sreg[48:48]),.I2(reorder_tvalid),.O(N_319));
defparam desc3622.INIT=8'hCA;
  LUT3 desc3623(.I0(buffer_sreg[47:47]),.I1(buffer_sreg[49:49]),.I2(reorder_tvalid),.O(N_320));
defparam desc3623.INIT=8'hCA;
  LUT3 desc3624(.I0(buffer_sreg[44:44]),.I1(buffer_sreg[46:46]),.I2(reorder_tvalid_0_rep2),.O(N_317));
defparam desc3624.INIT=8'hCA;
  LUT3 desc3625(.I0(buffer_sreg[45:45]),.I1(buffer_sreg[47:47]),.I2(reorder_tvalid_0_rep2),.O(N_318));
defparam desc3625.INIT=8'hCA;
  LUT3 desc3626(.I0(buffer_sreg[42:42]),.I1(buffer_sreg[44:44]),.I2(reorder_tvalid_0_rep2),.O(N_315));
defparam desc3626.INIT=8'hCA;
  LUT3 desc3627(.I0(buffer_sreg[43:43]),.I1(buffer_sreg[45:45]),.I2(reorder_tvalid_0_rep2),.O(N_316));
defparam desc3627.INIT=8'hCA;
  LUT3 desc3628(.I0(buffer_sreg[39:39]),.I1(buffer_sreg[41:41]),.I2(reorder_tvalid_0_rep2),.O(N_312));
defparam desc3628.INIT=8'hCA;
  LUT3 desc3629(.I0(buffer_sreg[40:40]),.I1(buffer_sreg[42:42]),.I2(reorder_tvalid_0_rep2),.O(N_313));
defparam desc3629.INIT=8'hCA;
  LUT3 desc3630(.I0(buffer_sreg[37:37]),.I1(buffer_sreg[39:39]),.I2(reorder_tvalid_0_rep2),.O(N_310));
defparam desc3630.INIT=8'hCA;
  LUT3 desc3631(.I0(buffer_sreg[38:38]),.I1(buffer_sreg[40:40]),.I2(reorder_tvalid_0_rep2),.O(N_311));
defparam desc3631.INIT=8'hCA;
  LUT3 desc3632(.I0(buffer_sreg[35:35]),.I1(buffer_sreg[37:37]),.I2(reorder_tvalid_0_rep2),.O(N_308));
defparam desc3632.INIT=8'hCA;
  LUT3 desc3633(.I0(buffer_sreg[36:36]),.I1(buffer_sreg[38:38]),.I2(reorder_tvalid_0_rep2),.O(N_309));
defparam desc3633.INIT=8'hCA;
  LUT3 desc3634(.I0(buffer_sreg[33:33]),.I1(buffer_sreg[35:35]),.I2(reorder_tvalid_0_rep2),.O(N_306));
defparam desc3634.INIT=8'hCA;
  LUT3 desc3635(.I0(buffer_sreg[34:34]),.I1(buffer_sreg[36:36]),.I2(reorder_tvalid_0_rep2),.O(N_307));
defparam desc3635.INIT=8'hCA;
  LUT3 desc3636(.I0(buffer_sreg[31:31]),.I1(buffer_sreg[33:33]),.I2(reorder_tvalid_0_rep2),.O(N_304));
defparam desc3636.INIT=8'hCA;
  LUT3 desc3637(.I0(buffer_sreg[32:32]),.I1(buffer_sreg[34:34]),.I2(reorder_tvalid_0_rep2),.O(N_305));
defparam desc3637.INIT=8'hCA;
  LUT3 desc3638(.I0(buffer_sreg[28:28]),.I1(buffer_sreg[30:30]),.I2(reorder_tvalid_0_rep2),.O(N_301));
defparam desc3638.INIT=8'hCA;
  LUT3 desc3639(.I0(buffer_sreg[29:29]),.I1(buffer_sreg[31:31]),.I2(reorder_tvalid_0_rep2),.O(N_302));
defparam desc3639.INIT=8'hCA;
  LUT3 desc3640(.I0(buffer_sreg[26:26]),.I1(buffer_sreg[28:28]),.I2(reorder_tvalid_0_rep2),.O(N_299));
defparam desc3640.INIT=8'hCA;
  LUT3 desc3641(.I0(buffer_sreg[27:27]),.I1(buffer_sreg[29:29]),.I2(reorder_tvalid_0_rep2),.O(N_300));
defparam desc3641.INIT=8'hCA;
  LUT3 desc3642(.I0(buffer_sreg[24:24]),.I1(buffer_sreg[26:26]),.I2(reorder_tvalid_0_rep2),.O(N_297));
defparam desc3642.INIT=8'hCA;
  LUT3 desc3643(.I0(buffer_sreg[25:25]),.I1(buffer_sreg[27:27]),.I2(reorder_tvalid_0_rep2),.O(N_298));
defparam desc3643.INIT=8'hCA;
  LUT3 desc3644(.I0(buffer_sreg[22:22]),.I1(buffer_sreg[24:24]),.I2(reorder_tvalid_0_rep2),.O(N_295));
defparam desc3644.INIT=8'hCA;
  LUT3 desc3645(.I0(buffer_sreg[23:23]),.I1(buffer_sreg[25:25]),.I2(reorder_tvalid_0_rep2),.O(N_296));
defparam desc3645.INIT=8'hCA;
  LUT3 desc3646(.I0(buffer_sreg[20:20]),.I1(buffer_sreg[22:22]),.I2(reorder_tvalid_0_rep2),.O(N_293));
defparam desc3646.INIT=8'hCA;
  LUT3 desc3647(.I0(buffer_sreg[21:21]),.I1(buffer_sreg[23:23]),.I2(reorder_tvalid_0_rep2),.O(N_294));
defparam desc3647.INIT=8'hCA;
  LUT3 desc3648(.I0(buffer_sreg[18:18]),.I1(buffer_sreg[20:20]),.I2(reorder_tvalid_0_rep2),.O(N_291));
defparam desc3648.INIT=8'hCA;
  LUT3 desc3649(.I0(buffer_sreg[19:19]),.I1(buffer_sreg[21:21]),.I2(reorder_tvalid_0_rep2),.O(N_292));
defparam desc3649.INIT=8'hCA;
  LUT3 desc3650(.I0(buffer_sreg[16:16]),.I1(buffer_sreg[18:18]),.I2(reorder_tvalid_0_rep2),.O(N_289));
defparam desc3650.INIT=8'hCA;
  LUT3 desc3651(.I0(buffer_sreg[17:17]),.I1(buffer_sreg[19:19]),.I2(reorder_tvalid_0_rep2),.O(N_290));
defparam desc3651.INIT=8'hCA;
  LUT3 desc3652(.I0(buffer_sreg[14:14]),.I1(buffer_sreg[16:16]),.I2(reorder_tvalid_0_rep2),.O(N_287));
defparam desc3652.INIT=8'hCA;
  LUT3 desc3653(.I0(buffer_sreg[15:15]),.I1(buffer_sreg[17:17]),.I2(reorder_tvalid_0_rep2),.O(N_288));
defparam desc3653.INIT=8'hCA;
  LUT3 desc3654(.I0(buffer_sreg[12:12]),.I1(buffer_sreg[14:14]),.I2(reorder_tvalid_0_rep2),.O(N_285));
defparam desc3654.INIT=8'hCA;
  LUT3 desc3655(.I0(buffer_sreg[13:13]),.I1(buffer_sreg[15:15]),.I2(reorder_tvalid_0_rep2),.O(N_286));
defparam desc3655.INIT=8'hCA;
  LUT3 desc3656(.I0(buffer_sreg[10:10]),.I1(buffer_sreg[12:12]),.I2(reorder_tvalid_0_rep2),.O(N_283));
defparam desc3656.INIT=8'hCA;
  LUT3 desc3657(.I0(buffer_sreg[11:11]),.I1(buffer_sreg[13:13]),.I2(reorder_tvalid_0_rep2),.O(N_284));
defparam desc3657.INIT=8'hCA;
  LUT3 desc3658(.I0(buffer_sreg[8:8]),.I1(buffer_sreg[10:10]),.I2(reorder_tvalid_0_rep2),.O(N_281));
defparam desc3658.INIT=8'hCA;
  LUT3 desc3659(.I0(buffer_sreg[9:9]),.I1(buffer_sreg[11:11]),.I2(reorder_tvalid_0_rep2),.O(N_282));
defparam desc3659.INIT=8'hCA;
  LUT3 desc3660(.I0(buffer_sreg[7:7]),.I1(buffer_sreg[9:9]),.I2(reorder_tvalid_0_rep2),.O(N_280));
defparam desc3660.INIT=8'hCA;
  LUT3 desc3661(.I0(buffer_sreg[41:41]),.I1(buffer_sreg[43:43]),.I2(reorder_tvalid_0_rep2),.O(N_314));
defparam desc3661.INIT=8'hCA;
  LUT3 desc3662(.I0(buffer_sreg[5:5]),.I1(buffer_sreg[7:7]),.I2(reorder_tvalid_0_rep2),.O(N_278));
defparam desc3662.INIT=8'hCA;
  LUT3 desc3663(.I0(buffer_sreg[6:6]),.I1(buffer_sreg[8:8]),.I2(reorder_tvalid_0_rep2),.O(N_279));
defparam desc3663.INIT=8'hCA;
  LUT3 desc3664(.I0(buffer_sreg[4:4]),.I1(buffer_sreg[6:6]),.I2(reorder_tvalid_0_rep2),.O(N_277));
defparam desc3664.INIT=8'hCA;
  LUT3 desc3665(.I0(buffer_sreg[30:30]),.I1(buffer_sreg[32:32]),.I2(reorder_tvalid_0_rep2),.O(N_303));
defparam desc3665.INIT=8'hCA;
  LUT3 desc3666(.I0(buffer_sreg[2:2]),.I1(buffer_sreg[4:4]),.I2(reorder_tvalid_0_rep2),.O(N_275));
defparam desc3666.INIT=8'hCA;
  LUT3 desc3667(.I0(buffer_sreg[3:3]),.I1(buffer_sreg[5:5]),.I2(reorder_tvalid_0_rep2),.O(N_276));
defparam desc3667.INIT=8'hCA;
  LUT3 desc3668(.I0(buffer_sreg[2:2]),.I1(reorder_tdata),.I2(reorder_tvalid_0_rep2),.O(N_273));
defparam desc3668.INIT=8'hAC;
  LUT3 desc3669(.I0(buffer_sreg[1:1]),.I1(buffer_sreg[3:3]),.I2(reorder_tvalid_0_rep2),.O(N_274));
defparam desc3669.INIT=8'hCA;
  LUT3 desc3670(.I0(buffer_sreg[95:95]),.I1(buffer_sreg[93:93]),.I2(reorder_tvalid),.O(N_271));
defparam desc3670.INIT=8'hAC;
  LUT3 desc3671(.I0(buffer_sreg[92:92]),.I1(buffer_sreg[94:94]),.I2(reorder_tvalid),.O(N_346));
defparam desc3671.INIT=8'hCA;
  LUT3 desc3672(.I0(buffer_sreg[89:89]),.I1(buffer_sreg[91:91]),.I2(reorder_tvalid),.O(N_269));
defparam desc3672.INIT=8'hCA;
  LUT3 desc3673(.I0(buffer_sreg[90:90]),.I1(buffer_sreg[92:92]),.I2(reorder_tvalid),.O(N_345));
defparam desc3673.INIT=8'hCA;
  LUT3 desc3674(.I0(buffer_sreg[87:87]),.I1(buffer_sreg[89:89]),.I2(reorder_tvalid),.O(N_268));
defparam desc3674.INIT=8'hCA;
  LUT3 desc3675(.I0(buffer_sreg[86:86]),.I1(buffer_sreg[88:88]),.I2(reorder_tvalid),.O(N_343));
defparam desc3675.INIT=8'hCA;
  LUT3 desc3676(.I0(buffer_sreg[85:85]),.I1(buffer_sreg[87:87]),.I2(reorder_tvalid),.O(N_267));
defparam desc3676.INIT=8'hCA;
  LUT3 desc3677(.I0(buffer_sreg[84:84]),.I1(buffer_sreg[86:86]),.I2(reorder_tvalid),.O(N_342));
defparam desc3677.INIT=8'hCA;
  LUT3 desc3678(.I0(buffer_sreg[83:83]),.I1(buffer_sreg[85:85]),.I2(reorder_tvalid),.O(N_266));
defparam desc3678.INIT=8'hCA;
  LUT3 desc3679(.I0(buffer_sreg[91:91]),.I1(buffer_sreg[93:93]),.I2(reorder_tvalid),.O(N_270));
defparam desc3679.INIT=8'hCA;
  LUT3 desc3680(.I0(buffer_sreg[81:81]),.I1(buffer_sreg[83:83]),.I2(reorder_tvalid),.O(N_265));
defparam desc3680.INIT=8'hCA;
  LUT3 desc3681(.I0(buffer_sreg[82:82]),.I1(buffer_sreg[84:84]),.I2(reorder_tvalid),.O(N_341));
defparam desc3681.INIT=8'hCA;
  LUT3 desc3682(.I0(buffer_sreg[79:79]),.I1(buffer_sreg[81:81]),.I2(reorder_tvalid),.O(N_264));
defparam desc3682.INIT=8'hCA;
  LUT3 desc3683(.I0(buffer_sreg[78:78]),.I1(buffer_sreg[80:80]),.I2(reorder_tvalid),.O(N_339));
defparam desc3683.INIT=8'hCA;
  LUT3 desc3684(.I0(buffer_sreg[77:77]),.I1(buffer_sreg[79:79]),.I2(reorder_tvalid),.O(N_263));
defparam desc3684.INIT=8'hCA;
  LUT3 desc3685(.I0(buffer_sreg[76:76]),.I1(buffer_sreg[78:78]),.I2(reorder_tvalid),.O(N_338));
defparam desc3685.INIT=8'hCA;
  LUT3 desc3686(.I0(buffer_sreg[75:75]),.I1(buffer_sreg[77:77]),.I2(reorder_tvalid),.O(N_262));
defparam desc3686.INIT=8'hCA;
  LUT3 desc3687(.I0(buffer_sreg[74:74]),.I1(buffer_sreg[76:76]),.I2(reorder_tvalid),.O(N_337));
defparam desc3687.INIT=8'hCA;
  LUT3 desc3688(.I0(buffer_sreg[71:71]),.I1(buffer_sreg[73:73]),.I2(reorder_tvalid),.O(N_260));
defparam desc3688.INIT=8'hCA;
  LUT3 desc3689(.I0(buffer_sreg[72:72]),.I1(buffer_sreg[74:74]),.I2(reorder_tvalid),.O(N_336));
defparam desc3689.INIT=8'hCA;
  LUT3 desc3690(.I0(buffer_sreg[69:69]),.I1(buffer_sreg[71:71]),.I2(reorder_tvalid),.O(N_259));
defparam desc3690.INIT=8'hCA;
  LUT3 desc3691(.I0(buffer_sreg[70:70]),.I1(buffer_sreg[72:72]),.I2(reorder_tvalid),.O(N_335));
defparam desc3691.INIT=8'hCA;
  LUT3 desc3692(.I0(buffer_sreg[67:67]),.I1(buffer_sreg[69:69]),.I2(reorder_tvalid),.O(N_258));
defparam desc3692.INIT=8'hCA;
  LUT3 desc3693(.I0(buffer_sreg[68:68]),.I1(buffer_sreg[70:70]),.I2(reorder_tvalid),.O(N_334));
defparam desc3693.INIT=8'hCA;
  LUT3 desc3694(.I0(buffer_sreg[65:65]),.I1(buffer_sreg[67:67]),.I2(reorder_tvalid),.O(N_257));
defparam desc3694.INIT=8'hCA;
  LUT3 desc3695(.I0(buffer_sreg[66:66]),.I1(buffer_sreg[68:68]),.I2(reorder_tvalid),.O(N_333));
defparam desc3695.INIT=8'hCA;
  LUT3 desc3696(.I0(buffer_sreg[63:63]),.I1(buffer_sreg[65:65]),.I2(reorder_tvalid),.O(N_256));
defparam desc3696.INIT=8'hCA;
  LUT3 desc3697(.I0(buffer_sreg[64:64]),.I1(buffer_sreg[66:66]),.I2(reorder_tvalid),.O(N_332));
defparam desc3697.INIT=8'hCA;
  LUT3 desc3698(.I0(buffer_sreg[61:61]),.I1(buffer_sreg[63:63]),.I2(reorder_tvalid),.O(N_255));
defparam desc3698.INIT=8'hCA;
  LUT3 desc3699(.I0(buffer_sreg[60:60]),.I1(buffer_sreg[62:62]),.I2(reorder_tvalid),.O(N_330));
defparam desc3699.INIT=8'hCA;
  LUT3 desc3700(.I0(buffer_sreg[59:59]),.I1(buffer_sreg[61:61]),.I2(reorder_tvalid),.O(N_254));
defparam desc3700.INIT=8'hCA;
  LUT3 desc3701(.I0(buffer_sreg[58:58]),.I1(buffer_sreg[60:60]),.I2(reorder_tvalid),.O(N_329));
defparam desc3701.INIT=8'hCA;
  LUT3 desc3702(.I0(buffer_sreg[57:57]),.I1(buffer_sreg[59:59]),.I2(reorder_tvalid),.O(N_253));
defparam desc3702.INIT=8'hCA;
  LUT3 desc3703(.I0(buffer_sreg[56:56]),.I1(buffer_sreg[58:58]),.I2(reorder_tvalid),.O(N_328));
defparam desc3703.INIT=8'hCA;
  LUT3 desc3704(.I0(buffer_sreg[55:55]),.I1(buffer_sreg[57:57]),.I2(reorder_tvalid),.O(N_252));
defparam desc3704.INIT=8'hCA;
  LUT3 desc3705(.I0(buffer_sreg[62:62]),.I1(buffer_sreg[64:64]),.I2(reorder_tvalid),.O(N_331));
defparam desc3705.INIT=8'hCA;
  LUT2 un1_buffer_cnt_1_s_6_RNIL8A01_o6(.I0(N_357),.I1(un1_buffer_cnt_1_s_6_0),.O(N_71_i));
defparam un1_buffer_cnt_1_s_6_RNIL8A01_o6.INIT=4'h4;
  LUT4 un1_buffer_cnt_1_s_6_RNIL8A01_o5(.I0(traceback_last_tuser),.I1(traceback_tvalid),.I2(reorder_tvalid_0_rep2),.I3(N_357),.O(send_output_rep2));
defparam un1_buffer_cnt_1_s_6_RNIL8A01_o5.INIT=16'h08F8;
  LUT2 un1_buffer_cnt_1_s_5_RNI91131_o6(.I0(N_357),.I1(un1_buffer_cnt_1_s_5_0),.O(N_69_i));
defparam un1_buffer_cnt_1_s_5_RNI91131_o6.INIT=4'h4;
  LUT4 un1_buffer_cnt_1_s_5_RNI91131_o5(.I0(reorder_tvalid_fast),.I1(traceback_last_tuser),.I2(traceback_tvalid),.I3(N_357),.O(send_output_fast));
defparam un1_buffer_cnt_1_s_5_RNI91131_o5.INIT=16'h40EA;
  LUT2 un1_buffer_cnt_1_s_4_RNII8A01_o6(.I0(N_357),.I1(un1_buffer_cnt_1_s_4_0),.O(N_67_i));
defparam un1_buffer_cnt_1_s_4_RNII8A01_o6.INIT=4'h4;
  LUT4 un1_buffer_cnt_1_s_4_RNII8A01_o5(.I0(traceback_last_tuser),.I1(traceback_tvalid),.I2(reorder_tvalid_0_rep1),.I3(N_357),.O(send_output_rep1));
defparam un1_buffer_cnt_1_s_4_RNII8A01_o5.INIT=16'h08F8;
  LUT2 un1_buffer_cnt_1_s_1_RNITRFF_o6(.I0(N_357),.I1(un1_buffer_cnt_1_s_1_0),.O(N_61_i));
defparam un1_buffer_cnt_1_s_1_RNITRFF_o6.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_1_RNITRFF_o5(.I0(N_357),.I1(un1_buffer_cnt_1_s_3_0),.O(N_65_i));
defparam un1_buffer_cnt_1_s_1_RNITRFF_o5.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_2_RNI3INF_o6(.I0(N_357),.I1(un1_buffer_cnt_1_s_2_0),.O(N_63_i));
defparam un1_buffer_cnt_1_s_2_RNI3INF_o6.INIT=4'h4;
  LUT2 un1_buffer_cnt_1_s_2_RNI3INF_o5(.I0(un1_buffer_cnt_1_axb_0),.I1(N_357),.O(N_59_i));
defparam un1_buffer_cnt_1_s_2_RNI3INF_o5.INIT=4'h2;
endmodule
module dec_viterbi_inj (aclk,aresetn,s_axis_input_tvalid,s_axis_input_tdata,s_axis_input_tlast,s_axis_input_tready,m_axis_output_tvalid,m_axis_output_tdata,m_axis_output_tlast,m_axis_output_tready,s_axis_ctrl_tvalid,s_axis_ctrl_tdata,s_axis_ctrl_tlast,s_axis_ctrl_tready,p_desc95_p_O_FDacsZ0_,p_desc96_p_O_FDacsZ0_,p_desc134_p_O_FDacsZ0_1_,p_desc135_p_O_FDacsZ0_1_,p_desc173_p_O_FDacsZ0_2_,p_desc174_p_O_FDacsZ0_2_,p_desc212_p_O_FDacsZ0_3_,p_desc213_p_O_FDacsZ0_3_,p_desc251_p_O_FDacsZ0_4_,p_desc252_p_O_FDacsZ0_4_,p_desc290_p_O_FDacsZ0_5_,p_desc291_p_O_FDacsZ0_5_,p_desc329_p_O_FDacsZ0_6_,p_desc330_p_O_FDacsZ0_6_,p_desc368_p_O_FDacsZ0_7_,p_desc369_p_O_FDacsZ0_7_,p_desc407_p_O_FDacsZ0_8_,p_desc408_p_O_FDacsZ0_8_,p_desc446_p_O_FDacsZ0_9_,p_desc447_p_O_FDacsZ0_9_,p_desc485_p_O_FDacsZ0_10_,p_desc486_p_O_FDacsZ0_10_,p_desc524_p_O_FDacsZ0_11_,p_desc525_p_O_FDacsZ0_11_,p_desc563_p_O_FDacsZ0_12_,p_desc564_p_O_FDacsZ0_12_,p_desc602_p_O_FDacsZ0_13_,p_desc603_p_O_FDacsZ0_13_,p_desc641_p_O_FDacsZ0_14_,p_desc642_p_O_FDacsZ0_14_,p_desc680_p_O_FDacsZ0_15_,p_desc681_p_O_FDacsZ0_15_,p_desc719_p_O_FDacsZ0_16_,p_desc720_p_O_FDacsZ0_16_,p_desc758_p_O_FDacsZ0_17_,p_desc759_p_O_FDacsZ0_17_,p_desc797_p_O_FDacsZ0_18_,p_desc798_p_O_FDacsZ0_18_,p_desc873_p_O_FDacsZ0_20_,p_desc874_p_O_FDacsZ0_20_,p_desc912_p_O_FDacsZ0_21_,p_desc913_p_O_FDacsZ0_21_,p_desc989_p_O_FDacsZ0_22_,p_desc990_p_O_FDacsZ0_22_,p_desc1028_p_O_FDacsZ0_23_,p_desc1029_p_O_FDacsZ0_23_,p_desc1067_p_O_FDacsZ0_24_,p_desc1068_p_O_FDacsZ0_24_,p_desc1106_p_O_FDacsZ0_25_,p_desc1107_p_O_FDacsZ0_25_,p_desc1145_p_O_FDacsZ0_26_,p_desc1146_p_O_FDacsZ0_26_,p_desc1184_p_O_FDacsZ0_27_,p_desc1185_p_O_FDacsZ0_27_,p_desc1223_p_O_FDacsZ0_28_,p_desc1224_p_O_FDacsZ0_28_,p_desc1262_p_O_FDacsZ0_29_,p_desc1263_p_O_FDacsZ0_29_,p_desc1301_p_O_FDacsZ0_30_,p_desc1302_p_O_FDacsZ0_30_,p_desc1340_p_O_FDacsZ0_31_,p_desc1341_p_O_FDacsZ0_31_,p_desc1379_p_O_FDacsZ0_32_,p_desc1380_p_O_FDacsZ0_32_,p_desc1418_p_O_FDacsZ0_33_,p_desc1419_p_O_FDacsZ0_33_,p_desc1457_p_O_FDacsZ0_34_,p_desc1458_p_O_FDacsZ0_34_,p_desc1496_p_O_FDacsZ0_35_,p_desc1497_p_O_FDacsZ0_35_,p_desc1535_p_O_FDacsZ0_36_,p_desc1536_p_O_FDacsZ0_36_,p_desc1574_p_O_FDacsZ0_37_,p_desc1575_p_O_FDacsZ0_37_,p_desc1613_p_O_FDacsZ0_38_,p_desc1614_p_O_FDacsZ0_38_,p_desc1652_p_O_FDacsZ0_39_,p_desc1653_p_O_FDacsZ0_39_,p_desc1691_p_O_FDacsZ0_40_,p_desc1692_p_O_FDacsZ0_40_,p_desc1730_p_O_FDacsZ0_41_,p_desc1731_p_O_FDacsZ0_41_,p_desc1769_p_O_FDacsZ0_42_,p_desc1770_p_O_FDacsZ0_42_,p_desc1808_p_O_FDacsZ0_43_,p_desc1809_p_O_FDacsZ0_43_,p_desc1847_p_O_FDacsZ0_44_,p_desc1848_p_O_FDacsZ0_44_,p_desc1886_p_O_FDacsZ0_45_,p_desc1887_p_O_FDacsZ0_45_,p_desc1925_p_O_FDacsZ0_46_,p_desc1926_p_O_FDacsZ0_46_,p_desc1964_p_O_FDacsZ0_47_,p_desc1965_p_O_FDacsZ0_47_,p_desc2003_p_O_FDacsZ0_48_,p_desc2004_p_O_FDacsZ0_48_,p_desc2042_p_O_FDacsZ0_49_,p_desc2043_p_O_FDacsZ0_49_,p_desc2081_p_O_FDacsZ0_50_,p_desc2082_p_O_FDacsZ0_50_,p_desc2120_p_O_FDacsZ0_51_,p_desc2121_p_O_FDacsZ0_51_,p_desc2159_p_O_FDacsZ0_52_,p_desc2160_p_O_FDacsZ0_52_,p_desc2198_p_O_FDacsZ0_53_,p_desc2199_p_O_FDacsZ0_53_,p_desc2237_p_O_FDacsZ0_54_,p_desc2238_p_O_FDacsZ0_54_,p_desc2276_p_O_FDacsZ0_55_,p_desc2277_p_O_FDacsZ0_55_,p_desc2315_p_O_FDacsZ0_56_,p_desc2316_p_O_FDacsZ0_56_,p_desc2354_p_O_FDacsZ0_57_,p_desc2355_p_O_FDacsZ0_57_,p_desc2393_p_O_FDacsZ0_58_,p_desc2394_p_O_FDacsZ0_58_,p_desc2432_p_O_FDacsZ0_59_,p_desc2433_p_O_FDacsZ0_59_,p_desc2471_p_O_FDacsZ0_60_,p_desc2472_p_O_FDacsZ0_60_,p_desc2510_p_O_FDacsZ0_61_,p_desc2511_p_O_FDacsZ0_61_,p_desc2549_p_O_FDacsZ0_62_,p_desc2550_p_O_FDacsZ0_62_,p_m_axis_output_tdata_0_rep2_Z_p_O_FDREbranch_distanceZ3_,p_m_axis_output_tdata_0_rep1_Z_p_O_FDREbranch_distanceZ3_,p_desc31_p_O_FDREbranch_distanceZ3_,p_desc32_p_O_FDREbranch_distanceZ3_,p_desc33_p_O_FDREbranch_distanceZ3_,p_desc34_p_O_FDREbranch_distanceZ3_,p_desc35_p_O_FDREbranch_distanceZ3_,p_desc36_p_O_FDREbranch_distanceZ3_,p_desc37_p_O_FDREbranch_distanceZ3_,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ2_,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ2_,p_desc39_p_O_FDREbranch_distanceZ2_,p_desc52_p_O_FDREbranch_distanceZ2_,p_desc53_p_O_FDREbranch_distanceZ2_,p_desc54_p_O_FDREbranch_distanceZ2_,p_desc55_p_O_FDREbranch_distanceZ2_,p_desc56_p_O_FDREbranch_distanceZ2_,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ0_,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ0_,p_desc63_p_O_FDREbranch_distanceZ0_,p_desc78_p_O_FDREbranch_distanceZ0_,p_desc79_p_O_FDREbranch_distanceZ0_,p_desc80_p_O_FDREbranch_distanceZ0_,p_desc81_p_O_FDREbranch_distanceZ0_,p_desc82_p_O_FDREbranch_distanceZ0_,p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ1_,p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ1_,p_desc83_p_O_FDREbranch_distanceZ1_,p_desc84_p_O_FDREbranch_distanceZ1_,p_desc85_p_O_FDREbranch_distanceZ1_,p_desc86_p_O_FDREbranch_distanceZ1_,p_desc87_p_O_FDREbranch_distanceZ1_,p_desc88_p_O_FDREbranch_distanceZ1_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_,p_desc125_p_O_FDREacsZ0_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_1_,p_desc164_p_O_FDREacsZ0_1_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_2_,p_desc203_p_O_FDREacsZ0_2_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_3_,p_desc242_p_O_FDREacsZ0_3_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_4_,p_desc281_p_O_FDREacsZ0_4_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_5_,p_desc320_p_O_FDREacsZ0_5_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_6_,p_desc359_p_O_FDREacsZ0_6_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_7_,p_desc398_p_O_FDREacsZ0_7_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_8_,p_desc437_p_O_FDREacsZ0_8_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_9_,p_desc476_p_O_FDREacsZ0_9_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_10_,p_desc515_p_O_FDREacsZ0_10_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_11_,p_desc554_p_O_FDREacsZ0_11_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_12_,p_desc593_p_O_FDREacsZ0_12_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_13_,p_desc632_p_O_FDREacsZ0_13_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_14_,p_desc671_p_O_FDREacsZ0_14_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_15_,p_desc710_p_O_FDREacsZ0_15_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_16_,p_desc749_p_O_FDREacsZ0_16_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_17_,p_desc788_p_O_FDREacsZ0_17_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_18_,p_desc827_p_O_FDREacsZ0_18_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_19_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_20_,p_desc903_p_O_FDREacsZ0_20_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_21_,p_desc942_p_O_FDREacsZ0_21_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_22_,p_desc1019_p_O_FDREacsZ0_22_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_23_,p_desc1058_p_O_FDREacsZ0_23_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_24_,p_desc1097_p_O_FDREacsZ0_24_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_25_,p_desc1136_p_O_FDREacsZ0_25_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_26_,p_desc1175_p_O_FDREacsZ0_26_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_27_,p_desc1214_p_O_FDREacsZ0_27_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_28_,p_desc1253_p_O_FDREacsZ0_28_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_29_,p_desc1292_p_O_FDREacsZ0_29_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_30_,p_desc1331_p_O_FDREacsZ0_30_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_31_,p_desc1370_p_O_FDREacsZ0_31_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_32_,p_desc1409_p_O_FDREacsZ0_32_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_33_,p_desc1448_p_O_FDREacsZ0_33_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_34_,p_desc1487_p_O_FDREacsZ0_34_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_35_,p_desc1526_p_O_FDREacsZ0_35_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_36_,p_desc1565_p_O_FDREacsZ0_36_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_37_,p_desc1604_p_O_FDREacsZ0_37_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_38_,p_desc1643_p_O_FDREacsZ0_38_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_39_,p_desc1682_p_O_FDREacsZ0_39_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_40_,p_desc1721_p_O_FDREacsZ0_40_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_41_,p_desc1760_p_O_FDREacsZ0_41_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_42_,p_desc1799_p_O_FDREacsZ0_42_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_43_,p_desc1838_p_O_FDREacsZ0_43_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_44_,p_desc1877_p_O_FDREacsZ0_44_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_45_,p_desc1916_p_O_FDREacsZ0_45_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_46_,p_desc1955_p_O_FDREacsZ0_46_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_47_,p_desc1994_p_O_FDREacsZ0_47_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_48_,p_desc2033_p_O_FDREacsZ0_48_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_49_,p_desc2072_p_O_FDREacsZ0_49_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_50_,p_desc2111_p_O_FDREacsZ0_50_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_51_,p_desc2150_p_O_FDREacsZ0_51_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_52_,p_desc2189_p_O_FDREacsZ0_52_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_53_,p_desc2228_p_O_FDREacsZ0_53_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_54_,p_desc2267_p_O_FDREacsZ0_54_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_55_,p_desc2306_p_O_FDREacsZ0_55_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_56_,p_desc2345_p_O_FDREacsZ0_56_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_57_,p_desc2384_p_O_FDREacsZ0_57_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_58_,p_desc2423_p_O_FDREacsZ0_58_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_59_,p_desc2462_p_O_FDREacsZ0_59_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_60_,p_desc2501_p_O_FDREacsZ0_60_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_61_,p_desc2540_p_O_FDREacsZ0_61_,p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_62_,p_desc2579_p_O_FDREacsZ0_62_);
input aclk ;
input aresetn ;
input s_axis_input_tvalid ;
input [31:0] s_axis_input_tdata ;
input s_axis_input_tlast ;
output s_axis_input_tready ;
output m_axis_output_tvalid ;
output m_axis_output_tdata ;
output m_axis_output_tlast ;
input m_axis_output_tready ;
input s_axis_ctrl_tvalid ;
input [31:0] s_axis_ctrl_tdata ;
input s_axis_ctrl_tlast ;
output s_axis_ctrl_tready ;
wire aclk ;
wire aresetn ;
wire s_axis_input_tvalid ;
wire s_axis_input_tlast ;
wire s_axis_input_tready ;
wire m_axis_output_tvalid ;
wire m_axis_output_tdata ;
wire m_axis_output_tlast ;
wire m_axis_output_tready ;
wire s_axis_ctrl_tvalid ;
wire s_axis_ctrl_tlast ;
wire s_axis_ctrl_tready ;
wire [11:0] buffer_tdata ;
wire [5:0] branch_tdata_3 ;
wire [5:0] branch_tdata_2 ;
wire branch_tvalid ;
wire [5:0] branch_tdata_0 ;
wire branch_tlast ;
wire [5:0] branch_tdata_1 ;
wire [8:0] acs_prob_tdata_50 ;
wire [8:0] acs_prob_tdata_51 ;
wire [8:0] acs_prob_tdata_57 ;
wire [63:0] acs_dec_tdata ;
wire [8:0] acs_prob_tdata_24 ;
wire [8:0] acs_prob_tdata_25 ;
wire [8:0] acs_prob_tdata_12 ;
wire [8:0] acs_prob_tdata_44 ;
wire [8:0] acs_prob_tdata_45 ;
wire [8:0] acs_prob_tdata_54 ;
wire [8:0] acs_prob_tdata_20 ;
wire [8:0] acs_prob_tdata_21 ;
wire [8:0] acs_prob_tdata_42 ;
wire [8:0] acs_prob_tdata_48 ;
wire [8:0] acs_prob_tdata_49 ;
wire [8:0] acs_prob_tdata_32 ;
wire [8:0] acs_prob_tdata_33 ;
wire [8:0] acs_prob_tdata_16 ;
wire [8:0] acs_prob_tdata_2 ;
wire [8:0] acs_prob_tdata_3 ;
wire [8:0] acs_prob_tdata_1 ;
wire [8:0] acs_prob_tdata_36 ;
wire [8:0] acs_prob_tdata_37 ;
wire [8:0] acs_prob_tdata_18 ;
wire [8:0] acs_prob_tdata_6 ;
wire [8:0] acs_prob_tdata_7 ;
wire [8:0] acs_prob_tdata_60 ;
wire [8:0] acs_prob_tdata_61 ;
wire [8:0] acs_prob_tdata_62 ;
wire [8:0] acs_prob_tdata_30 ;
wire [8:0] acs_prob_tdata_31 ;
wire [8:0] acs_prob_tdata_47 ;
wire [8:0] acs_prob_tdata_10 ;
wire [8:0] acs_prob_tdata_11 ;
wire [8:0] acs_prob_tdata_5 ;
wire [8:0] acs_prob_tdata_34 ;
wire [8:0] acs_prob_tdata_35 ;
wire [8:0] acs_prob_tdata_4 ;
wire [8:0] acs_prob_tdata_38 ;
wire [8:0] acs_prob_tdata_39 ;
wire [8:0] acs_prob_tdata_19 ;
wire [8:0] acs_prob_tdata_8 ;
wire [8:0] acs_prob_tdata_9 ;
wire [8:0] acs_prob_tdata_63 ;
wire [8:0] acs_prob_tdata_58 ;
wire [8:0] acs_prob_tdata_59 ;
wire [8:0] acs_prob_tdata_0 ;
wire acs_tvalid ;
wire acs_tlast ;
wire [8:0] acs_prob_tdata_28 ;
wire [8:0] acs_prob_tdata_29 ;
wire [8:0] acs_prob_tdata_46 ;
wire [8:0] acs_prob_tdata_40 ;
wire [8:0] acs_prob_tdata_41 ;
wire [8:0] acs_prob_tdata_52 ;
wire [8:0] acs_prob_tdata_22 ;
wire [8:0] acs_prob_tdata_14 ;
wire [8:0] acs_prob_tdata_15 ;
wire [8:0] acs_prob_tdata_43 ;
wire [8:0] acs_prob_tdata_53 ;
wire [8:0] acs_prob_tdata_23 ;
wire [8:0] acs_prob_tdata_17 ;
wire [8:0] acs_prob_tdata_13 ;
wire [8:0] acs_prob_tdata_26 ;
wire [8:0] acs_prob_tdata_55 ;
wire [8:0] acs_prob_tdata_27 ;
wire [8:0] acs_prob_tdata_56 ;
wire [1:0] ram_tvalid ;
wire [1:0] ram_tlast ;
wire [1:0] ram_window_tuser ;
wire [1:0] ram_last_tuser ;
wire [1:0] traceback_tvalid ;
wire [1:0] traceback_tdata ;
wire [1:0] traceback_tlast ;
wire [1:0] traceback_last_tuser ;
wire [1:0] reorder_last_tuser ;
wire reorder_tvalid ;
wire reorder_tdata ;
wire current_active ;
wire [2:0] \gen_inst_reorder.0.inst_reorder.buffer_cnt  ;
wire [2:0] \gen_inst_reorder.1.inst_reorder.buffer_cnt  ;
wire [4:0] \inst_ram_ctrl.write_ram_fsm  ;
wire [63:0] \inst_ram_ctrl.pr_buf_ram_output.0.ram_buffer_0_2  ;
wire [63:0] \inst_ram_ctrl.pr_buf_ram_output.1.ram_buffer_1_1  ;
wire [63:0] \inst_ram_ctrl.ram_buffer_0  ;
wire [63:0] \inst_ram_ctrl.ram_buffer_1  ;
wire [1:0] \inst_ram_ctrl.ram_buffer_full  ;
wire [3:1] buffer_tdata_i ;
wire current_active_0 ;
wire [1:0] reorder_tvalid_fast ;
wire branch_tdata_0_fast ;
wire branch_tdata_2_fast ;
wire branch_tdata_3_fast ;
wire branch_tdata_1_fast ;
wire buffer_tvalid ;
wire buffer_tlast ;
wire VCC ;
wire GND ;
wire \inst_axi4s_buffer.pr_reg.un1_output_accept  ;
wire \gen_inst_reorder.0.inst_reorder.last_window  ;
wire \gen_inst_reorder.1.inst_reorder.last_window  ;
wire \inst_ram_ctrl.pr_write_ram.un1_s_axis_input_tvalid  ;
wire N_104 ;
wire N_130 ;
wire \inst_ram_ctrl.N_1756_1  ;
wire \inst_ram_ctrl.un27_s_axis_input_tready_int  ;
wire N_129 ;
wire aresetn_i ;
wire N_2388_i ;
wire N_99 ;
wire \pr_buf_ram_output.1.un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5  ;
wire s_axis_inbranch_tlast_d_RNIIAVE1_O5 ;
wire reorder_tvalid_0_rep1 ;
wire reorder_tvalid_0_rep2 ;
wire \inst_ram_ctrl.write_ram_fsm_4_rep1  ;
wire \inst_ram_ctrl.write_ram_fsm_4_rep2  ;
wire \inst_ram_ctrl.write_ram_fsm_0_rep1  ;
wire \inst_ram_ctrl.write_ram_fsm_0_rep2  ;
wire branch_tdata_0_0_rep1 ;
wire branch_tdata_0_0_rep2 ;
wire \gen_branch_distance.2.inst_branch_distance.v_branch_result.v_branch_result_axb_0_i_fast  ;
wire branch_tdata_2_0_rep1 ;
wire branch_tdata_2_0_rep2 ;
wire branch_tdata_3_0_rep1 ;
wire branch_tdata_3_0_rep2 ;
wire \gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_fast  ;
wire branch_tdata_1_0_rep1 ;
wire \gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep1  ;
wire branch_tdata_1_0_rep2 ;
wire \gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep2  ;
wire reorder_tvalid_1_rep1 ;
wire \gen_inst_reorder.1.inst_reorder.send_output_rep1  ;
input p_desc95_p_O_FDacsZ0_ ;
input p_desc96_p_O_FDacsZ0_ ;
input p_desc134_p_O_FDacsZ0_1_ ;
input p_desc135_p_O_FDacsZ0_1_ ;
input p_desc173_p_O_FDacsZ0_2_ ;
input p_desc174_p_O_FDacsZ0_2_ ;
input p_desc212_p_O_FDacsZ0_3_ ;
input p_desc213_p_O_FDacsZ0_3_ ;
input p_desc251_p_O_FDacsZ0_4_ ;
input p_desc252_p_O_FDacsZ0_4_ ;
input p_desc290_p_O_FDacsZ0_5_ ;
input p_desc291_p_O_FDacsZ0_5_ ;
input p_desc329_p_O_FDacsZ0_6_ ;
input p_desc330_p_O_FDacsZ0_6_ ;
input p_desc368_p_O_FDacsZ0_7_ ;
input p_desc369_p_O_FDacsZ0_7_ ;
input p_desc407_p_O_FDacsZ0_8_ ;
input p_desc408_p_O_FDacsZ0_8_ ;
input p_desc446_p_O_FDacsZ0_9_ ;
input p_desc447_p_O_FDacsZ0_9_ ;
input p_desc485_p_O_FDacsZ0_10_ ;
input p_desc486_p_O_FDacsZ0_10_ ;
input p_desc524_p_O_FDacsZ0_11_ ;
input p_desc525_p_O_FDacsZ0_11_ ;
input p_desc563_p_O_FDacsZ0_12_ ;
input p_desc564_p_O_FDacsZ0_12_ ;
input p_desc602_p_O_FDacsZ0_13_ ;
input p_desc603_p_O_FDacsZ0_13_ ;
input p_desc641_p_O_FDacsZ0_14_ ;
input p_desc642_p_O_FDacsZ0_14_ ;
input p_desc680_p_O_FDacsZ0_15_ ;
input p_desc681_p_O_FDacsZ0_15_ ;
input p_desc719_p_O_FDacsZ0_16_ ;
input p_desc720_p_O_FDacsZ0_16_ ;
input p_desc758_p_O_FDacsZ0_17_ ;
input p_desc759_p_O_FDacsZ0_17_ ;
input p_desc797_p_O_FDacsZ0_18_ ;
input p_desc798_p_O_FDacsZ0_18_ ;
input p_desc873_p_O_FDacsZ0_20_ ;
input p_desc874_p_O_FDacsZ0_20_ ;
input p_desc912_p_O_FDacsZ0_21_ ;
input p_desc913_p_O_FDacsZ0_21_ ;
input p_desc989_p_O_FDacsZ0_22_ ;
input p_desc990_p_O_FDacsZ0_22_ ;
input p_desc1028_p_O_FDacsZ0_23_ ;
input p_desc1029_p_O_FDacsZ0_23_ ;
input p_desc1067_p_O_FDacsZ0_24_ ;
input p_desc1068_p_O_FDacsZ0_24_ ;
input p_desc1106_p_O_FDacsZ0_25_ ;
input p_desc1107_p_O_FDacsZ0_25_ ;
input p_desc1145_p_O_FDacsZ0_26_ ;
input p_desc1146_p_O_FDacsZ0_26_ ;
input p_desc1184_p_O_FDacsZ0_27_ ;
input p_desc1185_p_O_FDacsZ0_27_ ;
input p_desc1223_p_O_FDacsZ0_28_ ;
input p_desc1224_p_O_FDacsZ0_28_ ;
input p_desc1262_p_O_FDacsZ0_29_ ;
input p_desc1263_p_O_FDacsZ0_29_ ;
input p_desc1301_p_O_FDacsZ0_30_ ;
input p_desc1302_p_O_FDacsZ0_30_ ;
input p_desc1340_p_O_FDacsZ0_31_ ;
input p_desc1341_p_O_FDacsZ0_31_ ;
input p_desc1379_p_O_FDacsZ0_32_ ;
input p_desc1380_p_O_FDacsZ0_32_ ;
input p_desc1418_p_O_FDacsZ0_33_ ;
input p_desc1419_p_O_FDacsZ0_33_ ;
input p_desc1457_p_O_FDacsZ0_34_ ;
input p_desc1458_p_O_FDacsZ0_34_ ;
input p_desc1496_p_O_FDacsZ0_35_ ;
input p_desc1497_p_O_FDacsZ0_35_ ;
input p_desc1535_p_O_FDacsZ0_36_ ;
input p_desc1536_p_O_FDacsZ0_36_ ;
input p_desc1574_p_O_FDacsZ0_37_ ;
input p_desc1575_p_O_FDacsZ0_37_ ;
input p_desc1613_p_O_FDacsZ0_38_ ;
input p_desc1614_p_O_FDacsZ0_38_ ;
input p_desc1652_p_O_FDacsZ0_39_ ;
input p_desc1653_p_O_FDacsZ0_39_ ;
input p_desc1691_p_O_FDacsZ0_40_ ;
input p_desc1692_p_O_FDacsZ0_40_ ;
input p_desc1730_p_O_FDacsZ0_41_ ;
input p_desc1731_p_O_FDacsZ0_41_ ;
input p_desc1769_p_O_FDacsZ0_42_ ;
input p_desc1770_p_O_FDacsZ0_42_ ;
input p_desc1808_p_O_FDacsZ0_43_ ;
input p_desc1809_p_O_FDacsZ0_43_ ;
input p_desc1847_p_O_FDacsZ0_44_ ;
input p_desc1848_p_O_FDacsZ0_44_ ;
input p_desc1886_p_O_FDacsZ0_45_ ;
input p_desc1887_p_O_FDacsZ0_45_ ;
input p_desc1925_p_O_FDacsZ0_46_ ;
input p_desc1926_p_O_FDacsZ0_46_ ;
input p_desc1964_p_O_FDacsZ0_47_ ;
input p_desc1965_p_O_FDacsZ0_47_ ;
input p_desc2003_p_O_FDacsZ0_48_ ;
input p_desc2004_p_O_FDacsZ0_48_ ;
input p_desc2042_p_O_FDacsZ0_49_ ;
input p_desc2043_p_O_FDacsZ0_49_ ;
input p_desc2081_p_O_FDacsZ0_50_ ;
input p_desc2082_p_O_FDacsZ0_50_ ;
input p_desc2120_p_O_FDacsZ0_51_ ;
input p_desc2121_p_O_FDacsZ0_51_ ;
input p_desc2159_p_O_FDacsZ0_52_ ;
input p_desc2160_p_O_FDacsZ0_52_ ;
input p_desc2198_p_O_FDacsZ0_53_ ;
input p_desc2199_p_O_FDacsZ0_53_ ;
input p_desc2237_p_O_FDacsZ0_54_ ;
input p_desc2238_p_O_FDacsZ0_54_ ;
input p_desc2276_p_O_FDacsZ0_55_ ;
input p_desc2277_p_O_FDacsZ0_55_ ;
input p_desc2315_p_O_FDacsZ0_56_ ;
input p_desc2316_p_O_FDacsZ0_56_ ;
input p_desc2354_p_O_FDacsZ0_57_ ;
input p_desc2355_p_O_FDacsZ0_57_ ;
input p_desc2393_p_O_FDacsZ0_58_ ;
input p_desc2394_p_O_FDacsZ0_58_ ;
input p_desc2432_p_O_FDacsZ0_59_ ;
input p_desc2433_p_O_FDacsZ0_59_ ;
input p_desc2471_p_O_FDacsZ0_60_ ;
input p_desc2472_p_O_FDacsZ0_60_ ;
input p_desc2510_p_O_FDacsZ0_61_ ;
input p_desc2511_p_O_FDacsZ0_61_ ;
input p_desc2549_p_O_FDacsZ0_62_ ;
input p_desc2550_p_O_FDacsZ0_62_ ;
input p_m_axis_output_tdata_0_rep2_Z_p_O_FDREbranch_distanceZ3_ ;
input p_m_axis_output_tdata_0_rep1_Z_p_O_FDREbranch_distanceZ3_ ;
input p_desc31_p_O_FDREbranch_distanceZ3_ ;
input p_desc32_p_O_FDREbranch_distanceZ3_ ;
input p_desc33_p_O_FDREbranch_distanceZ3_ ;
input p_desc34_p_O_FDREbranch_distanceZ3_ ;
input p_desc35_p_O_FDREbranch_distanceZ3_ ;
input p_desc36_p_O_FDREbranch_distanceZ3_ ;
input p_desc37_p_O_FDREbranch_distanceZ3_ ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ2_ ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ2_ ;
input p_desc39_p_O_FDREbranch_distanceZ2_ ;
input p_desc52_p_O_FDREbranch_distanceZ2_ ;
input p_desc53_p_O_FDREbranch_distanceZ2_ ;
input p_desc54_p_O_FDREbranch_distanceZ2_ ;
input p_desc55_p_O_FDREbranch_distanceZ2_ ;
input p_desc56_p_O_FDREbranch_distanceZ2_ ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ0_ ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ0_ ;
input p_desc63_p_O_FDREbranch_distanceZ0_ ;
input p_desc78_p_O_FDREbranch_distanceZ0_ ;
input p_desc79_p_O_FDREbranch_distanceZ0_ ;
input p_desc80_p_O_FDREbranch_distanceZ0_ ;
input p_desc81_p_O_FDREbranch_distanceZ0_ ;
input p_desc82_p_O_FDREbranch_distanceZ0_ ;
input p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ1_ ;
input p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ1_ ;
input p_desc83_p_O_FDREbranch_distanceZ1_ ;
input p_desc84_p_O_FDREbranch_distanceZ1_ ;
input p_desc85_p_O_FDREbranch_distanceZ1_ ;
input p_desc86_p_O_FDREbranch_distanceZ1_ ;
input p_desc87_p_O_FDREbranch_distanceZ1_ ;
input p_desc88_p_O_FDREbranch_distanceZ1_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_ ;
input p_desc125_p_O_FDREacsZ0_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_1_ ;
input p_desc164_p_O_FDREacsZ0_1_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_2_ ;
input p_desc203_p_O_FDREacsZ0_2_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_3_ ;
input p_desc242_p_O_FDREacsZ0_3_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_4_ ;
input p_desc281_p_O_FDREacsZ0_4_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_5_ ;
input p_desc320_p_O_FDREacsZ0_5_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_6_ ;
input p_desc359_p_O_FDREacsZ0_6_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_7_ ;
input p_desc398_p_O_FDREacsZ0_7_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_8_ ;
input p_desc437_p_O_FDREacsZ0_8_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_9_ ;
input p_desc476_p_O_FDREacsZ0_9_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_10_ ;
input p_desc515_p_O_FDREacsZ0_10_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_11_ ;
input p_desc554_p_O_FDREacsZ0_11_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_12_ ;
input p_desc593_p_O_FDREacsZ0_12_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_13_ ;
input p_desc632_p_O_FDREacsZ0_13_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_14_ ;
input p_desc671_p_O_FDREacsZ0_14_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_15_ ;
input p_desc710_p_O_FDREacsZ0_15_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_16_ ;
input p_desc749_p_O_FDREacsZ0_16_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_17_ ;
input p_desc788_p_O_FDREacsZ0_17_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_18_ ;
input p_desc827_p_O_FDREacsZ0_18_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_19_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_20_ ;
input p_desc903_p_O_FDREacsZ0_20_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_21_ ;
input p_desc942_p_O_FDREacsZ0_21_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_22_ ;
input p_desc1019_p_O_FDREacsZ0_22_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_23_ ;
input p_desc1058_p_O_FDREacsZ0_23_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_24_ ;
input p_desc1097_p_O_FDREacsZ0_24_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_25_ ;
input p_desc1136_p_O_FDREacsZ0_25_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_26_ ;
input p_desc1175_p_O_FDREacsZ0_26_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_27_ ;
input p_desc1214_p_O_FDREacsZ0_27_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_28_ ;
input p_desc1253_p_O_FDREacsZ0_28_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_29_ ;
input p_desc1292_p_O_FDREacsZ0_29_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_30_ ;
input p_desc1331_p_O_FDREacsZ0_30_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_31_ ;
input p_desc1370_p_O_FDREacsZ0_31_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_32_ ;
input p_desc1409_p_O_FDREacsZ0_32_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_33_ ;
input p_desc1448_p_O_FDREacsZ0_33_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_34_ ;
input p_desc1487_p_O_FDREacsZ0_34_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_35_ ;
input p_desc1526_p_O_FDREacsZ0_35_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_36_ ;
input p_desc1565_p_O_FDREacsZ0_36_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_37_ ;
input p_desc1604_p_O_FDREacsZ0_37_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_38_ ;
input p_desc1643_p_O_FDREacsZ0_38_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_39_ ;
input p_desc1682_p_O_FDREacsZ0_39_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_40_ ;
input p_desc1721_p_O_FDREacsZ0_40_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_41_ ;
input p_desc1760_p_O_FDREacsZ0_41_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_42_ ;
input p_desc1799_p_O_FDREacsZ0_42_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_43_ ;
input p_desc1838_p_O_FDREacsZ0_43_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_44_ ;
input p_desc1877_p_O_FDREacsZ0_44_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_45_ ;
input p_desc1916_p_O_FDREacsZ0_45_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_46_ ;
input p_desc1955_p_O_FDREacsZ0_46_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_47_ ;
input p_desc1994_p_O_FDREacsZ0_47_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_48_ ;
input p_desc2033_p_O_FDREacsZ0_48_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_49_ ;
input p_desc2072_p_O_FDREacsZ0_49_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_50_ ;
input p_desc2111_p_O_FDREacsZ0_50_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_51_ ;
input p_desc2150_p_O_FDREacsZ0_51_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_52_ ;
input p_desc2189_p_O_FDREacsZ0_52_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_53_ ;
input p_desc2228_p_O_FDREacsZ0_53_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_54_ ;
input p_desc2267_p_O_FDREacsZ0_54_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_55_ ;
input p_desc2306_p_O_FDREacsZ0_55_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_56_ ;
input p_desc2345_p_O_FDREacsZ0_56_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_57_ ;
input p_desc2384_p_O_FDREacsZ0_57_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_58_ ;
input p_desc2423_p_O_FDREacsZ0_58_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_59_ ;
input p_desc2462_p_O_FDREacsZ0_59_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_60_ ;
input p_desc2501_p_O_FDREacsZ0_60_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_61_ ;
input p_desc2540_p_O_FDREacsZ0_61_ ;
input p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_62_ ;
input p_desc2579_p_O_FDREacsZ0_62_ ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  FDR desc3706(.Q(current_active),.D(current_active_0),.C(aclk),.R(aresetn_i));
  LUT6_L desc3707(.I0(m_axis_output_tready),.I1(reorder_last_tuser[0:0]),.I2(reorder_last_tuser[1:1]),.I3(current_active),.I4(reorder_tvalid_0_rep1),.I5(reorder_tvalid_1_rep1),.LO(current_active_0));
defparam desc3707.INIT=64'h5F885F00FF88FF00;
  axi4s_buffer_inj inst_axi4s_buffer(.buffer_tdata_i(buffer_tdata_i[3:1]),.acs_tvalid(acs_tvalid),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.s_axis_input_tdata_0(s_axis_input_tdata[0:0]),.s_axis_input_tdata_1(s_axis_input_tdata[1:1]),.s_axis_input_tdata_2(s_axis_input_tdata[2:2]),.s_axis_input_tdata_3(s_axis_input_tdata[3:3]),.s_axis_input_tdata_8(s_axis_input_tdata[8:8]),.s_axis_input_tdata_9(s_axis_input_tdata[9:9]),.s_axis_input_tdata_10(s_axis_input_tdata[10:10]),.s_axis_input_tdata_11(s_axis_input_tdata[11:11]),.buffer_tdata_3(buffer_tdata[3:3]),.buffer_tdata_2(buffer_tdata[2:2]),.buffer_tdata_1(buffer_tdata[1:1]),.buffer_tdata_10(buffer_tdata[10:10]),.buffer_tdata_9(buffer_tdata[9:9]),.buffer_tdata_11(buffer_tdata[11:11]),.buffer_tdata_8(buffer_tdata[8:8]),.buffer_tdata_0(buffer_tdata[0:0]),.s_axis_input_tready(s_axis_input_tready),.aclk(aclk),.aresetn_i(aresetn_i),.buffer_tvalid(buffer_tvalid),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.s_axis_input_tvalid(s_axis_input_tvalid),.s_axis_input_tlast(s_axis_input_tlast),.N_2388_i(N_2388_i),.buffer_tlast(buffer_tlast));
  branch_distanceZ3_inj desc3708(.branch_tdata_3_fast(branch_tdata_3_fast),.buffer_tdata_0(buffer_tdata[0:0]),.buffer_tdata_8(buffer_tdata[8:8]),.buffer_tdata_1(buffer_tdata[1:1]),.buffer_tdata_9(buffer_tdata[9:9]),.buffer_tdata_10(buffer_tdata[10:10]),.buffer_tdata_11(buffer_tdata[11:11]),.buffer_tdata_3(buffer_tdata[3:3]),.buffer_tdata_2(buffer_tdata[2:2]),.buffer_tdata_i(buffer_tdata_i[3:1]),.branch_tdata_3(branch_tdata_3[5:0]),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.aclk(aclk),.aresetn_i(aresetn_i),.un1_output_accept(\inst_axi4s_buffer.pr_reg.un1_output_accept ),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.N_2388_i(N_2388_i),.p_m_axis_output_tdata_0_rep2_Z_p_O_FDRE(p_m_axis_output_tdata_0_rep2_Z_p_O_FDREbranch_distanceZ3_),.p_m_axis_output_tdata_0_rep1_Z_p_O_FDRE(p_m_axis_output_tdata_0_rep1_Z_p_O_FDREbranch_distanceZ3_),.p_desc31_p_O_FDRE(p_desc31_p_O_FDREbranch_distanceZ3_),.p_desc32_p_O_FDRE(p_desc32_p_O_FDREbranch_distanceZ3_),.p_desc33_p_O_FDRE(p_desc33_p_O_FDREbranch_distanceZ3_),.p_desc34_p_O_FDRE(p_desc34_p_O_FDREbranch_distanceZ3_),.p_desc35_p_O_FDRE(p_desc35_p_O_FDREbranch_distanceZ3_),.p_desc36_p_O_FDRE(p_desc36_p_O_FDREbranch_distanceZ3_),.p_desc37_p_O_FDRE(p_desc37_p_O_FDREbranch_distanceZ3_));
  branch_distanceZ2_inj desc3709(.branch_tdata_2_fast(branch_tdata_2_fast),.buffer_tdata_0(buffer_tdata[0:0]),.buffer_tdata_8(buffer_tdata[8:8]),.buffer_tdata_11(buffer_tdata[11:11]),.buffer_tdata_3(buffer_tdata[3:3]),.buffer_tdata_2(buffer_tdata[2:2]),.buffer_tdata_10(buffer_tdata[10:10]),.buffer_tdata_1(buffer_tdata[1:1]),.buffer_tdata_9(buffer_tdata[9:9]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_0(branch_tdata_2[0:0]),.un10_v_branch_result_axb_0_i_rep2(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep2 ),.un10_v_branch_result_axb_0_i_fast(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_fast ),.un10_v_branch_result_axb_0_i_rep1(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep1 ),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.aclk(aclk),.aresetn_i(aresetn_i),.un1_output_accept(\inst_axi4s_buffer.pr_reg.un1_output_accept ),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.v_branch_result_axb_0_i_fast(\gen_branch_distance.2.inst_branch_distance.v_branch_result.v_branch_result_axb_0_i_fast ),.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ2_),.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ2_),.p_desc39_p_O_FDRE(p_desc39_p_O_FDREbranch_distanceZ2_),.p_desc52_p_O_FDRE(p_desc52_p_O_FDREbranch_distanceZ2_),.p_desc53_p_O_FDRE(p_desc53_p_O_FDREbranch_distanceZ2_),.p_desc54_p_O_FDRE(p_desc54_p_O_FDREbranch_distanceZ2_),.p_desc55_p_O_FDRE(p_desc55_p_O_FDREbranch_distanceZ2_),.p_desc56_p_O_FDRE(p_desc56_p_O_FDREbranch_distanceZ2_));
  branch_distanceZ0_inj desc3710(.branch_tlast(branch_tlast),.branch_tdata_0_fast(branch_tdata_0_fast),.buffer_tdata_11(buffer_tdata[11:11]),.buffer_tdata_3(buffer_tdata[3:3]),.buffer_tdata_2(buffer_tdata[2:2]),.buffer_tdata_10(buffer_tdata[10:10]),.buffer_tdata_1(buffer_tdata[1:1]),.buffer_tdata_9(buffer_tdata[9:9]),.buffer_tdata_0(buffer_tdata[0:0]),.buffer_tdata_8(buffer_tdata[8:8]),.acs_tvalid(acs_tvalid),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_0(branch_tdata_0[0:0]),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.un1_output_accept(\inst_axi4s_buffer.pr_reg.un1_output_accept ),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.buffer_tvalid(buffer_tvalid),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.buffer_tlast(buffer_tlast),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.s_axis_inbranch_tlast_d_RNIIAVE1_O5(s_axis_inbranch_tlast_d_RNIIAVE1_O5),.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ0_),.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ0_),.p_desc63_p_O_FDRE(p_desc63_p_O_FDREbranch_distanceZ0_),.p_desc78_p_O_FDRE(p_desc78_p_O_FDREbranch_distanceZ0_),.p_desc79_p_O_FDRE(p_desc79_p_O_FDREbranch_distanceZ0_),.p_desc80_p_O_FDRE(p_desc80_p_O_FDREbranch_distanceZ0_),.p_desc81_p_O_FDRE(p_desc81_p_O_FDREbranch_distanceZ0_),.p_desc82_p_O_FDRE(p_desc82_p_O_FDREbranch_distanceZ0_));
  branch_distanceZ1_inj desc3711(.branch_tdata_1_fast(branch_tdata_1_fast),.buffer_tdata_0(buffer_tdata[0:0]),.buffer_tdata_8(buffer_tdata[8:8]),.buffer_tdata_11(buffer_tdata[11:11]),.buffer_tdata_3(buffer_tdata[3:3]),.buffer_tdata_1(buffer_tdata[1:1]),.buffer_tdata_9(buffer_tdata[9:9]),.buffer_tdata_2(buffer_tdata[2:2]),.buffer_tdata_10(buffer_tdata[10:10]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_0(branch_tdata_1[0:0]),.v_branch_result_axb_0_i_fast(\gen_branch_distance.2.inst_branch_distance.v_branch_result.v_branch_result_axb_0_i_fast ),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.un10_v_branch_result_axb_0_i_rep2(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep2 ),.aclk(aclk),.aresetn_i(aresetn_i),.un1_output_accept(\inst_axi4s_buffer.pr_reg.un1_output_accept ),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.un10_v_branch_result_axb_0_i_rep1(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_rep1 ),.un10_v_branch_result_axb_0_i_fast(\gen_branch_distance.1.inst_branch_distance.un10_v_branch_result_axb_0_i_fast ),.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ1_),.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDRE(p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ1_),.p_desc83_p_O_FDRE(p_desc83_p_O_FDREbranch_distanceZ1_),.p_desc84_p_O_FDRE(p_desc84_p_O_FDREbranch_distanceZ1_),.p_desc85_p_O_FDRE(p_desc85_p_O_FDREbranch_distanceZ1_),.p_desc86_p_O_FDRE(p_desc86_p_O_FDREbranch_distanceZ1_),.p_desc87_p_O_FDRE(p_desc87_p_O_FDREbranch_distanceZ1_),.p_desc88_p_O_FDRE(p_desc88_p_O_FDREbranch_distanceZ1_));
  acsZ0_inj desc3712(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[57:57]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_50(acs_prob_tdata_50[8:0]),.acs_prob_tdata_51(acs_prob_tdata_51[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_57(acs_prob_tdata_57[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc95_p_O_FD(p_desc95_p_O_FDacsZ0_),.p_desc96_p_O_FD(p_desc96_p_O_FDacsZ0_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_),.p_desc125_p_O_FDRE(p_desc125_p_O_FDREacsZ0_));
  acsZ0_1_inj desc3713(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[12:12]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_25(acs_prob_tdata_25[8:0]),.acs_prob_tdata_24(acs_prob_tdata_24[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_12(acs_prob_tdata_12[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc134_p_O_FD(p_desc134_p_O_FDacsZ0_1_),.p_desc135_p_O_FD(p_desc135_p_O_FDacsZ0_1_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_1_),.p_desc164_p_O_FDRE(p_desc164_p_O_FDREacsZ0_1_));
  acsZ0_2_inj desc3714(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[54:54]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_45(acs_prob_tdata_45[8:0]),.acs_prob_tdata_44(acs_prob_tdata_44[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_54(acs_prob_tdata_54[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc173_p_O_FD(p_desc173_p_O_FDacsZ0_2_),.p_desc174_p_O_FD(p_desc174_p_O_FDacsZ0_2_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_2_),.p_desc203_p_O_FDRE(p_desc203_p_O_FDREacsZ0_2_));
  acsZ0_3_inj desc3715(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[42:42]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_21(acs_prob_tdata_21[8:0]),.acs_prob_tdata_20(acs_prob_tdata_20[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_42(acs_prob_tdata_42[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc212_p_O_FD(p_desc212_p_O_FDacsZ0_3_),.p_desc213_p_O_FD(p_desc213_p_O_FDacsZ0_3_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_3_),.p_desc242_p_O_FDRE(p_desc242_p_O_FDREacsZ0_3_));
  acsZ0_4_inj desc3716(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[24:24]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_49(acs_prob_tdata_49[8:0]),.acs_prob_tdata_48(acs_prob_tdata_48[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_24(acs_prob_tdata_24[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc251_p_O_FD(p_desc251_p_O_FDacsZ0_4_),.p_desc252_p_O_FD(p_desc252_p_O_FDacsZ0_4_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_4_),.p_desc281_p_O_FDRE(p_desc281_p_O_FDREacsZ0_4_));
  acsZ0_5_inj desc3717(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[25:25]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_51(acs_prob_tdata_51[8:0]),.acs_prob_tdata_50(acs_prob_tdata_50[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_25(acs_prob_tdata_25[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc290_p_O_FD(p_desc290_p_O_FDacsZ0_5_),.p_desc291_p_O_FD(p_desc291_p_O_FDacsZ0_5_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_5_),.p_desc320_p_O_FDRE(p_desc320_p_O_FDREacsZ0_5_));
  acsZ0_6_inj desc3718(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[16:16]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_33(acs_prob_tdata_33[8:0]),.acs_prob_tdata_32(acs_prob_tdata_32[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_16(acs_prob_tdata_16[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc329_p_O_FD(p_desc329_p_O_FDacsZ0_6_),.p_desc330_p_O_FD(p_desc330_p_O_FDacsZ0_6_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_6_),.p_desc359_p_O_FDRE(p_desc359_p_O_FDREacsZ0_6_));
  acsZ0_7_inj desc3719(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[1:1]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_3(acs_prob_tdata_3[8:0]),.acs_prob_tdata_2(acs_prob_tdata_2[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:0]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_1(acs_prob_tdata_1[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc368_p_O_FD(p_desc368_p_O_FDacsZ0_7_),.p_desc369_p_O_FD(p_desc369_p_O_FDacsZ0_7_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_7_),.p_desc398_p_O_FDRE(p_desc398_p_O_FDREacsZ0_7_));
  acsZ0_8_inj desc3720(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[33:33]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_3(acs_prob_tdata_3[8:0]),.acs_prob_tdata_2(acs_prob_tdata_2[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_33(acs_prob_tdata_33[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc407_p_O_FD(p_desc407_p_O_FDacsZ0_8_),.p_desc408_p_O_FD(p_desc408_p_O_FDacsZ0_8_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_8_),.p_desc437_p_O_FDRE(p_desc437_p_O_FDREacsZ0_8_));
  acsZ0_9_inj desc3721(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[18:18]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_37(acs_prob_tdata_37[8:0]),.acs_prob_tdata_36(acs_prob_tdata_36[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_18(acs_prob_tdata_18[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc446_p_O_FD(p_desc446_p_O_FDacsZ0_9_),.p_desc447_p_O_FD(p_desc447_p_O_FDacsZ0_9_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_9_),.p_desc476_p_O_FDRE(p_desc476_p_O_FDREacsZ0_9_));
  acsZ0_10_inj desc3722(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[3:3]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_7(acs_prob_tdata_7[8:0]),.acs_prob_tdata_6(acs_prob_tdata_6[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:0]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_3(acs_prob_tdata_3[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc485_p_O_FD(p_desc485_p_O_FDacsZ0_10_),.p_desc486_p_O_FD(p_desc486_p_O_FDacsZ0_10_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_10_),.p_desc515_p_O_FDRE(p_desc515_p_O_FDREacsZ0_10_));
  acsZ0_11_inj desc3723(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[62:62]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_61(acs_prob_tdata_61[8:0]),.acs_prob_tdata_60(acs_prob_tdata_60[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_62(acs_prob_tdata_62[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc524_p_O_FD(p_desc524_p_O_FDacsZ0_11_),.p_desc525_p_O_FD(p_desc525_p_O_FDacsZ0_11_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_11_),.p_desc554_p_O_FDRE(p_desc554_p_O_FDREacsZ0_11_));
  acsZ0_12_inj desc3724(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[47:47]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_31(acs_prob_tdata_31[8:0]),.acs_prob_tdata_30(acs_prob_tdata_30[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_47(acs_prob_tdata_47[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc563_p_O_FD(p_desc563_p_O_FDacsZ0_12_),.p_desc564_p_O_FD(p_desc564_p_O_FDacsZ0_12_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_12_),.p_desc593_p_O_FDRE(p_desc593_p_O_FDREacsZ0_12_));
  acsZ0_13_inj desc3725(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[5:5]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_11(acs_prob_tdata_11[8:0]),.acs_prob_tdata_10(acs_prob_tdata_10[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_5(acs_prob_tdata_5[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc602_p_O_FD(p_desc602_p_O_FDacsZ0_13_),.p_desc603_p_O_FD(p_desc603_p_O_FDacsZ0_13_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_13_),.p_desc632_p_O_FDRE(p_desc632_p_O_FDREacsZ0_13_));
  acsZ0_14_inj desc3726(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[37:37]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_11(acs_prob_tdata_11[8:0]),.acs_prob_tdata_10(acs_prob_tdata_10[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_37(acs_prob_tdata_37[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc641_p_O_FD(p_desc641_p_O_FDacsZ0_14_),.p_desc642_p_O_FD(p_desc642_p_O_FDacsZ0_14_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_14_),.p_desc671_p_O_FDRE(p_desc671_p_O_FDREacsZ0_14_));
  acsZ0_15_inj desc3727(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[49:49]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_34(acs_prob_tdata_34[8:0]),.acs_prob_tdata_35(acs_prob_tdata_35[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_49(acs_prob_tdata_49[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc680_p_O_FD(p_desc680_p_O_FDacsZ0_15_),.p_desc681_p_O_FD(p_desc681_p_O_FDacsZ0_15_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_15_),.p_desc710_p_O_FDRE(p_desc710_p_O_FDREacsZ0_15_));
  acsZ0_16_inj desc3728(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[34:34]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_5(acs_prob_tdata_5[8:0]),.acs_prob_tdata_4(acs_prob_tdata_4[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_34(acs_prob_tdata_34[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc719_p_O_FD(p_desc719_p_O_FDacsZ0_16_),.p_desc720_p_O_FD(p_desc720_p_O_FDacsZ0_16_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_16_),.p_desc749_p_O_FDRE(p_desc749_p_O_FDREacsZ0_16_));
  acsZ0_17_inj desc3729(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[19:19]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_39(acs_prob_tdata_39[8:0]),.acs_prob_tdata_38(acs_prob_tdata_38[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_19(acs_prob_tdata_19[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc758_p_O_FD(p_desc758_p_O_FDacsZ0_17_),.p_desc759_p_O_FD(p_desc759_p_O_FDacsZ0_17_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_17_),.p_desc788_p_O_FDRE(p_desc788_p_O_FDREacsZ0_17_));
  acsZ0_18_inj desc3730(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[4:4]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_9(acs_prob_tdata_9[8:0]),.acs_prob_tdata_8(acs_prob_tdata_8[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:0]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_4(acs_prob_tdata_4[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc797_p_O_FD(p_desc797_p_O_FDacsZ0_18_),.p_desc798_p_O_FD(p_desc798_p_O_FDacsZ0_18_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_18_),.p_desc827_p_O_FDRE(p_desc827_p_O_FDREacsZ0_18_));
  acsZ0_19_inj desc3731(.branch_tvalid(branch_tvalid),.acs_prob_tdata_63(acs_prob_tdata_63[8:0]),.acs_dec_tdata(acs_dec_tdata[63:63]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_62(acs_prob_tdata_62[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tlast(branch_tlast),.branch_tdata_0_fast(branch_tdata_0_fast),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_19_));
  acsZ0_20_inj desc3732(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[61:61]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_59(acs_prob_tdata_59[8:0]),.acs_prob_tdata_58(acs_prob_tdata_58[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_61(acs_prob_tdata_61[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc873_p_O_FD(p_desc873_p_O_FDacsZ0_20_),.p_desc874_p_O_FD(p_desc874_p_O_FDacsZ0_20_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_20_),.p_desc903_p_O_FDRE(p_desc903_p_O_FDREacsZ0_20_));
  acsZ0_21_inj desc3733(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[32:32]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_1(acs_prob_tdata_1[8:0]),.acs_prob_tdata_0(acs_prob_tdata_0[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_32(acs_prob_tdata_32[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc912_p_O_FD(p_desc912_p_O_FDacsZ0_21_),.p_desc913_p_O_FD(p_desc913_p_O_FDacsZ0_21_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_21_),.p_desc942_p_O_FDRE(p_desc942_p_O_FDREacsZ0_21_));
  acsZ1_inj desc3734(.acs_tvalid(acs_tvalid),.branch_tlast(branch_tlast),.branch_tvalid(branch_tvalid),.acs_prob_tdata_0(acs_prob_tdata_0[8:0]),.acs_dec_tdata(acs_dec_tdata[0:0]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_1(acs_prob_tdata_1[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_tlast(acs_tlast),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.un1_output_accept(\inst_axi4s_buffer.pr_reg.un1_output_accept ),.s_axis_inbranch_tlast_d_RNIIAVE1_O5(s_axis_inbranch_tlast_d_RNIIAVE1_O5),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.un1_s_axis_input_tvalid(\inst_ram_ctrl.pr_write_ram.un1_s_axis_input_tvalid ),.aresetn(aresetn));
  acsZ0_22_inj desc3735(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[46:46]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_29(acs_prob_tdata_29[8:0]),.acs_prob_tdata_28(acs_prob_tdata_28[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_46(acs_prob_tdata_46[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc989_p_O_FD(p_desc989_p_O_FDacsZ0_22_),.p_desc990_p_O_FD(p_desc990_p_O_FDacsZ0_22_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_22_),.p_desc1019_p_O_FDRE(p_desc1019_p_O_FDREacsZ0_22_));
  acsZ0_23_inj desc3736(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[9:9]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_19(acs_prob_tdata_19[8:0]),.acs_prob_tdata_18(acs_prob_tdata_18[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_9(acs_prob_tdata_9[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1028_p_O_FD(p_desc1028_p_O_FDacsZ0_23_),.p_desc1029_p_O_FD(p_desc1029_p_O_FDacsZ0_23_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_23_),.p_desc1058_p_O_FDRE(p_desc1058_p_O_FDREacsZ0_23_));
  acsZ0_24_inj desc3737(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[2:2]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_5(acs_prob_tdata_5[8:0]),.acs_prob_tdata_4(acs_prob_tdata_4[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:0]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_2(acs_prob_tdata_2[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1067_p_O_FD(p_desc1067_p_O_FDacsZ0_24_),.p_desc1068_p_O_FD(p_desc1068_p_O_FDacsZ0_24_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_24_),.p_desc1097_p_O_FDRE(p_desc1097_p_O_FDREacsZ0_24_));
  acsZ0_25_inj desc3738(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[52:52]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_41(acs_prob_tdata_41[8:0]),.acs_prob_tdata_40(acs_prob_tdata_40[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_52(acs_prob_tdata_52[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1106_p_O_FD(p_desc1106_p_O_FDacsZ0_25_),.p_desc1107_p_O_FD(p_desc1107_p_O_FDacsZ0_25_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_25_),.p_desc1136_p_O_FDRE(p_desc1136_p_O_FDREacsZ0_25_));
  acsZ0_26_inj desc3739(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[10:10]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_21(acs_prob_tdata_21[8:0]),.acs_prob_tdata_20(acs_prob_tdata_20[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_10(acs_prob_tdata_10[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1145_p_O_FD(p_desc1145_p_O_FDacsZ0_26_),.p_desc1146_p_O_FD(p_desc1146_p_O_FDacsZ0_26_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_26_),.p_desc1175_p_O_FDRE(p_desc1175_p_O_FDREacsZ0_26_));
  acsZ0_27_inj desc3740(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[22:22]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_45(acs_prob_tdata_45[8:0]),.acs_prob_tdata_44(acs_prob_tdata_44[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_22(acs_prob_tdata_22[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1184_p_O_FD(p_desc1184_p_O_FDacsZ0_27_),.p_desc1185_p_O_FD(p_desc1185_p_O_FDacsZ0_27_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_27_),.p_desc1214_p_O_FDRE(p_desc1214_p_O_FDREacsZ0_27_));
  acsZ0_28_inj desc3741(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[7:7]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_15(acs_prob_tdata_15[8:0]),.acs_prob_tdata_14(acs_prob_tdata_14[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_7(acs_prob_tdata_7[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1223_p_O_FD(p_desc1223_p_O_FDacsZ0_28_),.p_desc1224_p_O_FD(p_desc1224_p_O_FDacsZ0_28_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_28_),.p_desc1253_p_O_FDRE(p_desc1253_p_O_FDREacsZ0_28_));
  acsZ0_29_inj desc3742(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[39:39]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_15(acs_prob_tdata_15[8:0]),.acs_prob_tdata_14(acs_prob_tdata_14[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_39(acs_prob_tdata_39[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1262_p_O_FD(p_desc1262_p_O_FDacsZ0_29_),.p_desc1263_p_O_FD(p_desc1263_p_O_FDacsZ0_29_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_29_),.p_desc1292_p_O_FDRE(p_desc1292_p_O_FDREacsZ0_29_));
  acsZ0_30_inj desc3743(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[51:51]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_39(acs_prob_tdata_39[8:0]),.acs_prob_tdata_38(acs_prob_tdata_38[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_51(acs_prob_tdata_51[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1301_p_O_FD(p_desc1301_p_O_FDacsZ0_30_),.p_desc1302_p_O_FD(p_desc1302_p_O_FDacsZ0_30_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_30_),.p_desc1331_p_O_FDRE(p_desc1331_p_O_FDREacsZ0_30_));
  acsZ0_31_inj desc3744(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[36:36]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_9(acs_prob_tdata_9[8:0]),.acs_prob_tdata_8(acs_prob_tdata_8[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_36(acs_prob_tdata_36[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1340_p_O_FD(p_desc1340_p_O_FDacsZ0_31_),.p_desc1341_p_O_FD(p_desc1341_p_O_FDacsZ0_31_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_31_),.p_desc1370_p_O_FDRE(p_desc1370_p_O_FDREacsZ0_31_));
  acsZ0_32_inj desc3745(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[21:21]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_43(acs_prob_tdata_43[8:0]),.acs_prob_tdata_42(acs_prob_tdata_42[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_21(acs_prob_tdata_21[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1379_p_O_FD(p_desc1379_p_O_FDacsZ0_32_),.p_desc1380_p_O_FD(p_desc1380_p_O_FDacsZ0_32_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_32_),.p_desc1409_p_O_FDRE(p_desc1409_p_O_FDREacsZ0_32_));
  acsZ0_33_inj desc3746(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[53:53]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_43(acs_prob_tdata_43[8:0]),.acs_prob_tdata_42(acs_prob_tdata_42[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_53(acs_prob_tdata_53[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1418_p_O_FD(p_desc1418_p_O_FDacsZ0_33_),.p_desc1419_p_O_FD(p_desc1419_p_O_FDacsZ0_33_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_33_),.p_desc1448_p_O_FDRE(p_desc1448_p_O_FDREacsZ0_33_));
  acsZ0_34_inj desc3747(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[11:11]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_23(acs_prob_tdata_23[8:0]),.acs_prob_tdata_22(acs_prob_tdata_22[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_11(acs_prob_tdata_11[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1457_p_O_FD(p_desc1457_p_O_FDacsZ0_34_),.p_desc1458_p_O_FD(p_desc1458_p_O_FDacsZ0_34_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_34_),.p_desc1487_p_O_FDRE(p_desc1487_p_O_FDREacsZ0_34_));
  acsZ0_35_inj desc3748(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[23:23]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_47(acs_prob_tdata_47[8:0]),.acs_prob_tdata_46(acs_prob_tdata_46[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_23(acs_prob_tdata_23[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1496_p_O_FD(p_desc1496_p_O_FDacsZ0_35_),.p_desc1497_p_O_FD(p_desc1497_p_O_FDacsZ0_35_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_35_),.p_desc1526_p_O_FDRE(p_desc1526_p_O_FDREacsZ0_35_));
  acsZ0_36_inj desc3749(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[8:8]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_16(acs_prob_tdata_16[8:0]),.acs_prob_tdata_17(acs_prob_tdata_17[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_8(acs_prob_tdata_8[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1535_p_O_FD(p_desc1535_p_O_FDacsZ0_36_),.p_desc1536_p_O_FD(p_desc1536_p_O_FDacsZ0_36_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_36_),.p_desc1565_p_O_FDRE(p_desc1565_p_O_FDREacsZ0_36_));
  acsZ0_37_inj desc3750(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[40:40]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_17(acs_prob_tdata_17[8:0]),.acs_prob_tdata_16(acs_prob_tdata_16[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_40(acs_prob_tdata_40[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1574_p_O_FD(p_desc1574_p_O_FDacsZ0_37_),.p_desc1575_p_O_FD(p_desc1575_p_O_FDacsZ0_37_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_37_),.p_desc1604_p_O_FDRE(p_desc1604_p_O_FDREacsZ0_37_));
  acsZ0_38_inj desc3751(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[17:17]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_35(acs_prob_tdata_35[8:0]),.acs_prob_tdata_34(acs_prob_tdata_34[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_17(acs_prob_tdata_17[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1613_p_O_FD(p_desc1613_p_O_FDacsZ0_38_),.p_desc1614_p_O_FD(p_desc1614_p_O_FDacsZ0_38_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_38_),.p_desc1643_p_O_FDRE(p_desc1643_p_O_FDREacsZ0_38_));
  acsZ0_39_inj desc3752(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[50:50]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_37(acs_prob_tdata_37[8:0]),.acs_prob_tdata_36(acs_prob_tdata_36[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_50(acs_prob_tdata_50[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1652_p_O_FD(p_desc1652_p_O_FDacsZ0_39_),.p_desc1653_p_O_FD(p_desc1653_p_O_FDacsZ0_39_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_39_),.p_desc1682_p_O_FDRE(p_desc1682_p_O_FDREacsZ0_39_));
  acsZ0_40_inj desc3753(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[35:35]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_7(acs_prob_tdata_7[8:0]),.acs_prob_tdata_6(acs_prob_tdata_6[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_35(acs_prob_tdata_35[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1691_p_O_FD(p_desc1691_p_O_FDacsZ0_40_),.p_desc1692_p_O_FD(p_desc1692_p_O_FDacsZ0_40_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_40_),.p_desc1721_p_O_FDRE(p_desc1721_p_O_FDREacsZ0_40_));
  acsZ0_41_inj desc3754(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[6:6]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_13(acs_prob_tdata_13[8:0]),.acs_prob_tdata_12(acs_prob_tdata_12[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_6(acs_prob_tdata_6[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1730_p_O_FD(p_desc1730_p_O_FDacsZ0_41_),.p_desc1731_p_O_FD(p_desc1731_p_O_FDacsZ0_41_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_41_),.p_desc1760_p_O_FDRE(p_desc1760_p_O_FDREacsZ0_41_));
  acsZ0_42_inj desc3755(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[48:48]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_33(acs_prob_tdata_33[8:0]),.acs_prob_tdata_32(acs_prob_tdata_32[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_48(acs_prob_tdata_48[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1769_p_O_FD(p_desc1769_p_O_FDacsZ0_42_),.p_desc1770_p_O_FD(p_desc1770_p_O_FDacsZ0_42_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_42_),.p_desc1799_p_O_FDRE(p_desc1799_p_O_FDREacsZ0_42_));
  acsZ0_43_inj desc3756(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[20:20]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_41(acs_prob_tdata_41[8:0]),.acs_prob_tdata_40(acs_prob_tdata_40[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_20(acs_prob_tdata_20[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1808_p_O_FD(p_desc1808_p_O_FDacsZ0_43_),.p_desc1809_p_O_FD(p_desc1809_p_O_FDacsZ0_43_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_43_),.p_desc1838_p_O_FDRE(p_desc1838_p_O_FDREacsZ0_43_));
  acsZ0_44_inj desc3757(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[38:38]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_13(acs_prob_tdata_13[8:0]),.acs_prob_tdata_12(acs_prob_tdata_12[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_38(acs_prob_tdata_38[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1847_p_O_FD(p_desc1847_p_O_FDacsZ0_44_),.p_desc1848_p_O_FD(p_desc1848_p_O_FDacsZ0_44_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_44_),.p_desc1877_p_O_FDRE(p_desc1877_p_O_FDREacsZ0_44_));
  acsZ0_45_inj desc3758(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[41:41]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_19(acs_prob_tdata_19[8:0]),.acs_prob_tdata_18(acs_prob_tdata_18[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_41(acs_prob_tdata_41[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1886_p_O_FD(p_desc1886_p_O_FDacsZ0_45_),.p_desc1887_p_O_FD(p_desc1887_p_O_FDacsZ0_45_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_45_),.p_desc1916_p_O_FDRE(p_desc1916_p_O_FDREacsZ0_45_));
  acsZ0_46_inj desc3759(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[26:26]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_53(acs_prob_tdata_53[8:0]),.acs_prob_tdata_52(acs_prob_tdata_52[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_26(acs_prob_tdata_26[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1925_p_O_FD(p_desc1925_p_O_FDacsZ0_46_),.p_desc1926_p_O_FD(p_desc1926_p_O_FDacsZ0_46_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_46_),.p_desc1955_p_O_FDRE(p_desc1955_p_O_FDREacsZ0_46_));
  acsZ0_47_inj desc3760(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[58:58]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_53(acs_prob_tdata_53[8:0]),.acs_prob_tdata_52(acs_prob_tdata_52[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_58(acs_prob_tdata_58[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc1964_p_O_FD(p_desc1964_p_O_FDacsZ0_47_),.p_desc1965_p_O_FD(p_desc1965_p_O_FDacsZ0_47_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_47_),.p_desc1994_p_O_FDRE(p_desc1994_p_O_FDREacsZ0_47_));
  acsZ0_48_inj desc3761(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[43:43]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_23(acs_prob_tdata_23[8:0]),.acs_prob_tdata_22(acs_prob_tdata_22[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_43(acs_prob_tdata_43[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2003_p_O_FD(p_desc2003_p_O_FDacsZ0_48_),.p_desc2004_p_O_FD(p_desc2004_p_O_FDacsZ0_48_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_48_),.p_desc2033_p_O_FDRE(p_desc2033_p_O_FDREacsZ0_48_));
  acsZ0_49_inj desc3762(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[55:55]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_47(acs_prob_tdata_47[8:0]),.acs_prob_tdata_46(acs_prob_tdata_46[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_55(acs_prob_tdata_55[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2042_p_O_FD(p_desc2042_p_O_FDacsZ0_49_),.p_desc2043_p_O_FD(p_desc2043_p_O_FDacsZ0_49_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_49_),.p_desc2072_p_O_FDRE(p_desc2072_p_O_FDREacsZ0_49_));
  acsZ0_50_inj desc3763(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[13:13]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_27(acs_prob_tdata_27[8:0]),.acs_prob_tdata_26(acs_prob_tdata_26[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_13(acs_prob_tdata_13[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2081_p_O_FD(p_desc2081_p_O_FDacsZ0_50_),.p_desc2082_p_O_FD(p_desc2082_p_O_FDacsZ0_50_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_50_),.p_desc2111_p_O_FDRE(p_desc2111_p_O_FDREacsZ0_50_));
  acsZ0_51_inj desc3764(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[45:45]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_26(acs_prob_tdata_26[8:0]),.acs_prob_tdata_27(acs_prob_tdata_27[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_45(acs_prob_tdata_45[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2120_p_O_FD(p_desc2120_p_O_FDacsZ0_51_),.p_desc2121_p_O_FD(p_desc2121_p_O_FDacsZ0_51_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_51_),.p_desc2150_p_O_FDRE(p_desc2150_p_O_FDREacsZ0_51_));
  acsZ0_52_inj desc3765(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[30:30]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_61(acs_prob_tdata_61[8:0]),.acs_prob_tdata_60(acs_prob_tdata_60[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_30(acs_prob_tdata_30[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2159_p_O_FD(p_desc2159_p_O_FDacsZ0_52_),.p_desc2160_p_O_FD(p_desc2160_p_O_FDacsZ0_52_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_52_),.p_desc2189_p_O_FDRE(p_desc2189_p_O_FDREacsZ0_52_));
  acsZ0_53_inj desc3766(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[15:15]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_31(acs_prob_tdata_31[8:0]),.acs_prob_tdata_30(acs_prob_tdata_30[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_15(acs_prob_tdata_15[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2198_p_O_FD(p_desc2198_p_O_FDacsZ0_53_),.p_desc2199_p_O_FD(p_desc2199_p_O_FDacsZ0_53_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_53_),.p_desc2228_p_O_FDRE(p_desc2228_p_O_FDREacsZ0_53_));
  acsZ0_54_inj desc3767(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[27:27]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_55(acs_prob_tdata_55[8:0]),.acs_prob_tdata_54(acs_prob_tdata_54[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_27(acs_prob_tdata_27[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2237_p_O_FD(p_desc2237_p_O_FDacsZ0_54_),.p_desc2238_p_O_FD(p_desc2238_p_O_FDacsZ0_54_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_54_),.p_desc2267_p_O_FDRE(p_desc2267_p_O_FDREacsZ0_54_));
  acsZ0_55_inj desc3768(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[59:59]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_55(acs_prob_tdata_55[8:0]),.acs_prob_tdata_54(acs_prob_tdata_54[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_59(acs_prob_tdata_59[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2276_p_O_FD(p_desc2276_p_O_FDacsZ0_55_),.p_desc2277_p_O_FD(p_desc2277_p_O_FDacsZ0_55_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_55_),.p_desc2306_p_O_FDRE(p_desc2306_p_O_FDREacsZ0_55_));
  acsZ0_56_inj desc3769(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[44:44]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_25(acs_prob_tdata_25[8:0]),.acs_prob_tdata_24(acs_prob_tdata_24[8:0]),.write_ram_fsm_3(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_44(acs_prob_tdata_44[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2315_p_O_FD(p_desc2315_p_O_FDacsZ0_56_),.p_desc2316_p_O_FD(p_desc2316_p_O_FDacsZ0_56_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_56_),.p_desc2345_p_O_FDRE(p_desc2345_p_O_FDREacsZ0_56_));
  acsZ0_57_inj desc3770(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[56:56]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_49(acs_prob_tdata_49[8:0]),.acs_prob_tdata_48(acs_prob_tdata_48[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_56(acs_prob_tdata_56[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2354_p_O_FD(p_desc2354_p_O_FDacsZ0_57_),.p_desc2355_p_O_FD(p_desc2355_p_O_FDacsZ0_57_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_57_),.p_desc2384_p_O_FDRE(p_desc2384_p_O_FDREacsZ0_57_));
  acsZ0_58_inj desc3771(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[14:14]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_29(acs_prob_tdata_29[8:0]),.acs_prob_tdata_28(acs_prob_tdata_28[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_0_fast(branch_tdata_0_fast),.acs_prob_tdata_14(acs_prob_tdata_14[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_3_0_rep1(branch_tdata_3_0_rep1),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2393_p_O_FD(p_desc2393_p_O_FDacsZ0_58_),.p_desc2394_p_O_FD(p_desc2394_p_O_FDacsZ0_58_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_58_),.p_desc2423_p_O_FDRE(p_desc2423_p_O_FDREacsZ0_58_));
  acsZ0_59_inj desc3772(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[31:31]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_63(acs_prob_tdata_63[8:0]),.acs_prob_tdata_62(acs_prob_tdata_62[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_31(acs_prob_tdata_31[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2432_p_O_FD(p_desc2432_p_O_FDacsZ0_59_),.p_desc2433_p_O_FD(p_desc2433_p_O_FDacsZ0_59_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_59_),.p_desc2462_p_O_FDRE(p_desc2462_p_O_FDREacsZ0_59_));
  acsZ0_60_inj desc3773(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[28:28]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_57(acs_prob_tdata_57[8:0]),.acs_prob_tdata_56(acs_prob_tdata_56[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_2_fast(branch_tdata_2_fast),.acs_prob_tdata_28(acs_prob_tdata_28[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_1_0_rep1(branch_tdata_1_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2471_p_O_FD(p_desc2471_p_O_FDacsZ0_60_),.p_desc2472_p_O_FD(p_desc2472_p_O_FDacsZ0_60_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_60_),.p_desc2501_p_O_FDRE(p_desc2501_p_O_FDREacsZ0_60_));
  acsZ0_61_inj desc3774(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[29:29]),.branch_tdata_0_1(branch_tdata_0[1:1]),.branch_tdata_0_2(branch_tdata_0[2:2]),.branch_tdata_0_3(branch_tdata_0[3:3]),.branch_tdata_0_5(branch_tdata_0[5:5]),.branch_tdata_0_0(branch_tdata_0[0:0]),.branch_tdata_3(branch_tdata_3[5:0]),.acs_prob_tdata_59(acs_prob_tdata_59[8:0]),.acs_prob_tdata_58(acs_prob_tdata_58[8:0]),.write_ram_fsm(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_3_fast(branch_tdata_3_fast),.acs_prob_tdata_29(acs_prob_tdata_29[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_0_0_rep2(branch_tdata_0_0_rep2),.branch_tdata_3_0_rep2(branch_tdata_3_0_rep2),.branch_tdata_0_0_rep1(branch_tdata_0_0_rep1),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2510_p_O_FD(p_desc2510_p_O_FDacsZ0_61_),.p_desc2511_p_O_FD(p_desc2511_p_O_FDacsZ0_61_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_61_),.p_desc2540_p_O_FDRE(p_desc2540_p_O_FDREacsZ0_61_));
  acsZ0_62_inj desc3775(.branch_tlast(branch_tlast),.acs_dec_tdata(acs_dec_tdata[60:60]),.branch_tdata_1_1(branch_tdata_1[1:1]),.branch_tdata_1_2(branch_tdata_1[2:2]),.branch_tdata_1_3(branch_tdata_1[3:3]),.branch_tdata_1_5(branch_tdata_1[5:5]),.branch_tdata_1_0(branch_tdata_1[0:0]),.branch_tdata_2_1(branch_tdata_2[1:1]),.branch_tdata_2_2(branch_tdata_2[2:2]),.branch_tdata_2_3(branch_tdata_2[3:3]),.branch_tdata_2_5(branch_tdata_2[5:5]),.branch_tdata_2_0(branch_tdata_2[0:0]),.acs_prob_tdata_57(acs_prob_tdata_57[8:0]),.acs_prob_tdata_56(acs_prob_tdata_56[8:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.branch_tvalid(branch_tvalid),.branch_tdata_1_fast(branch_tdata_1_fast),.acs_prob_tdata_60(acs_prob_tdata_60[8:0]),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ),.aclk(aclk),.aresetn_i(aresetn_i),.branch_tdata_1_0_rep2(branch_tdata_1_0_rep2),.branch_tdata_2_0_rep2(branch_tdata_2_0_rep2),.branch_tdata_2_0_rep1(branch_tdata_2_0_rep1),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.aresetn(aresetn),.p_desc2549_p_O_FD(p_desc2549_p_O_FDacsZ0_62_),.p_desc2550_p_O_FD(p_desc2550_p_O_FDacsZ0_62_),.p_m_axis_outdec_tdata_Z_p_O_FDRE(p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_62_),.p_desc2579_p_O_FDRE(p_desc2579_p_O_FDREacsZ0_62_));
  ram_ctrl_inj inst_ram_ctrl(.acs_tlast(acs_tlast),.acs_tvalid(acs_tvalid),.write_ram_fsm_1(\inst_ram_ctrl.write_ram_fsm [1:1]),.write_ram_fsm_0(\inst_ram_ctrl.write_ram_fsm [0:0]),.write_ram_fsm_4(\inst_ram_ctrl.write_ram_fsm [4:4]),.ram_tlast(ram_tlast[1:0]),.ram_last_tuser(ram_last_tuser[1:0]),.s_axis_ctrl_tdata_16(s_axis_ctrl_tdata[16:16]),.s_axis_ctrl_tdata_17(s_axis_ctrl_tdata[17:17]),.s_axis_ctrl_tdata_18(s_axis_ctrl_tdata[18:18]),.s_axis_ctrl_tdata_19(s_axis_ctrl_tdata[19:19]),.s_axis_ctrl_tdata_20(s_axis_ctrl_tdata[20:20]),.s_axis_ctrl_tdata_21(s_axis_ctrl_tdata[21:21]),.s_axis_ctrl_tdata_22(s_axis_ctrl_tdata[22:22]),.s_axis_ctrl_tdata_0(s_axis_ctrl_tdata[0:0]),.s_axis_ctrl_tdata_1(s_axis_ctrl_tdata[1:1]),.s_axis_ctrl_tdata_2(s_axis_ctrl_tdata[2:2]),.s_axis_ctrl_tdata_3(s_axis_ctrl_tdata[3:3]),.s_axis_ctrl_tdata_4(s_axis_ctrl_tdata[4:4]),.s_axis_ctrl_tdata_5(s_axis_ctrl_tdata[5:5]),.s_axis_ctrl_tdata_6(s_axis_ctrl_tdata[6:6]),.ram_buffer_full(\inst_ram_ctrl.ram_buffer_full [1:0]),.traceback_tvalid(traceback_tvalid[1:0]),.ram_tvalid(ram_tvalid[1:0]),.ram_buffer_1_1(\inst_ram_ctrl.pr_buf_ram_output.1.ram_buffer_1_1 [63:0]),.ram_buffer_0_2(\inst_ram_ctrl.pr_buf_ram_output.0.ram_buffer_0_2 [63:0]),.ram_window_tuser(ram_window_tuser[1:0]),.reorder_tvalid_fast(reorder_tvalid_fast[1:0]),.ram_buffer_0(\inst_ram_ctrl.ram_buffer_0 [63:0]),.ram_buffer_1(\inst_ram_ctrl.ram_buffer_1 [63:0]),.acs_dec_tdata(acs_dec_tdata[63:0]),.aresetn(aresetn),.reorder_tvalid_1_rep1(reorder_tvalid_1_rep1),.un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5(\pr_buf_ram_output.1.un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ),.un1_s_axis_input_tvalid(\inst_ram_ctrl.pr_write_ram.un1_s_axis_input_tvalid ),.aclk(aclk),.write_ram_fsm_0_rep1(\inst_ram_ctrl.write_ram_fsm_0_rep1 ),.write_ram_fsm_0_rep2(\inst_ram_ctrl.write_ram_fsm_0_rep2 ),.write_ram_fsm_4_rep1(\inst_ram_ctrl.write_ram_fsm_4_rep1 ),.write_ram_fsm_4_rep2(\inst_ram_ctrl.write_ram_fsm_4_rep2 ),.aresetn_i(aresetn_i),.N_1756_1(\inst_ram_ctrl.N_1756_1 ),.reorder_tvalid_0_rep1(reorder_tvalid_0_rep1),.reorder_tvalid_0_rep2(reorder_tvalid_0_rep2),.N_99(N_99),.s_axis_ctrl_tvalid(s_axis_ctrl_tvalid),.s_axis_ctrl_tready(s_axis_ctrl_tready),.un27_s_axis_input_tready_int(\inst_ram_ctrl.un27_s_axis_input_tready_int ));
  trellis_traceback_inj desc3776(.ram_window_tuser(ram_window_tuser[0:0]),.ram_tvalid(ram_tvalid[0:0]),.traceback_tvalid(traceback_tvalid[0:0]),.traceback_tdata(traceback_tdata[0:0]),.buffer_cnt(\gen_inst_reorder.0.inst_reorder.buffer_cnt [2:0]),.ram_last_tuser(ram_last_tuser[0:0]),.buffer_cnt_0(\gen_inst_reorder.1.inst_reorder.buffer_cnt [2:0]),.ram_buffer_full(\inst_ram_ctrl.ram_buffer_full [0:0]),.ram_buffer_0(\inst_ram_ctrl.ram_buffer_0 [63:0]),.ram_buffer_0_2(\inst_ram_ctrl.pr_buf_ram_output.0.ram_buffer_0_2 [63:0]),.traceback_last_tuser(traceback_last_tuser[0:0]),.traceback_tlast(traceback_tlast[0:0]),.ram_tlast(ram_tlast[0:0]),.reorder_tvalid_0_rep1(reorder_tvalid_0_rep1),.reorder_tvalid_0_rep2(reorder_tvalid_0_rep2),.aclk(aclk),.aresetn_i(aresetn_i),.N_129(N_129),.last_window(\gen_inst_reorder.0.inst_reorder.last_window ),.aresetn(aresetn),.N_130(N_130),.last_window_0(\gen_inst_reorder.1.inst_reorder.last_window ),.m_axis_output_tlast(m_axis_output_tlast));
  trellis_traceback_1_inj desc3777(.traceback_last_tuser(traceback_last_tuser[1:1]),.ram_tvalid(ram_tvalid[1:1]),.traceback_tvalid(traceback_tvalid[1:1]),.traceback_tdata(traceback_tdata[1:1]),.ram_last_tuser(ram_last_tuser[1:1]),.ram_window_tuser(ram_window_tuser[1:1]),.ram_buffer_full(\inst_ram_ctrl.ram_buffer_full [1:1]),.ram_buffer_1(\inst_ram_ctrl.ram_buffer_1 [63:0]),.ram_buffer_1_1(\inst_ram_ctrl.pr_buf_ram_output.1.ram_buffer_1_1 [63:0]),.traceback_tlast(traceback_tlast[1:1]),.ram_tlast(ram_tlast[1:1]),.reorder_tvalid_1_rep1(reorder_tvalid_1_rep1),.N_104(N_104),.send_output_rep1(\gen_inst_reorder.1.inst_reorder.send_output_rep1 ),.aclk(aclk),.aresetn_i(aresetn_i),.aresetn(aresetn),.un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5(\pr_buf_ram_output.1.un21_m_axis_output_tvalid_int_0_a2_lut6_2_O5 ));
  reorder_inj desc3778(.traceback_last_tuser(traceback_last_tuser[1:1]),.traceback_tvalid(traceback_tvalid[1:1]),.reorder_tvalid_fast(reorder_tvalid_fast[1:1]),.reorder_tvalid_0(reorder_tvalid),.traceback_tlast(traceback_tlast[1:1]),.current_active(current_active),.reorder_last_tuser(reorder_last_tuser[1:1]),.buffer_cnt_1(\gen_inst_reorder.1.inst_reorder.buffer_cnt [1:1]),.buffer_cnt_2(\gen_inst_reorder.1.inst_reorder.buffer_cnt [2:2]),.buffer_cnt_0(\gen_inst_reorder.1.inst_reorder.buffer_cnt [0:0]),.reorder_tdata_0(reorder_tdata),.traceback_tdata(traceback_tdata[1:1]),.N_104(N_104),.m_axis_output_tvalid(m_axis_output_tvalid),.aresetn(aresetn),.reorder_tvalid_1_rep1(reorder_tvalid_1_rep1),.m_axis_output_tready(m_axis_output_tready),.aclk(aclk),.aresetn_i(aresetn_i),.last_window(\gen_inst_reorder.1.inst_reorder.last_window ),.send_output_rep1(\gen_inst_reorder.1.inst_reorder.send_output_rep1 ),.m_axis_output_tdata(m_axis_output_tdata),.N_130(N_130));
  reorder_1_inj desc3779(.traceback_last_tuser(traceback_last_tuser[0:0]),.traceback_tvalid(traceback_tvalid[0:0]),.reorder_tvalid_fast(reorder_tvalid_fast[0:0]),.reorder_tvalid(reorder_tvalid),.reorder_tdata(reorder_tdata),.current_active(current_active),.traceback_tlast(traceback_tlast[0:0]),.reorder_last_tuser(reorder_last_tuser[0:0]),.buffer_cnt_1(\gen_inst_reorder.0.inst_reorder.buffer_cnt [1:1]),.buffer_cnt_2(\gen_inst_reorder.0.inst_reorder.buffer_cnt [2:2]),.buffer_cnt_0(\gen_inst_reorder.0.inst_reorder.buffer_cnt [0:0]),.traceback_tdata(traceback_tdata[0:0]),.reorder_tvalid_0_rep1(reorder_tvalid_0_rep1),.reorder_tvalid_0_rep2(reorder_tvalid_0_rep2),.m_axis_output_tready(m_axis_output_tready),.N_99(N_99),.aresetn(aresetn),.aclk(aclk),.aresetn_i(aresetn_i),.last_window(\gen_inst_reorder.0.inst_reorder.last_window ),.N_129(N_129));
endmodule
