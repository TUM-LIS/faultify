`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[110:0] testVector;
output[201:0] resultVector;
input[1439:0] injectionVector;
qr_wrapper_wrapper_inj toplevel_instance (
.IN0A0R(testVector [47:0]),
.IN0A0I(testVector [95:48]),
.SIGMA0IN(testVector [107:96]),
.OUT0Q0R(resultVector [47:0]),
.OUT0Q0I(resultVector [95:48]),
.OUT0R0R(resultVector [143:96]),
.OUT0R0I(resultVector [191:144]),
.PERMUT(resultVector [199:192]),
.CLK(clk),
.RST(rst),
.REDUCED0MATRIX(testVector[108]),
.START(testVector[109]),
.REQUEST0OUT(testVector[110]),
.VALID0OUT(resultVector[200]),
.READY(resultVector[201]),
.p_desc0_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[0]),
.p_desc1_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1]),
.p_desc2_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[2]),
.p_desc3_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[3]),
.p_desc4_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[4]),
.p_desc5_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[5]),
.p_desc6_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[6]),
.p_desc7_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[7]),
.p_desc8_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[8]),
.p_desc9_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[9]),
.p_desc10_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[10]),
.p_desc11_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[11]),
.p_desc12_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[12]),
.p_desc13_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[13]),
.p_desc14_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[14]),
.p_desc15_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[15]),
.p_desc16_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[16]),
.p_desc17_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[17]),
.p_desc18_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[18]),
.p_desc19_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[19]),
.p_desc20_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[20]),
.p_desc21_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[21]),
.p_desc22_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[22]),
.p_desc23_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[23]),
.p_desc24_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[24]),
.p_desc25_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[25]),
.p_desc26_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[26]),
.p_desc27_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[27]),
.p_desc28_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[28]),
.p_desc29_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[29]),
.p_desc30_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[30]),
.p_desc31_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[31]),
.p_desc32_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[32]),
.p_desc33_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[33]),
.p_desc34_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[34]),
.p_desc35_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[35]),
.p_desc36_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[36]),
.p_desc37_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[37]),
.p_desc38_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[38]),
.p_desc39_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[39]),
.p_desc40_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[40]),
.p_desc41_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[41]),
.p_desc42_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[42]),
.p_desc43_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[43]),
.p_desc44_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[44]),
.p_desc45_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[45]),
.p_desc46_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[46]),
.p_desc47_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[47]),
.p_desc48_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[48]),
.p_desc49_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[49]),
.p_desc50_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[50]),
.p_desc51_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[51]),
.p_desc52_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[52]),
.p_desc53_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[53]),
.p_desc54_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[54]),
.p_desc55_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[55]),
.p_desc56_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[56]),
.p_desc57_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[57]),
.p_desc58_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[58]),
.p_desc59_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[59]),
.p_desc60_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[60]),
.p_desc61_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[61]),
.p_desc62_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[62]),
.p_desc63_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[63]),
.p_desc64_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[64]),
.p_desc65_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[65]),
.p_desc66_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[66]),
.p_desc67_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[67]),
.p_desc68_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[68]),
.p_desc69_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[69]),
.p_desc70_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[70]),
.p_desc71_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[71]),
.p_desc72_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[72]),
.p_desc73_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[73]),
.p_desc74_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[74]),
.p_desc75_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[75]),
.p_desc76_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[76]),
.p_desc77_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[77]),
.p_desc78_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[78]),
.p_desc79_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[79]),
.p_desc80_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[80]),
.p_desc81_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[81]),
.p_desc82_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[82]),
.p_desc83_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[83]),
.p_desc84_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[84]),
.p_desc85_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[85]),
.p_desc86_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[86]),
.p_desc87_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[87]),
.p_desc88_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[88]),
.p_desc89_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[89]),
.p_desc90_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[90]),
.p_desc91_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[91]),
.p_desc92_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[92]),
.p_desc93_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[93]),
.p_desc94_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[94]),
.p_desc95_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[95]),
.p_desc96_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[96]),
.p_desc97_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[97]),
.p_desc98_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[98]),
.p_desc99_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[99]),
.p_desc100_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[100]),
.p_desc101_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[101]),
.p_desc102_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[102]),
.p_desc103_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[103]),
.p_desc104_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[104]),
.p_desc105_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[105]),
.p_desc106_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[106]),
.p_desc107_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[107]),
.p_desc108_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[108]),
.p_desc109_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[109]),
.p_desc110_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[110]),
.p_desc111_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[111]),
.p_desc112_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[112]),
.p_desc113_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[113]),
.p_desc114_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[114]),
.p_desc115_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[115]),
.p_desc116_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[116]),
.p_desc117_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[117]),
.p_desc118_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[118]),
.p_desc119_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[119]),
.p_desc120_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[120]),
.p_desc121_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[121]),
.p_desc122_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[122]),
.p_desc123_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[123]),
.p_desc124_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[124]),
.p_desc125_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[125]),
.p_desc126_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[126]),
.p_desc127_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[127]),
.p_desc128_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[128]),
.p_desc129_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[129]),
.p_desc130_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[130]),
.p_desc131_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[131]),
.p_desc132_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[132]),
.p_desc133_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[133]),
.p_desc134_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[134]),
.p_desc135_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[135]),
.p_desc136_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[136]),
.p_desc137_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[137]),
.p_desc138_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[138]),
.p_desc139_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[139]),
.p_desc140_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[140]),
.p_desc141_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[141]),
.p_desc142_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[142]),
.p_desc143_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[143]),
.p_desc144_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[144]),
.p_desc145_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[145]),
.p_desc146_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[146]),
.p_desc147_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[147]),
.p_desc148_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[148]),
.p_desc149_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[149]),
.p_desc150_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[150]),
.p_desc151_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[151]),
.p_desc152_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[152]),
.p_desc153_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[153]),
.p_desc154_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[154]),
.p_desc155_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[155]),
.p_desc156_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[156]),
.p_desc157_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[157]),
.p_desc158_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[158]),
.p_desc159_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[159]),
.p_desc160_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[160]),
.p_desc161_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[161]),
.p_desc162_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[162]),
.p_desc163_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[163]),
.p_desc164_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[164]),
.p_desc165_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[165]),
.p_desc166_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[166]),
.p_desc167_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[167]),
.p_desc168_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[168]),
.p_desc169_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[169]),
.p_desc170_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[170]),
.p_desc171_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[171]),
.p_desc172_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[172]),
.p_desc173_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[173]),
.p_desc174_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[174]),
.p_desc175_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[175]),
.p_desc176_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[176]),
.p_desc177_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[177]),
.p_desc178_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[178]),
.p_desc179_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[179]),
.p_desc180_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[180]),
.p_desc181_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[181]),
.p_desc182_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[182]),
.p_desc183_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[183]),
.p_desc184_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[184]),
.p_desc185_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[185]),
.p_desc186_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[186]),
.p_desc187_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[187]),
.p_desc188_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[188]),
.p_desc189_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[189]),
.p_desc190_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[190]),
.p_desc191_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[191]),
.p_desc192_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[192]),
.p_desc193_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[193]),
.p_desc194_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[194]),
.p_desc195_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[195]),
.p_desc196_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[196]),
.p_desc197_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[197]),
.p_desc198_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[198]),
.p_desc199_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[199]),
.p_desc200_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[200]),
.p_desc201_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[201]),
.p_desc202_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[202]),
.p_desc203_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[203]),
.p_desc204_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[204]),
.p_desc205_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[205]),
.p_desc206_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[206]),
.p_desc207_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[207]),
.p_desc208_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[208]),
.p_desc209_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[209]),
.p_desc210_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[210]),
.p_desc211_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[211]),
.p_desc212_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[212]),
.p_desc213_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[213]),
.p_desc214_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[214]),
.p_desc215_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[215]),
.p_desc216_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[216]),
.p_desc217_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[217]),
.p_desc218_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[218]),
.p_desc219_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[219]),
.p_desc220_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[220]),
.p_desc221_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[221]),
.p_desc222_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[222]),
.p_desc223_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[223]),
.p_desc224_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[224]),
.p_desc225_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[225]),
.p_desc226_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[226]),
.p_desc227_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[227]),
.p_desc228_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[228]),
.p_desc229_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[229]),
.p_desc230_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[230]),
.p_desc231_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[231]),
.p_desc232_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[232]),
.p_desc233_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[233]),
.p_desc234_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[234]),
.p_desc235_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[235]),
.p_desc236_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[236]),
.p_desc237_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[237]),
.p_desc238_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[238]),
.p_desc239_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[239]),
.p_desc240_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[240]),
.p_desc241_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[241]),
.p_desc242_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[242]),
.p_desc243_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[243]),
.p_desc244_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[244]),
.p_desc245_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[245]),
.p_desc246_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[246]),
.p_desc247_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[247]),
.p_desc248_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[248]),
.p_desc249_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[249]),
.p_desc250_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[250]),
.p_desc251_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[251]),
.p_desc252_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[252]),
.p_desc253_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[253]),
.p_desc254_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[254]),
.p_desc255_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[255]),
.p_desc256_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[256]),
.p_desc257_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[257]),
.p_desc258_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[258]),
.p_desc259_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[259]),
.p_desc260_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[260]),
.p_desc261_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[261]),
.p_desc262_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[262]),
.p_desc263_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[263]),
.p_desc264_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[264]),
.p_desc265_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[265]),
.p_desc266_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[266]),
.p_desc267_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[267]),
.p_desc268_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[268]),
.p_desc269_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[269]),
.p_desc270_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[270]),
.p_desc271_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[271]),
.p_desc272_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[272]),
.p_desc273_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[273]),
.p_desc274_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[274]),
.p_desc275_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[275]),
.p_desc276_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[276]),
.p_desc277_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[277]),
.p_desc278_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[278]),
.p_desc279_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[279]),
.p_desc280_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[280]),
.p_desc281_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[281]),
.p_desc282_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[282]),
.p_desc283_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[283]),
.p_desc284_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[284]),
.p_desc285_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[285]),
.p_desc286_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[286]),
.p_desc287_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[287]),
.p_desc288_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[288]),
.p_desc289_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[289]),
.p_desc290_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[290]),
.p_desc291_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[291]),
.p_desc292_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[292]),
.p_desc293_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[293]),
.p_desc294_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[294]),
.p_desc295_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[295]),
.p_desc296_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[296]),
.p_desc297_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[297]),
.p_desc298_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[298]),
.p_desc299_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[299]),
.p_desc300_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[300]),
.p_desc301_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[301]),
.p_desc302_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[302]),
.p_desc303_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[303]),
.p_desc304_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[304]),
.p_desc305_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[305]),
.p_desc306_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[306]),
.p_desc307_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[307]),
.p_desc308_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[308]),
.p_desc309_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[309]),
.p_desc310_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[310]),
.p_desc311_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[311]),
.p_desc312_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[312]),
.p_desc313_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[313]),
.p_desc314_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[314]),
.p_desc315_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[315]),
.p_desc316_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[316]),
.p_desc317_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[317]),
.p_desc318_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[318]),
.p_desc319_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[319]),
.p_desc320_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[320]),
.p_desc321_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[321]),
.p_desc322_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[322]),
.p_desc323_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[323]),
.p_desc324_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[324]),
.p_desc325_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[325]),
.p_desc326_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[326]),
.p_desc327_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[327]),
.p_desc328_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[328]),
.p_desc329_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[329]),
.p_desc330_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[330]),
.p_desc331_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[331]),
.p_desc332_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[332]),
.p_desc333_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[333]),
.p_desc334_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[334]),
.p_desc335_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[335]),
.p_desc336_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[336]),
.p_desc337_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[337]),
.p_desc338_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[338]),
.p_desc339_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[339]),
.p_desc340_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[340]),
.p_desc341_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[341]),
.p_desc342_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[342]),
.p_desc343_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[343]),
.p_desc344_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[344]),
.p_desc345_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[345]),
.p_desc346_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[346]),
.p_desc347_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[347]),
.p_desc348_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[348]),
.p_desc349_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[349]),
.p_desc350_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[350]),
.p_desc351_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[351]),
.p_desc352_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[352]),
.p_desc353_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[353]),
.p_desc354_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[354]),
.p_desc355_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[355]),
.p_desc356_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[356]),
.p_desc357_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[357]),
.p_desc358_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[358]),
.p_desc359_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[359]),
.p_desc360_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[360]),
.p_desc361_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[361]),
.p_desc362_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[362]),
.p_desc363_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[363]),
.p_desc364_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[364]),
.p_desc365_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[365]),
.p_desc366_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[366]),
.p_desc367_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[367]),
.p_desc368_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[368]),
.p_desc369_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[369]),
.p_desc370_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[370]),
.p_desc371_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[371]),
.p_desc372_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[372]),
.p_desc373_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[373]),
.p_desc374_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[374]),
.p_desc375_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[375]),
.p_desc376_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[376]),
.p_desc377_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[377]),
.p_desc378_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[378]),
.p_desc379_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[379]),
.p_desc380_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[380]),
.p_desc381_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[381]),
.p_desc382_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[382]),
.p_desc383_p_O_DFFX1mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[383]),
.p_desc384_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[384]),
.p_desc385_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[385]),
.p_desc386_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[386]),
.p_desc387_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[387]),
.p_desc388_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[388]),
.p_desc389_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[389]),
.p_desc390_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[390]),
.p_desc391_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[391]),
.p_desc392_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[392]),
.p_desc393_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[393]),
.p_desc394_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[394]),
.p_desc395_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[395]),
.p_desc396_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[396]),
.p_desc397_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[397]),
.p_desc398_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[398]),
.p_desc399_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[399]),
.p_desc400_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[400]),
.p_desc401_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[401]),
.p_desc402_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[402]),
.p_desc403_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[403]),
.p_desc404_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[404]),
.p_desc405_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[405]),
.p_desc406_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[406]),
.p_desc407_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[407]),
.p_desc408_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[408]),
.p_desc409_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[409]),
.p_desc410_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[410]),
.p_desc411_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[411]),
.p_desc412_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[412]),
.p_desc413_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[413]),
.p_desc414_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[414]),
.p_desc415_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[415]),
.p_desc416_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[416]),
.p_desc417_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[417]),
.p_desc418_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[418]),
.p_desc419_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[419]),
.p_desc420_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[420]),
.p_desc421_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[421]),
.p_desc422_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[422]),
.p_desc423_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[423]),
.p_desc424_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[424]),
.p_desc425_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[425]),
.p_desc426_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[426]),
.p_desc427_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[427]),
.p_desc428_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[428]),
.p_desc429_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[429]),
.p_desc430_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[430]),
.p_desc431_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[431]),
.p_desc432_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[432]),
.p_desc433_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[433]),
.p_desc434_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[434]),
.p_desc435_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[435]),
.p_desc436_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[436]),
.p_desc437_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[437]),
.p_desc438_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[438]),
.p_desc439_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[439]),
.p_desc440_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[440]),
.p_desc441_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[441]),
.p_desc442_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[442]),
.p_desc443_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[443]),
.p_desc444_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[444]),
.p_desc445_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[445]),
.p_desc446_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[446]),
.p_desc447_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[447]),
.p_desc448_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[448]),
.p_desc449_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[449]),
.p_desc450_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[450]),
.p_desc451_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[451]),
.p_desc452_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[452]),
.p_desc453_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[453]),
.p_desc454_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[454]),
.p_desc455_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[455]),
.p_desc456_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[456]),
.p_desc457_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[457]),
.p_desc458_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[458]),
.p_desc459_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[459]),
.p_desc460_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[460]),
.p_desc461_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[461]),
.p_desc462_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[462]),
.p_desc463_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[463]),
.p_desc464_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[464]),
.p_desc465_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[465]),
.p_desc466_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[466]),
.p_desc467_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[467]),
.p_desc468_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[468]),
.p_desc469_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[469]),
.p_desc470_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[470]),
.p_desc471_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[471]),
.p_desc472_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[472]),
.p_desc473_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[473]),
.p_desc474_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[474]),
.p_desc475_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[475]),
.p_desc476_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[476]),
.p_desc477_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[477]),
.p_desc478_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[478]),
.p_desc479_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[479]),
.p_desc480_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[480]),
.p_desc481_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[481]),
.p_desc482_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[482]),
.p_desc483_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[483]),
.p_desc484_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[484]),
.p_desc485_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[485]),
.p_desc486_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[486]),
.p_desc487_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[487]),
.p_desc488_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[488]),
.p_desc489_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[489]),
.p_desc490_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[490]),
.p_desc491_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[491]),
.p_desc492_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[492]),
.p_desc493_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[493]),
.p_desc494_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[494]),
.p_desc495_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[495]),
.p_desc496_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[496]),
.p_desc497_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[497]),
.p_desc498_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[498]),
.p_desc499_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[499]),
.p_desc500_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[500]),
.p_desc501_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[501]),
.p_desc502_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[502]),
.p_desc503_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[503]),
.p_desc504_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[504]),
.p_desc505_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[505]),
.p_desc506_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[506]),
.p_desc507_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[507]),
.p_desc508_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[508]),
.p_desc509_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[509]),
.p_desc510_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[510]),
.p_desc511_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[511]),
.p_desc512_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[512]),
.p_desc513_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[513]),
.p_desc514_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[514]),
.p_desc515_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[515]),
.p_desc516_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[516]),
.p_desc517_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[517]),
.p_desc518_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[518]),
.p_desc519_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[519]),
.p_desc520_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[520]),
.p_desc521_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[521]),
.p_desc522_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[522]),
.p_desc523_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[523]),
.p_desc524_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[524]),
.p_desc525_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[525]),
.p_desc526_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[526]),
.p_desc527_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[527]),
.p_desc528_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[528]),
.p_desc529_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[529]),
.p_desc530_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[530]),
.p_desc531_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[531]),
.p_desc532_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[532]),
.p_desc533_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[533]),
.p_desc534_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[534]),
.p_desc535_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[535]),
.p_desc536_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[536]),
.p_desc537_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[537]),
.p_desc538_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[538]),
.p_desc539_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[539]),
.p_desc540_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[540]),
.p_desc541_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[541]),
.p_desc542_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[542]),
.p_desc543_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[543]),
.p_desc544_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[544]),
.p_desc545_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[545]),
.p_desc546_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[546]),
.p_desc547_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[547]),
.p_desc548_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[548]),
.p_desc549_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[549]),
.p_desc550_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[550]),
.p_desc551_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[551]),
.p_desc552_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[552]),
.p_desc553_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[553]),
.p_desc554_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[554]),
.p_desc555_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[555]),
.p_desc556_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[556]),
.p_desc557_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[557]),
.p_desc558_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[558]),
.p_desc559_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[559]),
.p_desc560_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[560]),
.p_desc561_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[561]),
.p_desc562_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[562]),
.p_desc563_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[563]),
.p_desc564_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[564]),
.p_desc565_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[565]),
.p_desc566_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[566]),
.p_desc567_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[567]),
.p_desc568_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[568]),
.p_desc569_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[569]),
.p_desc570_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[570]),
.p_desc571_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[571]),
.p_desc572_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[572]),
.p_desc573_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[573]),
.p_desc574_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[574]),
.p_desc575_p_O_DFFX1r_mat_regs_WORD_WIDTH12_N4_LOG2_N2_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[575]),
.p_desc576_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[576]),
.p_desc577_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[577]),
.p_desc578_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[578]),
.p_desc579_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[579]),
.p_desc580_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[580]),
.p_desc581_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[581]),
.p_desc582_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[582]),
.p_desc583_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[583]),
.p_desc584_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[584]),
.p_desc585_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[585]),
.p_desc586_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[586]),
.p_desc587_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[587]),
.p_desc588_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[588]),
.p_desc589_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[589]),
.p_desc590_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[590]),
.p_desc591_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[591]),
.p_desc592_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[592]),
.p_desc593_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[593]),
.p_desc594_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[594]),
.p_desc595_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[595]),
.p_desc596_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[596]),
.p_desc597_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[597]),
.p_desc598_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[598]),
.p_desc599_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_19_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[599]),
.p_desc600_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[600]),
.p_desc601_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[601]),
.p_desc602_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[602]),
.p_desc603_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[603]),
.p_desc604_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[604]),
.p_desc605_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[605]),
.p_desc606_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[606]),
.p_desc607_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[607]),
.p_desc608_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[608]),
.p_desc609_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[609]),
.p_desc610_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[610]),
.p_desc611_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[611]),
.p_desc612_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[612]),
.p_desc613_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[613]),
.p_desc614_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[614]),
.p_desc615_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[615]),
.p_desc616_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[616]),
.p_desc617_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[617]),
.p_desc618_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[618]),
.p_desc619_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[619]),
.p_desc620_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[620]),
.p_desc621_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[621]),
.p_desc622_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[622]),
.p_desc623_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_18_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[623]),
.p_desc624_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[624]),
.p_desc625_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[625]),
.p_desc626_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[626]),
.p_desc627_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[627]),
.p_desc628_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[628]),
.p_desc629_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[629]),
.p_desc630_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[630]),
.p_desc631_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[631]),
.p_desc632_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[632]),
.p_desc633_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[633]),
.p_desc634_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[634]),
.p_desc635_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[635]),
.p_desc636_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[636]),
.p_desc637_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[637]),
.p_desc638_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[638]),
.p_desc639_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[639]),
.p_desc640_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[640]),
.p_desc641_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[641]),
.p_desc642_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[642]),
.p_desc643_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[643]),
.p_desc644_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[644]),
.p_desc645_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[645]),
.p_desc646_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[646]),
.p_desc647_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_17_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[647]),
.p_desc648_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[648]),
.p_desc649_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[649]),
.p_desc650_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[650]),
.p_desc651_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[651]),
.p_desc652_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[652]),
.p_desc653_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[653]),
.p_desc654_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[654]),
.p_desc655_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[655]),
.p_desc656_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[656]),
.p_desc657_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[657]),
.p_desc658_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[658]),
.p_desc659_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[659]),
.p_desc660_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[660]),
.p_desc661_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[661]),
.p_desc662_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[662]),
.p_desc663_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[663]),
.p_desc664_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[664]),
.p_desc665_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[665]),
.p_desc666_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[666]),
.p_desc667_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[667]),
.p_desc668_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[668]),
.p_desc669_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[669]),
.p_desc670_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[670]),
.p_desc671_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_16_complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[671]),
.p_desc672_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[672]),
.p_desc673_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[673]),
.p_desc674_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[674]),
.p_desc675_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[675]),
.p_desc676_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[676]),
.p_desc677_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[677]),
.p_desc678_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[678]),
.p_desc679_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[679]),
.p_desc680_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[680]),
.p_desc681_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[681]),
.p_desc682_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[682]),
.p_desc683_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[683]),
.p_desc684_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[684]),
.p_desc685_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[685]),
.p_desc686_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[686]),
.p_desc687_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[687]),
.p_desc688_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[688]),
.p_desc689_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[689]),
.p_desc690_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[690]),
.p_desc691_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[691]),
.p_desc692_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[692]),
.p_desc693_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[693]),
.p_desc694_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[694]),
.p_desc695_p_O_DFFX1complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_inner_prod_INT_BITS4_WORD_WIDTH12_N4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[695]),
.p_desc776_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[696]),
.p_desc777_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[697]),
.p_desc778_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[698]),
.p_desc779_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[699]),
.p_desc780_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[700]),
.p_desc781_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[701]),
.p_desc782_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[702]),
.p_desc783_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[703]),
.p_desc784_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[704]),
.p_desc785_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[705]),
.p_desc786_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[706]),
.p_desc787_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[707]),
.p_desc788_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[708]),
.p_desc789_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[709]),
.p_desc790_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[710]),
.p_desc791_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[711]),
.p_desc792_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[712]),
.p_desc793_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[713]),
.p_desc794_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[714]),
.p_desc795_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[715]),
.p_desc796_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[716]),
.p_desc797_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[717]),
.p_desc798_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[718]),
.p_desc799_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_15_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[719]),
.p_desc800_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[720]),
.p_desc801_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[721]),
.p_desc802_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[722]),
.p_desc803_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[723]),
.p_desc804_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[724]),
.p_desc805_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[725]),
.p_desc806_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[726]),
.p_desc807_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[727]),
.p_desc808_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[728]),
.p_desc809_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[729]),
.p_desc810_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[730]),
.p_desc811_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[731]),
.p_desc812_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[732]),
.p_desc813_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[733]),
.p_desc814_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[734]),
.p_desc815_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[735]),
.p_desc816_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[736]),
.p_desc817_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[737]),
.p_desc818_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[738]),
.p_desc819_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[739]),
.p_desc820_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[740]),
.p_desc821_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[741]),
.p_desc822_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[742]),
.p_desc823_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_14_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[743]),
.p_desc824_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[744]),
.p_desc825_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[745]),
.p_desc826_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[746]),
.p_desc827_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[747]),
.p_desc828_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[748]),
.p_desc829_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[749]),
.p_desc830_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[750]),
.p_desc831_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[751]),
.p_desc832_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[752]),
.p_desc833_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[753]),
.p_desc834_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[754]),
.p_desc835_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[755]),
.p_desc836_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[756]),
.p_desc837_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[757]),
.p_desc838_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[758]),
.p_desc839_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[759]),
.p_desc840_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[760]),
.p_desc841_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[761]),
.p_desc842_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[762]),
.p_desc843_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[763]),
.p_desc844_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[764]),
.p_desc845_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[765]),
.p_desc846_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[766]),
.p_desc847_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_13_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[767]),
.p_desc848_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[768]),
.p_desc849_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[769]),
.p_desc850_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[770]),
.p_desc851_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[771]),
.p_desc852_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[772]),
.p_desc853_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[773]),
.p_desc854_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[774]),
.p_desc855_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[775]),
.p_desc856_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[776]),
.p_desc857_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[777]),
.p_desc858_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[778]),
.p_desc859_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[779]),
.p_desc860_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[780]),
.p_desc861_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[781]),
.p_desc862_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[782]),
.p_desc863_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[783]),
.p_desc864_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[784]),
.p_desc865_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[785]),
.p_desc866_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[786]),
.p_desc867_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[787]),
.p_desc868_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[788]),
.p_desc869_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[789]),
.p_desc870_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[790]),
.p_desc871_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_12_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[791]),
.p_desc872_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[792]),
.p_desc873_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[793]),
.p_desc874_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[794]),
.p_desc875_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[795]),
.p_desc876_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[796]),
.p_desc877_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[797]),
.p_desc878_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[798]),
.p_desc879_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[799]),
.p_desc880_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[800]),
.p_desc881_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[801]),
.p_desc882_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[802]),
.p_desc883_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[803]),
.p_desc884_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[804]),
.p_desc885_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[805]),
.p_desc886_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[806]),
.p_desc887_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[807]),
.p_desc888_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[808]),
.p_desc889_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[809]),
.p_desc890_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[810]),
.p_desc891_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[811]),
.p_desc892_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[812]),
.p_desc893_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[813]),
.p_desc894_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[814]),
.p_desc895_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[815]),
.p_desc896_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[816]),
.p_desc897_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[817]),
.p_desc898_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[818]),
.p_desc899_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[819]),
.p_desc900_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[820]),
.p_desc901_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[821]),
.p_desc902_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[822]),
.p_desc903_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[823]),
.p_desc904_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[824]),
.p_desc905_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[825]),
.p_desc906_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[826]),
.p_desc907_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[827]),
.p_desc908_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[828]),
.p_desc909_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[829]),
.p_desc910_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[830]),
.p_desc911_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[831]),
.p_desc912_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[832]),
.p_desc913_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[833]),
.p_desc914_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[834]),
.p_desc915_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[835]),
.p_desc916_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[836]),
.p_desc917_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[837]),
.p_desc918_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[838]),
.p_desc919_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_11_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[839]),
.p_desc920_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[840]),
.p_desc921_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[841]),
.p_desc922_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[842]),
.p_desc923_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[843]),
.p_desc924_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[844]),
.p_desc925_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[845]),
.p_desc926_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[846]),
.p_desc927_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[847]),
.p_desc928_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[848]),
.p_desc929_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[849]),
.p_desc930_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[850]),
.p_desc931_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[851]),
.p_desc932_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[852]),
.p_desc933_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[853]),
.p_desc934_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[854]),
.p_desc935_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[855]),
.p_desc936_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[856]),
.p_desc937_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[857]),
.p_desc938_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[858]),
.p_desc939_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[859]),
.p_desc940_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[860]),
.p_desc941_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[861]),
.p_desc942_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[862]),
.p_desc943_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_10_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[863]),
.p_desc944_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[864]),
.p_desc945_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[865]),
.p_desc946_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[866]),
.p_desc947_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[867]),
.p_desc948_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[868]),
.p_desc949_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[869]),
.p_desc950_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[870]),
.p_desc951_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[871]),
.p_desc952_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[872]),
.p_desc953_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[873]),
.p_desc954_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[874]),
.p_desc955_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[875]),
.p_desc956_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[876]),
.p_desc957_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[877]),
.p_desc958_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[878]),
.p_desc959_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[879]),
.p_desc960_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[880]),
.p_desc961_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[881]),
.p_desc962_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[882]),
.p_desc963_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[883]),
.p_desc964_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[884]),
.p_desc965_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[885]),
.p_desc966_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[886]),
.p_desc967_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_9_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[887]),
.p_desc968_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[888]),
.p_desc969_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[889]),
.p_desc970_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[890]),
.p_desc971_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[891]),
.p_desc972_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[892]),
.p_desc973_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[893]),
.p_desc974_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[894]),
.p_desc975_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[895]),
.p_desc976_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[896]),
.p_desc977_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[897]),
.p_desc978_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[898]),
.p_desc979_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[899]),
.p_desc980_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[900]),
.p_desc981_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[901]),
.p_desc982_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[902]),
.p_desc983_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[903]),
.p_desc984_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[904]),
.p_desc985_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[905]),
.p_desc986_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[906]),
.p_desc987_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[907]),
.p_desc988_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[908]),
.p_desc989_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[909]),
.p_desc990_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[910]),
.p_desc991_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_8_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[911]),
.p_desc992_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[912]),
.p_desc993_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[913]),
.p_desc994_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[914]),
.p_desc995_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[915]),
.p_desc996_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[916]),
.p_desc997_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[917]),
.p_desc998_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[918]),
.p_desc999_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[919]),
.p_desc1000_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[920]),
.p_desc1001_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[921]),
.p_desc1002_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[922]),
.p_desc1003_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[923]),
.p_desc1004_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[924]),
.p_desc1005_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[925]),
.p_desc1006_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[926]),
.p_desc1007_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[927]),
.p_desc1008_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[928]),
.p_desc1009_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[929]),
.p_desc1010_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[930]),
.p_desc1011_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[931]),
.p_desc1012_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[932]),
.p_desc1013_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[933]),
.p_desc1014_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[934]),
.p_desc1015_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[935]),
.p_desc1016_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[936]),
.p_desc1017_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[937]),
.p_desc1018_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[938]),
.p_desc1019_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[939]),
.p_desc1020_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[940]),
.p_desc1021_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[941]),
.p_desc1022_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[942]),
.p_desc1023_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[943]),
.p_desc1024_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[944]),
.p_desc1025_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[945]),
.p_desc1026_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[946]),
.p_desc1027_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[947]),
.p_desc1028_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[948]),
.p_desc1029_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[949]),
.p_desc1030_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[950]),
.p_desc1031_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[951]),
.p_desc1032_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[952]),
.p_desc1033_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[953]),
.p_desc1034_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[954]),
.p_desc1035_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[955]),
.p_desc1036_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[956]),
.p_desc1037_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[957]),
.p_desc1038_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[958]),
.p_desc1039_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_7_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[959]),
.p_desc1040_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[960]),
.p_desc1041_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[961]),
.p_desc1042_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[962]),
.p_desc1043_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[963]),
.p_desc1044_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[964]),
.p_desc1045_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[965]),
.p_desc1046_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[966]),
.p_desc1047_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[967]),
.p_desc1048_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[968]),
.p_desc1049_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[969]),
.p_desc1050_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[970]),
.p_desc1051_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[971]),
.p_desc1052_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[972]),
.p_desc1053_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[973]),
.p_desc1054_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[974]),
.p_desc1055_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[975]),
.p_desc1056_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[976]),
.p_desc1057_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[977]),
.p_desc1058_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[978]),
.p_desc1059_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[979]),
.p_desc1060_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[980]),
.p_desc1061_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[981]),
.p_desc1062_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[982]),
.p_desc1063_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_6_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[983]),
.p_desc1064_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[984]),
.p_desc1065_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[985]),
.p_desc1066_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[986]),
.p_desc1067_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[987]),
.p_desc1068_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[988]),
.p_desc1069_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[989]),
.p_desc1070_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[990]),
.p_desc1071_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[991]),
.p_desc1072_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[992]),
.p_desc1073_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[993]),
.p_desc1074_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[994]),
.p_desc1075_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[995]),
.p_desc1076_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[996]),
.p_desc1077_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[997]),
.p_desc1078_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[998]),
.p_desc1079_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[999]),
.p_desc1080_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1000]),
.p_desc1081_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1001]),
.p_desc1082_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1002]),
.p_desc1083_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1003]),
.p_desc1084_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1004]),
.p_desc1085_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1005]),
.p_desc1086_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1006]),
.p_desc1087_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_5_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1007]),
.p_desc1088_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1008]),
.p_desc1089_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1009]),
.p_desc1090_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1010]),
.p_desc1091_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1011]),
.p_desc1092_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1012]),
.p_desc1093_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1013]),
.p_desc1094_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1014]),
.p_desc1095_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1015]),
.p_desc1096_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1016]),
.p_desc1097_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1017]),
.p_desc1098_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1018]),
.p_desc1099_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1019]),
.p_desc1100_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1020]),
.p_desc1101_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1021]),
.p_desc1102_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1022]),
.p_desc1103_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1023]),
.p_desc1104_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1024]),
.p_desc1105_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1025]),
.p_desc1106_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1026]),
.p_desc1107_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1027]),
.p_desc1108_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1028]),
.p_desc1109_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1029]),
.p_desc1110_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1030]),
.p_desc1111_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_4_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1031]),
.p_desc1112_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1032]),
.p_desc1113_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1033]),
.p_desc1114_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1034]),
.p_desc1115_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1035]),
.p_desc1116_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1036]),
.p_desc1117_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1037]),
.p_desc1118_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1038]),
.p_desc1119_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1039]),
.p_desc1120_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1040]),
.p_desc1121_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1041]),
.p_desc1122_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1042]),
.p_desc1123_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1043]),
.p_desc1124_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1044]),
.p_desc1125_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1045]),
.p_desc1126_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1046]),
.p_desc1127_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1047]),
.p_desc1128_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1048]),
.p_desc1129_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1049]),
.p_desc1130_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1050]),
.p_desc1131_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1051]),
.p_desc1132_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1052]),
.p_desc1133_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1053]),
.p_desc1134_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1054]),
.p_desc1135_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1055]),
.p_desc1136_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1056]),
.p_desc1137_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1057]),
.p_desc1138_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1058]),
.p_desc1139_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1059]),
.p_desc1140_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1060]),
.p_desc1141_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1061]),
.p_desc1142_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1062]),
.p_desc1143_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1063]),
.p_desc1144_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1064]),
.p_desc1145_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1065]),
.p_desc1146_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1066]),
.p_desc1147_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1067]),
.p_desc1148_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1068]),
.p_desc1149_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1069]),
.p_desc1150_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1070]),
.p_desc1151_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1071]),
.p_desc1152_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1072]),
.p_desc1153_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1073]),
.p_desc1154_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1074]),
.p_desc1155_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1075]),
.p_desc1156_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1076]),
.p_desc1157_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1077]),
.p_desc1158_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1078]),
.p_desc1159_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_3_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1079]),
.p_desc1160_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1080]),
.p_desc1161_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1081]),
.p_desc1162_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1082]),
.p_desc1163_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1083]),
.p_desc1164_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1084]),
.p_desc1165_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1085]),
.p_desc1166_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1086]),
.p_desc1167_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1087]),
.p_desc1168_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1088]),
.p_desc1169_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1089]),
.p_desc1170_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1090]),
.p_desc1171_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1091]),
.p_desc1172_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1092]),
.p_desc1173_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1093]),
.p_desc1174_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1094]),
.p_desc1175_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1095]),
.p_desc1176_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1096]),
.p_desc1177_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1097]),
.p_desc1178_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1098]),
.p_desc1179_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1099]),
.p_desc1180_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1100]),
.p_desc1181_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1101]),
.p_desc1182_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1102]),
.p_desc1183_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_2_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1103]),
.p_desc1184_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1104]),
.p_desc1185_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1105]),
.p_desc1186_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1106]),
.p_desc1187_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1107]),
.p_desc1188_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1108]),
.p_desc1189_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1109]),
.p_desc1190_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1110]),
.p_desc1191_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1111]),
.p_desc1192_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1112]),
.p_desc1193_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1113]),
.p_desc1194_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1114]),
.p_desc1195_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1115]),
.p_desc1196_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1116]),
.p_desc1197_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1117]),
.p_desc1198_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1118]),
.p_desc1199_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1119]),
.p_desc1200_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1120]),
.p_desc1201_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1121]),
.p_desc1202_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1122]),
.p_desc1203_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1123]),
.p_desc1204_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1124]),
.p_desc1205_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1125]),
.p_desc1206_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1126]),
.p_desc1207_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_1_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1127]),
.p_desc1208_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1128]),
.p_desc1209_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1129]),
.p_desc1210_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1130]),
.p_desc1211_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1131]),
.p_desc1212_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1132]),
.p_desc1213_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1133]),
.p_desc1214_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1134]),
.p_desc1215_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1135]),
.p_desc1216_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1136]),
.p_desc1217_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1137]),
.p_desc1218_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1138]),
.p_desc1219_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1139]),
.p_desc1220_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1140]),
.p_desc1221_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1141]),
.p_desc1222_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1142]),
.p_desc1223_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1143]),
.p_desc1224_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1144]),
.p_desc1225_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1145]),
.p_desc1226_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1146]),
.p_desc1227_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1147]),
.p_desc1228_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1148]),
.p_desc1229_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1149]),
.p_desc1230_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1150]),
.p_desc1231_p_O_DFFX1mult_pipe_WORD_WIDTH12_INT_BITS4_0_complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1151]),
.p_desc1232_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1152]),
.p_desc1233_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1153]),
.p_desc1234_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1154]),
.p_desc1235_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1155]),
.p_desc1236_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1156]),
.p_desc1237_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1157]),
.p_desc1238_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1158]),
.p_desc1239_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1159]),
.p_desc1240_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1160]),
.p_desc1241_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1161]),
.p_desc1242_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1162]),
.p_desc1243_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1163]),
.p_desc1244_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1164]),
.p_desc1245_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1165]),
.p_desc1246_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1166]),
.p_desc1247_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1167]),
.p_desc1248_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1168]),
.p_desc1249_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1169]),
.p_desc1250_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1170]),
.p_desc1251_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1171]),
.p_desc1252_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1172]),
.p_desc1253_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1173]),
.p_desc1254_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1174]),
.p_desc1255_p_O_DFFX1complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1175]),
.p_desc1256_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1176]),
.p_desc1257_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1177]),
.p_desc1258_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1178]),
.p_desc1259_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1179]),
.p_desc1260_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1180]),
.p_desc1261_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1181]),
.p_desc1262_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1182]),
.p_desc1263_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1183]),
.p_desc1264_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1184]),
.p_desc1265_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1185]),
.p_desc1266_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1186]),
.p_desc1267_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1187]),
.p_desc1268_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1188]),
.p_desc1269_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1189]),
.p_desc1270_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1190]),
.p_desc1271_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1191]),
.p_desc1272_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1192]),
.p_desc1273_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1193]),
.p_desc1274_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1194]),
.p_desc1275_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1195]),
.p_desc1276_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1196]),
.p_desc1277_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1197]),
.p_desc1278_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1198]),
.p_desc1279_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1199]),
.p_desc1280_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1200]),
.p_desc1281_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1201]),
.p_desc1282_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1202]),
.p_desc1283_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1203]),
.p_desc1284_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1204]),
.p_desc1285_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1205]),
.p_desc1286_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1206]),
.p_desc1287_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1207]),
.p_desc1288_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1208]),
.p_desc1289_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1209]),
.p_desc1290_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1210]),
.p_desc1291_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1211]),
.p_desc1292_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1212]),
.p_desc1293_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1213]),
.p_desc1294_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1214]),
.p_desc1295_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1215]),
.p_desc1296_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1216]),
.p_desc1297_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1217]),
.p_desc1298_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1218]),
.p_desc1299_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1219]),
.p_desc1300_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1220]),
.p_desc1301_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1221]),
.p_desc1302_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1222]),
.p_desc1303_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1223]),
.p_desc1304_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1224]),
.p_desc1305_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1225]),
.p_desc1306_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1226]),
.p_desc1307_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1227]),
.p_desc1308_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1228]),
.p_desc1309_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1229]),
.p_desc1310_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1230]),
.p_desc1311_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1231]),
.p_desc1312_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1232]),
.p_desc1313_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1233]),
.p_desc1314_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1234]),
.p_desc1315_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1235]),
.p_desc1316_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1236]),
.p_desc1317_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1237]),
.p_desc1318_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1238]),
.p_desc1319_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1239]),
.p_desc1320_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1240]),
.p_desc1321_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1241]),
.p_desc1322_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1242]),
.p_desc1323_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1243]),
.p_desc1324_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1244]),
.p_desc1325_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1245]),
.p_desc1326_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1246]),
.p_desc1327_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1247]),
.p_desc1328_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1248]),
.p_desc1329_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1249]),
.p_desc1330_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1250]),
.p_desc1331_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1251]),
.p_desc1332_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1252]),
.p_desc1333_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1253]),
.p_desc1334_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1254]),
.p_desc1335_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1255]),
.p_desc1336_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1256]),
.p_desc1337_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1257]),
.p_desc1338_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1258]),
.p_desc1339_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1259]),
.p_desc1340_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1260]),
.p_desc1341_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1261]),
.p_desc1342_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1262]),
.p_desc1343_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1263]),
.p_desc1344_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1264]),
.p_desc1345_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1265]),
.p_desc1346_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1266]),
.p_desc1347_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1267]),
.p_desc1348_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1268]),
.p_desc1349_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1269]),
.p_desc1350_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1270]),
.p_desc1351_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1271]),
.p_desc1352_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1272]),
.p_desc1353_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1273]),
.p_desc1354_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1274]),
.p_desc1355_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1275]),
.p_desc1356_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1276]),
.p_desc1357_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1277]),
.p_desc1358_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1278]),
.p_desc1359_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1279]),
.p_desc1360_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1280]),
.p_desc1361_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1281]),
.p_desc1363_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1282]),
.p_desc1364_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1283]),
.p_desc1365_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1284]),
.p_desc1366_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1285]),
.p_desc1367_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1286]),
.p_desc1368_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1287]),
.p_desc1369_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1288]),
.p_desc1370_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1289]),
.p_desc1371_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1290]),
.p_desc1372_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1291]),
.p_desc1373_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1292]),
.p_desc1374_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1293]),
.p_desc1375_p_O_DFFX1vec_mult_N4_WORD_WIDTH12_INT_BITS4_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1294]),
.p_desc1376_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1295]),
.p_desc1377_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1296]),
.p_desc1378_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1297]),
.p_desc1379_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1298]),
.p_desc1380_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1299]),
.p_desc1381_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1300]),
.p_desc1382_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1301]),
.p_desc1383_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1302]),
.p_desc1384_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1303]),
.p_desc1385_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1304]),
.p_desc1386_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1305]),
.p_desc1387_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1306]),
.p_desc1388_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1307]),
.p_desc1389_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1308]),
.p_desc1390_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1309]),
.p_desc1391_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1310]),
.p_desc1392_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1311]),
.p_desc1393_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1312]),
.p_desc1394_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1313]),
.p_desc1395_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1314]),
.p_desc1396_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1315]),
.p_desc1397_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1316]),
.p_desc1398_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1317]),
.p_desc1399_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1318]),
.p_desc1400_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1319]),
.p_desc1401_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1320]),
.p_desc1402_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1321]),
.p_desc1403_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1322]),
.p_desc1404_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1323]),
.p_desc1405_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1324]),
.p_desc1406_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1325]),
.p_desc1407_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1326]),
.p_desc1408_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1327]),
.p_desc1409_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1328]),
.p_desc1410_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1329]),
.p_desc1411_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1330]),
.p_desc1412_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1331]),
.p_desc1413_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1332]),
.p_desc1414_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1333]),
.p_desc1415_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1334]),
.p_desc1416_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1335]),
.p_desc1417_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1336]),
.p_desc1418_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1337]),
.p_desc1419_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1338]),
.p_desc1420_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1339]),
.p_desc1421_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1340]),
.p_desc1422_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1341]),
.p_desc1423_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1342]),
.p_desc1424_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1343]),
.p_desc1425_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1344]),
.p_desc1426_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1345]),
.p_desc1427_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1346]),
.p_desc1428_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1347]),
.p_desc1429_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1348]),
.p_desc1430_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1349]),
.p_desc1431_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1350]),
.p_desc1432_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1351]),
.p_desc1433_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1352]),
.p_desc1434_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1353]),
.p_desc1435_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1354]),
.p_desc1436_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1355]),
.p_desc1437_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1356]),
.p_desc1438_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1357]),
.p_desc1439_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1358]),
.p_desc1440_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1359]),
.p_desc1441_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1360]),
.p_desc1442_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1361]),
.p_desc1443_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1362]),
.p_desc1444_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1363]),
.p_desc1445_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1364]),
.p_desc1446_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1365]),
.p_desc1447_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1366]),
.p_desc1448_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1367]),
.p_desc1449_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1368]),
.p_desc1450_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1369]),
.p_desc1451_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1370]),
.p_desc1452_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1371]),
.p_desc1453_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1372]),
.p_desc1454_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1373]),
.p_desc1455_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1374]),
.p_desc1456_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1375]),
.p_desc1457_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1376]),
.p_desc1458_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1377]),
.p_desc1459_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1378]),
.p_desc1460_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1379]),
.p_desc1461_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1380]),
.p_desc1462_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1381]),
.p_desc1463_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1382]),
.p_desc1464_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1383]),
.p_desc1465_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1384]),
.p_desc1466_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1385]),
.p_desc1467_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1386]),
.p_desc1468_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1387]),
.p_desc1469_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1388]),
.p_desc1470_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1389]),
.p_desc1471_p_O_DFFX1vec_sub_N4_WORD_WIDTH12_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1390]),
.p_desc1472_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1391]),
.p_desc1473_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1392]),
.p_desc1474_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1393]),
.p_desc1475_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1394]),
.p_desc1476_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1395]),
.p_desc1477_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1396]),
.p_desc1478_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1397]),
.p_desc1479_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1398]),
.p_desc1480_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1399]),
.p_desc1481_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1400]),
.p_desc1482_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1401]),
.p_desc1483_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1402]),
.p_desc1484_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1403]),
.p_desc1485_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1404]),
.p_desc1486_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1405]),
.p_desc1487_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1406]),
.p_desc1488_p_O_DFFX1mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1407]),
.p_desc1493_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1408]),
.p_desc1494_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1409]),
.p_desc1495_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1410]),
.p_desc1496_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1411]),
.p_desc1497_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1412]),
.p_desc1498_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1413]),
.p_desc1499_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1414]),
.p_desc1500_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1415]),
.p_desc1501_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1416]),
.p_desc1502_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1417]),
.p_desc1503_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1418]),
.p_desc1504_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1419]),
.p_desc1505_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1420]),
.p_desc1506_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1421]),
.p_desc1507_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1422]),
.p_desc1510_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1423]),
.p_desc1511_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1424]),
.p_desc1514_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1425]),
.p_desc1515_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1426]),
.p_desc1516_p_O_DFFX1inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1427]),
.p_desc1521_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1428]),
.p_desc1522_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1429]),
.p_desc1523_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1430]),
.p_desc1524_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1431]),
.p_desc1525_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1432]),
.p_desc1526_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1433]),
.p_desc1527_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1434]),
.p_desc1528_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1435]),
.p_desc1529_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1436]),
.p_desc1530_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1437]),
.p_desc1531_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1438]),
.p_desc1532_p_O_DFFX1qr_decomp_ctl_1_qr_decomp_USE_NEWTON1_qr_wrapper_1_(injectionVector[1439]));
endmodule