`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[31:0] testVector;
output[53:0] resultVector;
input[215:0] injectionVector;
b14_inj toplevel_instance (
.clock(clk),
.reset(rst),
.addr(resultVector [19:0]),
.datai(testVector [31:0]),
.datao(resultVector [51:20]),
.rd(resultVector[52]),
.wr(resultVector[53]),
.p_b_Z_p_O_FDC(injectionVector[0]),
.p_desc52_p_O_FDC(injectionVector[1]),
.p_desc53_p_O_FDC(injectionVector[2]),
.p_desc54_p_O_FDC(injectionVector[3]),
.p_desc55_p_O_FDC(injectionVector[4]),
.p_desc56_p_O_FDC(injectionVector[5]),
.p_desc57_p_O_FDC(injectionVector[6]),
.p_desc58_p_O_FDC(injectionVector[7]),
.p_desc59_p_O_FDC(injectionVector[8]),
.p_desc60_p_O_FDC(injectionVector[9]),
.p_desc61_p_O_FDC(injectionVector[10]),
.p_desc62_p_O_FDC(injectionVector[11]),
.p_desc63_p_O_FDC(injectionVector[12]),
.p_desc64_p_O_FDC(injectionVector[13]),
.p_desc65_p_O_FDC(injectionVector[14]),
.p_desc66_p_O_FDC(injectionVector[15]),
.p_desc67_p_O_FDC(injectionVector[16]),
.p_desc68_p_O_FDC(injectionVector[17]),
.p_desc69_p_O_FDC(injectionVector[18]),
.p_desc70_p_O_FDC(injectionVector[19]),
.p_desc71_p_O_FDC(injectionVector[20]),
.p_desc72_p_O_FDC(injectionVector[21]),
.p_desc73_p_O_FDC(injectionVector[22]),
.p_desc74_p_O_FDC(injectionVector[23]),
.p_desc75_p_O_FDC(injectionVector[24]),
.p_desc76_p_O_FDC(injectionVector[25]),
.p_desc77_p_O_FDC(injectionVector[26]),
.p_desc78_p_O_FDC(injectionVector[27]),
.p_desc79_p_O_FDC(injectionVector[28]),
.p_desc80_p_O_FDC(injectionVector[29]),
.p_desc81_p_O_FDC(injectionVector[30]),
.p_desc82_p_O_FDC(injectionVector[31]),
.p_desc83_p_O_FDC(injectionVector[32]),
.p_rd_Z_p_O_FDC(injectionVector[33]),
.p_desc261_p_O_FDC(injectionVector[34]),
.p_wr_Z_p_O_FDC(injectionVector[35]),
.p_desc262_p_O_FDC(injectionVector[36]),
.p_desc50_p_O_FDCE(injectionVector[37]),
.p_desc51_p_O_FDCE(injectionVector[38]),
.p_desc84_p_O_FDCE(injectionVector[39]),
.p_desc85_p_O_FDCE(injectionVector[40]),
.p_desc86_p_O_FDCE(injectionVector[41]),
.p_desc87_p_O_FDCE(injectionVector[42]),
.p_desc88_p_O_FDCE(injectionVector[43]),
.p_desc89_p_O_FDCE(injectionVector[44]),
.p_desc90_p_O_FDCE(injectionVector[45]),
.p_desc91_p_O_FDCE(injectionVector[46]),
.p_desc92_p_O_FDCE(injectionVector[47]),
.p_desc93_p_O_FDCE(injectionVector[48]),
.p_desc94_p_O_FDCE(injectionVector[49]),
.p_desc95_p_O_FDCE(injectionVector[50]),
.p_desc96_p_O_FDCE(injectionVector[51]),
.p_desc97_p_O_FDCE(injectionVector[52]),
.p_desc98_p_O_FDCE(injectionVector[53]),
.p_desc99_p_O_FDCE(injectionVector[54]),
.p_desc100_p_O_FDCE(injectionVector[55]),
.p_desc101_p_O_FDCE(injectionVector[56]),
.p_desc102_p_O_FDCE(injectionVector[57]),
.p_desc103_p_O_FDCE(injectionVector[58]),
.p_desc104_p_O_FDCE(injectionVector[59]),
.p_desc105_p_O_FDCE(injectionVector[60]),
.p_desc106_p_O_FDCE(injectionVector[61]),
.p_desc107_p_O_FDCE(injectionVector[62]),
.p_desc108_p_O_FDCE(injectionVector[63]),
.p_desc109_p_O_FDCE(injectionVector[64]),
.p_desc110_p_O_FDCE(injectionVector[65]),
.p_desc111_p_O_FDCE(injectionVector[66]),
.p_desc112_p_O_FDCE(injectionVector[67]),
.p_desc113_p_O_FDCE(injectionVector[68]),
.p_desc114_p_O_FDCE(injectionVector[69]),
.p_desc115_p_O_FDCE(injectionVector[70]),
.p_desc116_p_O_FDCE(injectionVector[71]),
.p_desc117_p_O_FDCE(injectionVector[72]),
.p_desc118_p_O_FDCE(injectionVector[73]),
.p_desc119_p_O_FDCE(injectionVector[74]),
.p_desc120_p_O_FDCE(injectionVector[75]),
.p_desc121_p_O_FDCE(injectionVector[76]),
.p_desc122_p_O_FDCE(injectionVector[77]),
.p_desc123_p_O_FDCE(injectionVector[78]),
.p_desc124_p_O_FDCE(injectionVector[79]),
.p_desc125_p_O_FDCE(injectionVector[80]),
.p_desc126_p_O_FDCE(injectionVector[81]),
.p_desc127_p_O_FDCE(injectionVector[82]),
.p_desc128_p_O_FDCE(injectionVector[83]),
.p_desc129_p_O_FDCE(injectionVector[84]),
.p_desc130_p_O_FDCE(injectionVector[85]),
.p_desc131_p_O_FDCE(injectionVector[86]),
.p_desc132_p_O_FDCE(injectionVector[87]),
.p_desc133_p_O_FDCE(injectionVector[88]),
.p_desc134_p_O_FDCE(injectionVector[89]),
.p_desc135_p_O_FDCE(injectionVector[90]),
.p_desc136_p_O_FDCE(injectionVector[91]),
.p_desc137_p_O_FDCE(injectionVector[92]),
.p_desc138_p_O_FDCE(injectionVector[93]),
.p_desc139_p_O_FDCE(injectionVector[94]),
.p_desc140_p_O_FDCE(injectionVector[95]),
.p_desc141_p_O_FDCE(injectionVector[96]),
.p_desc142_p_O_FDCE(injectionVector[97]),
.p_desc143_p_O_FDCE(injectionVector[98]),
.p_desc144_p_O_FDCE(injectionVector[99]),
.p_desc145_p_O_FDCE(injectionVector[100]),
.p_desc146_p_O_FDCE(injectionVector[101]),
.p_desc147_p_O_FDCE(injectionVector[102]),
.p_desc148_p_O_FDCE(injectionVector[103]),
.p_desc149_p_O_FDCE(injectionVector[104]),
.p_desc150_p_O_FDCE(injectionVector[105]),
.p_desc151_p_O_FDCE(injectionVector[106]),
.p_desc152_p_O_FDCE(injectionVector[107]),
.p_desc153_p_O_FDCE(injectionVector[108]),
.p_desc154_p_O_FDCE(injectionVector[109]),
.p_desc155_p_O_FDCE(injectionVector[110]),
.p_desc156_p_O_FDCE(injectionVector[111]),
.p_desc157_p_O_FDCE(injectionVector[112]),
.p_desc158_p_O_FDCE(injectionVector[113]),
.p_desc159_p_O_FDCE(injectionVector[114]),
.p_desc160_p_O_FDCE(injectionVector[115]),
.p_desc161_p_O_FDCE(injectionVector[116]),
.p_desc162_p_O_FDCE(injectionVector[117]),
.p_desc163_p_O_FDCE(injectionVector[118]),
.p_desc164_p_O_FDCE(injectionVector[119]),
.p_desc165_p_O_FDCE(injectionVector[120]),
.p_desc166_p_O_FDCE(injectionVector[121]),
.p_desc167_p_O_FDCE(injectionVector[122]),
.p_desc168_p_O_FDCE(injectionVector[123]),
.p_desc169_p_O_FDCE(injectionVector[124]),
.p_desc170_p_O_FDCE(injectionVector[125]),
.p_desc171_p_O_FDCE(injectionVector[126]),
.p_desc172_p_O_FDCE(injectionVector[127]),
.p_desc173_p_O_FDCE(injectionVector[128]),
.p_desc174_p_O_FDCE(injectionVector[129]),
.p_desc175_p_O_FDCE(injectionVector[130]),
.p_desc176_p_O_FDCE(injectionVector[131]),
.p_desc177_p_O_FDCE(injectionVector[132]),
.p_desc178_p_O_FDCE(injectionVector[133]),
.p_desc179_p_O_FDCE(injectionVector[134]),
.p_desc180_p_O_FDCE(injectionVector[135]),
.p_desc181_p_O_FDCE(injectionVector[136]),
.p_desc182_p_O_FDCE(injectionVector[137]),
.p_desc183_p_O_FDCE(injectionVector[138]),
.p_desc184_p_O_FDCE(injectionVector[139]),
.p_desc185_p_O_FDCE(injectionVector[140]),
.p_desc186_p_O_FDCE(injectionVector[141]),
.p_desc187_p_O_FDCE(injectionVector[142]),
.p_desc188_p_O_FDCE(injectionVector[143]),
.p_desc189_p_O_FDCE(injectionVector[144]),
.p_desc190_p_O_FDCE(injectionVector[145]),
.p_desc191_p_O_FDCE(injectionVector[146]),
.p_desc192_p_O_FDCE(injectionVector[147]),
.p_desc193_p_O_FDCE(injectionVector[148]),
.p_desc194_p_O_FDCE(injectionVector[149]),
.p_desc195_p_O_FDCE(injectionVector[150]),
.p_desc196_p_O_FDCE(injectionVector[151]),
.p_desc197_p_O_FDCE(injectionVector[152]),
.p_desc198_p_O_FDCE(injectionVector[153]),
.p_desc199_p_O_FDCE(injectionVector[154]),
.p_desc200_p_O_FDCE(injectionVector[155]),
.p_desc201_p_O_FDCE(injectionVector[156]),
.p_desc202_p_O_FDCE(injectionVector[157]),
.p_desc203_p_O_FDCE(injectionVector[158]),
.p_desc204_p_O_FDCE(injectionVector[159]),
.p_desc205_p_O_FDCE(injectionVector[160]),
.p_desc206_p_O_FDCE(injectionVector[161]),
.p_desc207_p_O_FDCE(injectionVector[162]),
.p_desc208_p_O_FDCE(injectionVector[163]),
.p_desc209_p_O_FDCE(injectionVector[164]),
.p_desc210_p_O_FDCE(injectionVector[165]),
.p_desc211_p_O_FDCE(injectionVector[166]),
.p_desc212_p_O_FDCE(injectionVector[167]),
.p_desc213_p_O_FDCE(injectionVector[168]),
.p_desc214_p_O_FDCE(injectionVector[169]),
.p_desc215_p_O_FDCE(injectionVector[170]),
.p_desc216_p_O_FDCE(injectionVector[171]),
.p_desc217_p_O_FDCE(injectionVector[172]),
.p_desc218_p_O_FDCE(injectionVector[173]),
.p_desc219_p_O_FDCE(injectionVector[174]),
.p_desc220_p_O_FDCE(injectionVector[175]),
.p_desc221_p_O_FDCE(injectionVector[176]),
.p_desc222_p_O_FDCE(injectionVector[177]),
.p_desc223_p_O_FDCE(injectionVector[178]),
.p_desc224_p_O_FDCE(injectionVector[179]),
.p_desc225_p_O_FDCE(injectionVector[180]),
.p_desc226_p_O_FDCE(injectionVector[181]),
.p_desc227_p_O_FDCE(injectionVector[182]),
.p_desc228_p_O_FDCE(injectionVector[183]),
.p_desc229_p_O_FDCE(injectionVector[184]),
.p_desc230_p_O_FDCE(injectionVector[185]),
.p_desc231_p_O_FDCE(injectionVector[186]),
.p_desc232_p_O_FDCE(injectionVector[187]),
.p_desc233_p_O_FDCE(injectionVector[188]),
.p_desc234_p_O_FDCE(injectionVector[189]),
.p_desc235_p_O_FDCE(injectionVector[190]),
.p_desc236_p_O_FDCE(injectionVector[191]),
.p_desc237_p_O_FDCE(injectionVector[192]),
.p_desc238_p_O_FDCE(injectionVector[193]),
.p_desc239_p_O_FDCE(injectionVector[194]),
.p_desc240_p_O_FDCE(injectionVector[195]),
.p_desc241_p_O_FDCE(injectionVector[196]),
.p_desc242_p_O_FDCE(injectionVector[197]),
.p_desc243_p_O_FDCE(injectionVector[198]),
.p_desc244_p_O_FDCE(injectionVector[199]),
.p_desc245_p_O_FDCE(injectionVector[200]),
.p_desc246_p_O_FDCE(injectionVector[201]),
.p_desc247_p_O_FDCE(injectionVector[202]),
.p_desc248_p_O_FDCE(injectionVector[203]),
.p_desc249_p_O_FDCE(injectionVector[204]),
.p_desc250_p_O_FDCE(injectionVector[205]),
.p_desc251_p_O_FDCE(injectionVector[206]),
.p_desc252_p_O_FDCE(injectionVector[207]),
.p_desc253_p_O_FDCE(injectionVector[208]),
.p_desc254_p_O_FDCE(injectionVector[209]),
.p_desc255_p_O_FDCE(injectionVector[210]),
.p_desc256_p_O_FDCE(injectionVector[211]),
.p_desc257_p_O_FDCE(injectionVector[212]),
.p_desc258_p_O_FDCE(injectionVector[213]),
.p_desc259_p_O_FDCE(injectionVector[214]),
.p_desc260_p_O_FDCE(injectionVector[215]));
endmodule