`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[7:0] testVector;
output[7:0] resultVector;
input[104:0] injectionVector;
fir_inj toplevel_instance (
.x_in(testVector [7:0]),
.clk(clk),
.y(resultVector [7:0]),
.p_desc0_p_O_FD(injectionVector[0]),
.p_desc1_p_O_FD(injectionVector[1]),
.p_desc2_p_O_FD(injectionVector[2]),
.p_desc3_p_O_FD(injectionVector[3]),
.p_desc4_p_O_FD(injectionVector[4]),
.p_desc5_p_O_FD(injectionVector[5]),
.p_desc6_p_O_FD(injectionVector[6]),
.p_desc7_p_O_FD(injectionVector[7]),
.p_desc8_p_O_FD(injectionVector[8]),
.p_desc9_p_O_FD(injectionVector[9]),
.p_desc10_p_O_FD(injectionVector[10]),
.p_desc11_p_O_FD(injectionVector[11]),
.p_desc12_p_O_FD(injectionVector[12]),
.p_desc13_p_O_FD(injectionVector[13]),
.p_desc14_p_O_FD(injectionVector[14]),
.p_desc15_p_O_FD(injectionVector[15]),
.p_desc16_p_O_FD(injectionVector[16]),
.p_desc17_p_O_FD(injectionVector[17]),
.p_desc18_p_O_FD(injectionVector[18]),
.p_desc19_p_O_FD(injectionVector[19]),
.p_desc20_p_O_FD(injectionVector[20]),
.p_desc21_p_O_FD(injectionVector[21]),
.p_desc22_p_O_FD(injectionVector[22]),
.p_desc23_p_O_FD(injectionVector[23]),
.p_desc24_p_O_FD(injectionVector[24]),
.p_desc25_p_O_FD(injectionVector[25]),
.p_desc26_p_O_FD(injectionVector[26]),
.p_desc27_p_O_FD(injectionVector[27]),
.p_desc28_p_O_FD(injectionVector[28]),
.p_desc29_p_O_FD(injectionVector[29]),
.p_desc30_p_O_FD(injectionVector[30]),
.p_desc31_p_O_FD(injectionVector[31]),
.p_desc32_p_O_FD(injectionVector[32]),
.p_x_14_pipe_0_Z_p_O_FD(injectionVector[33]),
.p_x_14_pipe_9_Z_p_O_FD(injectionVector[34]),
.p_x_14_pipe_10_Z_p_O_FD(injectionVector[35]),
.p_x_14_pipe_11_Z_p_O_FD(injectionVector[36]),
.p_x_14_pipe_12_Z_p_O_FD(injectionVector[37]),
.p_x_14_pipe_13_Z_p_O_FD(injectionVector[38]),
.p_x_14_pipe_14_Z_p_O_FD(injectionVector[39]),
.p_x_14_pipe_15_Z_p_O_FD(injectionVector[40]),
.p_x_14_pipe_16_Z_p_O_FD(injectionVector[41]),
.p_x_14_pipe_17_Z_p_O_FD(injectionVector[42]),
.p_x_9_pipe_1_Z_p_O_FD(injectionVector[43]),
.p_x_9_pipe_2_Z_p_O_FD(injectionVector[44]),
.p_x_9_pipe_3_Z_p_O_FD(injectionVector[45]),
.p_x_9_pipe_4_Z_p_O_FD(injectionVector[46]),
.p_x_9_pipe_5_Z_p_O_FD(injectionVector[47]),
.p_x_9_pipe_6_Z_p_O_FD(injectionVector[48]),
.p_x_9_pipe_7_Z_p_O_FD(injectionVector[49]),
.p_x_9_pipe_8_Z_p_O_FD(injectionVector[50]),
.p_x_15_pipe_0_0_15_Z_p_O_FD(injectionVector[51]),
.p_x_15_pipe_0_0_16_Z_p_O_FD(injectionVector[52]),
.p_x_15_pipe_0_0_17_Z_p_O_FD(injectionVector[53]),
.p_x_15_pipe_0_0_18_Z_p_O_FD(injectionVector[54]),
.p_x_15_pipe_0_0_19_Z_p_O_FD(injectionVector[55]),
.p_x_15_pipe_0_0_20_Z_p_O_FD(injectionVector[56]),
.p_x_15_pipe_0_0_21_Z_p_O_FD(injectionVector[57]),
.p_x_15_pipe_0_0_22_Z_p_O_FD(injectionVector[58]),
.p_x_15_pipe_0_0_23_Z_p_O_FD(injectionVector[59]),
.p_x_15_pipe_0_0_24_Z_p_O_FD(injectionVector[60]),
.p_x_15_pipe_0_0_25_Z_p_O_FD(injectionVector[61]),
.p_x_15_pipe_0_0_26_Z_p_O_FD(injectionVector[62]),
.p_x_15_pipe_0_0_27_Z_p_O_FD(injectionVector[63]),
.p_x_15_pipe_0_0_28_Z_p_O_FD(injectionVector[64]),
.p_x_15_pipe_0_0_29_Z_p_O_FD(injectionVector[65]),
.p_x_16_pipe_0_0_0_Z_p_O_FD(injectionVector[66]),
.p_x_16_pipe_0_0_1_Z_p_O_FD(injectionVector[67]),
.p_x_16_pipe_0_0_2_Z_p_O_FD(injectionVector[68]),
.p_x_16_pipe_0_0_3_Z_p_O_FD(injectionVector[69]),
.p_x_16_pipe_0_0_4_Z_p_O_FD(injectionVector[70]),
.p_x_16_pipe_0_0_5_Z_p_O_FD(injectionVector[71]),
.p_x_16_pipe_0_0_6_Z_p_O_FD(injectionVector[72]),
.p_x_16_pipe_0_0_7_Z_p_O_FD(injectionVector[73]),
.p_x_16_pipe_0_0_8_Z_p_O_FD(injectionVector[74]),
.p_x_16_pipe_0_0_9_Z_p_O_FD(injectionVector[75]),
.p_x_16_pipe_0_0_10_Z_p_O_FD(injectionVector[76]),
.p_x_16_pipe_0_0_11_Z_p_O_FD(injectionVector[77]),
.p_x_16_pipe_0_0_12_Z_p_O_FD(injectionVector[78]),
.p_x_16_pipe_0_0_13_Z_p_O_FD(injectionVector[79]),
.p_x_16_pipe_0_0_14_Z_p_O_FD(injectionVector[80]),
.p_desc33_p_O_FD(injectionVector[81]),
.p_desc34_p_O_FD(injectionVector[82]),
.p_desc35_p_O_FD(injectionVector[83]),
.p_desc36_p_O_FD(injectionVector[84]),
.p_desc37_p_O_FD(injectionVector[85]),
.p_desc38_p_O_FD(injectionVector[86]),
.p_desc39_p_O_FD(injectionVector[87]),
.p_desc40_p_O_FD(injectionVector[88]),
.p_desc41_p_O_FD(injectionVector[89]),
.p_desc42_p_O_FD(injectionVector[90]),
.p_desc43_p_O_FD(injectionVector[91]),
.p_desc44_p_O_FD(injectionVector[92]),
.p_desc45_p_O_FD(injectionVector[93]),
.p_desc46_p_O_FD(injectionVector[94]),
.p_desc47_p_O_FD(injectionVector[95]),
.p_desc48_p_O_FD(injectionVector[96]),
.p_desc49_p_O_FD(injectionVector[97]),
.p_desc50_p_O_FD(injectionVector[98]),
.p_desc51_p_O_FD(injectionVector[99]),
.p_desc52_p_O_FD(injectionVector[100]),
.p_desc53_p_O_FD(injectionVector[101]),
.p_desc54_p_O_FD(injectionVector[102]),
.p_desc55_p_O_FD(injectionVector[103]),
.p_desc56_p_O_FD(injectionVector[104]));
endmodule