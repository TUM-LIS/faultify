`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[141:0] injectionVector;
fpu_inj toplevel_instance (
.clk_i(clk),
.opa_i(testVector [31:0]),
.opb_i(testVector [63:32]),
.fpu_op_i(testVector [66:64]),
.rmode_i(testVector [68:67]),
.output_o(resultVector [31:0]),
.start_i(testVector[69]),
.ready_o(resultVector[32]),
.ine_o(resultVector[33]),
.overflow_o(resultVector[34]),
.underflow_o(resultVector[35]),
.div_zero_o(resultVector[36]),
.inf_o(resultVector[37]),
.zero_o(resultVector[38]),
.qnan_o(resultVector[39]),
.snan_o(resultVector[40]),
.p_desc595_p_O_FDpre_norm_mul_(injectionVector[0]),
.p_desc596_p_O_FDpre_norm_mul_(injectionVector[1]),
.p_desc597_p_O_FDpre_norm_mul_(injectionVector[2]),
.p_desc598_p_O_FDpre_norm_mul_(injectionVector[3]),
.p_desc599_p_O_FDpre_norm_mul_(injectionVector[4]),
.p_desc600_p_O_FDpre_norm_mul_(injectionVector[5]),
.p_desc601_p_O_FDpre_norm_mul_(injectionVector[6]),
.p_desc602_p_O_FDpre_norm_mul_(injectionVector[7]),
.p_desc603_p_O_FDpre_norm_mul_(injectionVector[8]),
.p_desc604_p_O_FDpre_norm_mul_(injectionVector[9]),
.p_desc1070_p_O_FDpost_norm_mul_(injectionVector[10]),
.p_desc1071_p_O_FDpost_norm_mul_(injectionVector[11]),
.p_desc1072_p_O_FDpost_norm_mul_(injectionVector[12]),
.p_desc1073_p_O_FDpost_norm_mul_(injectionVector[13]),
.p_desc1074_p_O_FDpost_norm_mul_(injectionVector[14]),
.p_desc1075_p_O_FDpost_norm_mul_(injectionVector[15]),
.p_desc1076_p_O_FDpost_norm_mul_(injectionVector[16]),
.p_desc1077_p_O_FDpost_norm_mul_(injectionVector[17]),
.p_desc1078_p_O_FDpost_norm_mul_(injectionVector[18]),
.p_desc1079_p_O_FDpost_norm_mul_(injectionVector[19]),
.p_desc1080_p_O_FDpost_norm_mul_(injectionVector[20]),
.p_desc1081_p_O_FDpost_norm_mul_(injectionVector[21]),
.p_desc1082_p_O_FDpost_norm_mul_(injectionVector[22]),
.p_desc1083_p_O_FDpost_norm_mul_(injectionVector[23]),
.p_desc1084_p_O_FDpost_norm_mul_(injectionVector[24]),
.p_desc1085_p_O_FDpost_norm_mul_(injectionVector[25]),
.p_desc1086_p_O_FDpost_norm_mul_(injectionVector[26]),
.p_desc1087_p_O_FDpost_norm_mul_(injectionVector[27]),
.p_desc1088_p_O_FDpost_norm_mul_(injectionVector[28]),
.p_desc1089_p_O_FDpost_norm_mul_(injectionVector[29]),
.p_desc1090_p_O_FDpost_norm_mul_(injectionVector[30]),
.p_desc1091_p_O_FDpost_norm_mul_(injectionVector[31]),
.p_desc1092_p_O_FDpost_norm_mul_(injectionVector[32]),
.p_desc1163_p_O_FDpost_norm_mul_(injectionVector[33]),
.p_desc1164_p_O_FDpost_norm_mul_(injectionVector[34]),
.p_desc1165_p_O_FDpost_norm_mul_(injectionVector[35]),
.p_desc1166_p_O_FDpost_norm_mul_(injectionVector[36]),
.p_desc1167_p_O_FDpost_norm_mul_(injectionVector[37]),
.p_desc1168_p_O_FDpost_norm_mul_(injectionVector[38]),
.p_desc1169_p_O_FDpost_norm_mul_(injectionVector[39]),
.p_desc1170_p_O_FDpost_norm_mul_(injectionVector[40]),
.p_desc1171_p_O_FDpost_norm_mul_(injectionVector[41]),
.p_desc1172_p_O_FDpost_norm_mul_(injectionVector[42]),
.p_desc1173_p_O_FDpost_norm_mul_(injectionVector[43]),
.p_desc1174_p_O_FDpost_norm_mul_(injectionVector[44]),
.p_desc1175_p_O_FDpost_norm_mul_(injectionVector[45]),
.p_desc1176_p_O_FDpost_norm_mul_(injectionVector[46]),
.p_desc1177_p_O_FDpost_norm_mul_(injectionVector[47]),
.p_desc1178_p_O_FDpost_norm_mul_(injectionVector[48]),
.p_desc1179_p_O_FDpost_norm_mul_(injectionVector[49]),
.p_desc1180_p_O_FDpost_norm_mul_(injectionVector[50]),
.p_desc1181_p_O_FDpost_norm_mul_(injectionVector[51]),
.p_desc1182_p_O_FDpost_norm_mul_(injectionVector[52]),
.p_desc1183_p_O_FDpost_norm_mul_(injectionVector[53]),
.p_desc1184_p_O_FDpost_norm_mul_(injectionVector[54]),
.p_desc1185_p_O_FDpost_norm_mul_(injectionVector[55]),
.p_desc1186_p_O_FDpost_norm_mul_(injectionVector[56]),
.p_desc1187_p_O_FDpost_norm_mul_(injectionVector[57]),
.p_desc1188_p_O_FDpost_norm_mul_(injectionVector[58]),
.p_desc1189_p_O_FDpost_norm_mul_(injectionVector[59]),
.p_desc1190_p_O_FDpost_norm_mul_(injectionVector[60]),
.p_desc1191_p_O_FDpost_norm_mul_(injectionVector[61]),
.p_desc1192_p_O_FDpost_norm_mul_(injectionVector[62]),
.p_desc1193_p_O_FDpost_norm_mul_(injectionVector[63]),
.p_desc1194_p_O_FDpost_norm_mul_(injectionVector[64]),
.p_desc1195_p_O_FDpost_norm_mul_(injectionVector[65]),
.p_desc1196_p_O_FDpost_norm_mul_(injectionVector[66]),
.p_desc1197_p_O_FDpost_norm_mul_(injectionVector[67]),
.p_desc1198_p_O_FDpost_norm_mul_(injectionVector[68]),
.p_desc1199_p_O_FDpost_norm_mul_(injectionVector[69]),
.p_desc1200_p_O_FDpost_norm_mul_(injectionVector[70]),
.p_desc1201_p_O_FDpost_norm_mul_(injectionVector[71]),
.p_desc1202_p_O_FDpost_norm_mul_(injectionVector[72]),
.p_desc1203_p_O_FDpost_norm_mul_(injectionVector[73]),
.p_desc1204_p_O_FDpost_norm_mul_(injectionVector[74]),
.p_desc1205_p_O_FDpost_norm_mul_(injectionVector[75]),
.p_desc1206_p_O_FDpost_norm_mul_(injectionVector[76]),
.p_desc1207_p_O_FDpost_norm_mul_(injectionVector[77]),
.p_desc1208_p_O_FDpost_norm_mul_(injectionVector[78]),
.p_desc1209_p_O_FDpost_norm_mul_(injectionVector[79]),
.p_desc1210_p_O_FDpost_norm_mul_(injectionVector[80]),
.p_desc1211_p_O_FDpost_norm_mul_(injectionVector[81]),
.p_desc1212_p_O_FDpost_norm_mul_(injectionVector[82]),
.p_desc1213_p_O_FDpost_norm_mul_(injectionVector[83]),
.p_desc1214_p_O_FDpost_norm_mul_(injectionVector[84]),
.p_desc1215_p_O_FDpost_norm_mul_(injectionVector[85]),
.p_desc1216_p_O_FDpost_norm_mul_(injectionVector[86]),
.p_desc1217_p_O_FDpost_norm_mul_(injectionVector[87]),
.p_desc1218_p_O_FDpost_norm_mul_(injectionVector[88]),
.p_desc1219_p_O_FDpost_norm_mul_(injectionVector[89]),
.p_desc1220_p_O_FDpost_norm_mul_(injectionVector[90]),
.p_desc1221_p_O_FDpost_norm_mul_(injectionVector[91]),
.p_s_sign_i_Z_p_O_FDpost_norm_mul_(injectionVector[92]),
.p_ine_o_Z_p_O_FDpost_norm_mul_(injectionVector[93]),
.p_desc1244_p_O_FDpost_norm_mul_(injectionVector[94]),
.p_desc1245_p_O_FDpost_norm_mul_(injectionVector[95]),
.p_desc1246_p_O_FDpost_norm_mul_(injectionVector[96]),
.p_desc1247_p_O_FDpost_norm_mul_(injectionVector[97]),
.p_desc1248_p_O_FDpost_norm_mul_(injectionVector[98]),
.p_desc1249_p_O_FDpost_norm_mul_(injectionVector[99]),
.p_desc1250_p_O_FDpost_norm_mul_(injectionVector[100]),
.p_desc1251_p_O_FDpost_norm_mul_(injectionVector[101]),
.p_desc1252_p_O_FDpost_norm_mul_(injectionVector[102]),
.p_desc1253_p_O_FDpost_norm_mul_(injectionVector[103]),
.p_desc1254_p_O_FDpost_norm_mul_(injectionVector[104]),
.p_desc1255_p_O_FDpost_norm_mul_(injectionVector[105]),
.p_desc1256_p_O_FDpost_norm_mul_(injectionVector[106]),
.p_desc1257_p_O_FDpost_norm_mul_(injectionVector[107]),
.p_desc1258_p_O_FDpost_norm_mul_(injectionVector[108]),
.p_desc1259_p_O_FDpost_norm_mul_(injectionVector[109]),
.p_desc1260_p_O_FDpost_norm_mul_(injectionVector[110]),
.p_desc1261_p_O_FDpost_norm_mul_(injectionVector[111]),
.p_desc1262_p_O_FDpost_norm_mul_(injectionVector[112]),
.p_desc1263_p_O_FDpost_norm_mul_(injectionVector[113]),
.p_desc1264_p_O_FDpost_norm_mul_(injectionVector[114]),
.p_desc1265_p_O_FDpost_norm_mul_(injectionVector[115]),
.p_desc1266_p_O_FDpost_norm_mul_(injectionVector[116]),
.p_desc1267_p_O_FDpost_norm_mul_(injectionVector[117]),
.p_desc1268_p_O_FDpost_norm_mul_(injectionVector[118]),
.p_desc1269_p_O_FDpost_norm_mul_(injectionVector[119]),
.p_desc1270_p_O_FDpost_norm_mul_(injectionVector[120]),
.p_desc1271_p_O_FDpost_norm_mul_(injectionVector[121]),
.p_desc1272_p_O_FDpost_norm_mul_(injectionVector[122]),
.p_desc1273_p_O_FDpost_norm_mul_(injectionVector[123]),
.p_desc1274_p_O_FDpost_norm_mul_(injectionVector[124]),
.p_desc1275_p_O_FDpost_norm_mul_(injectionVector[125]),
.p_desc1276_p_O_FDpost_norm_mul_(injectionVector[126]),
.p_desc1277_p_O_FDpost_norm_mul_(injectionVector[127]),
.p_desc1278_p_O_FDpost_norm_mul_(injectionVector[128]),
.p_desc1279_p_O_FDpost_norm_mul_(injectionVector[129]),
.p_desc1280_p_O_FDpost_norm_mul_(injectionVector[130]),
.p_desc1281_p_O_FDpost_norm_mul_(injectionVector[131]),
.p_desc1282_p_O_FDpost_norm_mul_(injectionVector[132]),
.p_desc1283_p_O_FDpost_norm_mul_(injectionVector[133]),
.p_desc1284_p_O_FDpost_norm_mul_(injectionVector[134]),
.p_desc1285_p_O_FDpost_norm_mul_(injectionVector[135]),
.p_desc1286_p_O_FDpost_norm_mul_(injectionVector[136]),
.p_desc1287_p_O_FDpost_norm_mul_(injectionVector[137]),
.p_desc1288_p_O_FDpost_norm_mul_(injectionVector[138]),
.p_desc1289_p_O_FDpost_norm_mul_(injectionVector[139]),
.p_desc1290_p_O_FDpost_norm_mul_(injectionVector[140]),
.p_desc1291_p_O_FDpost_norm_mul_(injectionVector[141]));
endmodule