`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[630:0] injectionVector;
fpu_inj toplevel_instance (
.OPA0I(testVector [31:0]),
.OPB0I(testVector [63:32]),
.FPU0OP0I(testVector [66:64]),
.RMODE0I(testVector [68:67]),
.OUTPUT0O(resultVector [31:0]),
.CLK0I(clk),
.START0I(testVector[69]),
.READY0O(resultVector[32]),
.INE0O(resultVector[33]),
.OVERFLOW0O(resultVector[34]),
.UNDERFLOW0O(resultVector[35]),
.DIV0ZERO0O(resultVector[36]),
.INF0O(resultVector[37]),
.ZERO0O(resultVector[38]),
.QNAN0O(resultVector[39]),
.SNAN0O(resultVector[40]),
.p_desc180_p_O_DFFX1pre_norm_mul_1_(injectionVector[0]),
.p_desc181_p_O_DFFX1pre_norm_mul_1_(injectionVector[1]),
.p_desc182_p_O_DFFX1pre_norm_mul_1_(injectionVector[2]),
.p_desc183_p_O_DFFX1pre_norm_mul_1_(injectionVector[3]),
.p_desc184_p_O_DFFX1pre_norm_mul_1_(injectionVector[4]),
.p_desc185_p_O_DFFX1pre_norm_mul_1_(injectionVector[5]),
.p_desc186_p_O_DFFX1pre_norm_mul_1_(injectionVector[6]),
.p_desc187_p_O_DFFX1pre_norm_mul_1_(injectionVector[7]),
.p_desc188_p_O_DFFX1pre_norm_mul_1_(injectionVector[8]),
.p_desc189_p_O_DFFX1pre_norm_mul_1_(injectionVector[9]),
.p_desc190_p_O_DFFX1mul_24_1_(injectionVector[10]),
.p_desc191_p_O_DFFX1mul_24_1_(injectionVector[11]),
.p_desc192_p_O_DFFX1mul_24_1_(injectionVector[12]),
.p_desc193_p_O_DFFX1mul_24_1_(injectionVector[13]),
.p_desc194_p_O_DFFX1mul_24_1_(injectionVector[14]),
.p_desc195_p_O_DFFX1mul_24_1_(injectionVector[15]),
.p_desc196_p_O_DFFX1mul_24_1_(injectionVector[16]),
.p_desc197_p_O_DFFX1mul_24_1_(injectionVector[17]),
.p_desc198_p_O_DFFX1mul_24_1_(injectionVector[18]),
.p_desc199_p_O_DFFX1mul_24_1_(injectionVector[19]),
.p_desc200_p_O_DFFX1mul_24_1_(injectionVector[20]),
.p_desc201_p_O_DFFX1mul_24_1_(injectionVector[21]),
.p_desc202_p_O_DFFX1mul_24_1_(injectionVector[22]),
.p_desc203_p_O_DFFX1mul_24_1_(injectionVector[23]),
.p_desc204_p_O_DFFX1mul_24_1_(injectionVector[24]),
.p_desc205_p_O_DFFX1mul_24_1_(injectionVector[25]),
.p_desc206_p_O_DFFX1mul_24_1_(injectionVector[26]),
.p_desc207_p_O_DFFX1mul_24_1_(injectionVector[27]),
.p_desc208_p_O_DFFX1mul_24_1_(injectionVector[28]),
.p_desc209_p_O_DFFX1mul_24_1_(injectionVector[29]),
.p_desc210_p_O_DFFX1mul_24_1_(injectionVector[30]),
.p_desc211_p_O_DFFX1mul_24_1_(injectionVector[31]),
.p_desc212_p_O_DFFX1mul_24_1_(injectionVector[32]),
.p_desc213_p_O_DFFX1mul_24_1_(injectionVector[33]),
.p_desc214_p_O_DFFX1mul_24_1_(injectionVector[34]),
.p_desc215_p_O_DFFX1mul_24_1_(injectionVector[35]),
.p_desc216_p_O_DFFX1mul_24_1_(injectionVector[36]),
.p_desc217_p_O_DFFX1mul_24_1_(injectionVector[37]),
.p_desc218_p_O_DFFX1mul_24_1_(injectionVector[38]),
.p_desc219_p_O_DFFX1mul_24_1_(injectionVector[39]),
.p_desc220_p_O_DFFX1mul_24_1_(injectionVector[40]),
.p_desc221_p_O_DFFX1mul_24_1_(injectionVector[41]),
.p_desc222_p_O_DFFX1mul_24_1_(injectionVector[42]),
.p_desc223_p_O_DFFX1mul_24_1_(injectionVector[43]),
.p_desc224_p_O_DFFX1mul_24_1_(injectionVector[44]),
.p_desc225_p_O_DFFX1mul_24_1_(injectionVector[45]),
.p_desc226_p_O_DFFX1mul_24_1_(injectionVector[46]),
.p_desc227_p_O_DFFX1mul_24_1_(injectionVector[47]),
.p_desc228_p_O_DFFX1mul_24_1_(injectionVector[48]),
.p_desc229_p_O_DFFX1mul_24_1_(injectionVector[49]),
.p_desc230_p_O_DFFX1mul_24_1_(injectionVector[50]),
.p_desc231_p_O_DFFX1mul_24_1_(injectionVector[51]),
.p_desc232_p_O_DFFX1mul_24_1_(injectionVector[52]),
.p_desc233_p_O_DFFX1mul_24_1_(injectionVector[53]),
.p_desc234_p_O_DFFX1mul_24_1_(injectionVector[54]),
.p_desc235_p_O_DFFX1mul_24_1_(injectionVector[55]),
.p_desc236_p_O_DFFX1mul_24_1_(injectionVector[56]),
.p_desc237_p_O_DFFX1mul_24_1_(injectionVector[57]),
.p_s_signa_i_reg_p_O_DFFX1mul_24_1_(injectionVector[58]),
.p_s_signb_i_reg_p_O_DFFX1mul_24_1_(injectionVector[59]),
.p_s_start_i_reg_p_O_DFFX1mul_24_1_(injectionVector[60]),
.p_desc238_p_O_DFFX1mul_24_1_(injectionVector[61]),
.p_s_state_reg_p_O_DFFX1mul_24_1_(injectionVector[62]),
.p_s_ready_o_reg_p_O_DFFX1mul_24_1_(injectionVector[63]),
.p_desc239_p_O_DFFX1mul_24_1_(injectionVector[64]),
.p_desc240_p_O_DFFX1mul_24_1_(injectionVector[65]),
.p_desc241_p_O_DFFX1mul_24_1_(injectionVector[66]),
.p_desc242_p_O_DFFX1mul_24_1_(injectionVector[67]),
.p_desc243_p_O_DFFX1mul_24_1_(injectionVector[68]),
.p_desc244_p_O_DFFX1mul_24_1_(injectionVector[69]),
.p_desc245_p_O_DFFX1mul_24_1_(injectionVector[70]),
.p_desc246_p_O_DFFX1mul_24_1_(injectionVector[71]),
.p_desc247_p_O_DFFX1mul_24_1_(injectionVector[72]),
.p_desc248_p_O_DFFX1mul_24_1_(injectionVector[73]),
.p_desc249_p_O_DFFX1mul_24_1_(injectionVector[74]),
.p_desc250_p_O_DFFX1mul_24_1_(injectionVector[75]),
.p_desc251_p_O_DFFX1mul_24_1_(injectionVector[76]),
.p_desc252_p_O_DFFX1mul_24_1_(injectionVector[77]),
.p_desc253_p_O_DFFX1mul_24_1_(injectionVector[78]),
.p_desc254_p_O_DFFX1mul_24_1_(injectionVector[79]),
.p_desc255_p_O_DFFX1mul_24_1_(injectionVector[80]),
.p_desc256_p_O_DFFX1mul_24_1_(injectionVector[81]),
.p_desc257_p_O_DFFX1mul_24_1_(injectionVector[82]),
.p_desc258_p_O_DFFX1mul_24_1_(injectionVector[83]),
.p_desc259_p_O_DFFX1mul_24_1_(injectionVector[84]),
.p_desc260_p_O_DFFX1mul_24_1_(injectionVector[85]),
.p_desc261_p_O_DFFX1mul_24_1_(injectionVector[86]),
.p_desc262_p_O_DFFX1mul_24_1_(injectionVector[87]),
.p_desc263_p_O_DFFX1mul_24_1_(injectionVector[88]),
.p_desc264_p_O_DFFX1mul_24_1_(injectionVector[89]),
.p_desc265_p_O_DFFX1mul_24_1_(injectionVector[90]),
.p_desc266_p_O_DFFX1mul_24_1_(injectionVector[91]),
.p_desc267_p_O_DFFX1mul_24_1_(injectionVector[92]),
.p_desc268_p_O_DFFX1mul_24_1_(injectionVector[93]),
.p_desc269_p_O_DFFX1mul_24_1_(injectionVector[94]),
.p_desc270_p_O_DFFX1mul_24_1_(injectionVector[95]),
.p_desc271_p_O_DFFX1mul_24_1_(injectionVector[96]),
.p_desc272_p_O_DFFX1mul_24_1_(injectionVector[97]),
.p_desc273_p_O_DFFX1mul_24_1_(injectionVector[98]),
.p_desc274_p_O_DFFX1mul_24_1_(injectionVector[99]),
.p_desc275_p_O_DFFX1mul_24_1_(injectionVector[100]),
.p_desc276_p_O_DFFX1mul_24_1_(injectionVector[101]),
.p_desc277_p_O_DFFX1mul_24_1_(injectionVector[102]),
.p_desc278_p_O_DFFX1mul_24_1_(injectionVector[103]),
.p_desc279_p_O_DFFX1mul_24_1_(injectionVector[104]),
.p_desc280_p_O_DFFX1mul_24_1_(injectionVector[105]),
.p_desc281_p_O_DFFX1mul_24_1_(injectionVector[106]),
.p_desc282_p_O_DFFX1mul_24_1_(injectionVector[107]),
.p_desc283_p_O_DFFX1mul_24_1_(injectionVector[108]),
.p_desc284_p_O_DFFX1mul_24_1_(injectionVector[109]),
.p_desc285_p_O_DFFX1mul_24_1_(injectionVector[110]),
.p_desc286_p_O_DFFX1mul_24_1_(injectionVector[111]),
.p_desc287_p_O_DFFX1mul_24_1_(injectionVector[112]),
.p_desc288_p_O_DFFX1mul_24_1_(injectionVector[113]),
.p_desc289_p_O_DFFX1mul_24_1_(injectionVector[114]),
.p_desc290_p_O_DFFX1mul_24_1_(injectionVector[115]),
.p_desc291_p_O_DFFX1mul_24_1_(injectionVector[116]),
.p_desc292_p_O_DFFX1mul_24_1_(injectionVector[117]),
.p_desc293_p_O_DFFX1mul_24_1_(injectionVector[118]),
.p_desc294_p_O_DFFX1mul_24_1_(injectionVector[119]),
.p_desc295_p_O_DFFX1mul_24_1_(injectionVector[120]),
.p_desc296_p_O_DFFX1mul_24_1_(injectionVector[121]),
.p_desc297_p_O_DFFX1mul_24_1_(injectionVector[122]),
.p_desc298_p_O_DFFX1mul_24_1_(injectionVector[123]),
.p_desc299_p_O_DFFX1mul_24_1_(injectionVector[124]),
.p_desc300_p_O_DFFX1mul_24_1_(injectionVector[125]),
.p_desc301_p_O_DFFX1mul_24_1_(injectionVector[126]),
.p_desc302_p_O_DFFX1mul_24_1_(injectionVector[127]),
.p_desc303_p_O_DFFX1mul_24_1_(injectionVector[128]),
.p_desc304_p_O_DFFX1mul_24_1_(injectionVector[129]),
.p_desc305_p_O_DFFX1mul_24_1_(injectionVector[130]),
.p_desc306_p_O_DFFX1mul_24_1_(injectionVector[131]),
.p_desc307_p_O_DFFX1mul_24_1_(injectionVector[132]),
.p_desc308_p_O_DFFX1mul_24_1_(injectionVector[133]),
.p_desc309_p_O_DFFX1mul_24_1_(injectionVector[134]),
.p_desc310_p_O_DFFX1mul_24_1_(injectionVector[135]),
.p_desc311_p_O_DFFX1mul_24_1_(injectionVector[136]),
.p_desc312_p_O_DFFX1mul_24_1_(injectionVector[137]),
.p_desc313_p_O_DFFX1mul_24_1_(injectionVector[138]),
.p_desc314_p_O_DFFX1mul_24_1_(injectionVector[139]),
.p_desc315_p_O_DFFX1mul_24_1_(injectionVector[140]),
.p_desc316_p_O_DFFX1mul_24_1_(injectionVector[141]),
.p_desc317_p_O_DFFX1mul_24_1_(injectionVector[142]),
.p_desc318_p_O_DFFX1mul_24_1_(injectionVector[143]),
.p_desc319_p_O_DFFX1mul_24_1_(injectionVector[144]),
.p_desc320_p_O_DFFX1mul_24_1_(injectionVector[145]),
.p_desc321_p_O_DFFX1mul_24_1_(injectionVector[146]),
.p_desc322_p_O_DFFX1mul_24_1_(injectionVector[147]),
.p_desc323_p_O_DFFX1mul_24_1_(injectionVector[148]),
.p_desc324_p_O_DFFX1mul_24_1_(injectionVector[149]),
.p_desc325_p_O_DFFX1mul_24_1_(injectionVector[150]),
.p_desc326_p_O_DFFX1mul_24_1_(injectionVector[151]),
.p_desc327_p_O_DFFX1mul_24_1_(injectionVector[152]),
.p_desc328_p_O_DFFX1mul_24_1_(injectionVector[153]),
.p_desc329_p_O_DFFX1mul_24_1_(injectionVector[154]),
.p_desc330_p_O_DFFX1mul_24_1_(injectionVector[155]),
.p_desc331_p_O_DFFX1mul_24_1_(injectionVector[156]),
.p_desc332_p_O_DFFX1mul_24_1_(injectionVector[157]),
.p_desc333_p_O_DFFX1mul_24_1_(injectionVector[158]),
.p_desc334_p_O_DFFX1mul_24_1_(injectionVector[159]),
.p_desc335_p_O_DFFX1mul_24_1_(injectionVector[160]),
.p_desc336_p_O_DFFX1mul_24_1_(injectionVector[161]),
.p_desc337_p_O_DFFX1mul_24_1_(injectionVector[162]),
.p_desc338_p_O_DFFX1mul_24_1_(injectionVector[163]),
.p_desc339_p_O_DFFX1mul_24_1_(injectionVector[164]),
.p_desc340_p_O_DFFX1mul_24_1_(injectionVector[165]),
.p_desc341_p_O_DFFX1mul_24_1_(injectionVector[166]),
.p_desc342_p_O_DFFX1mul_24_1_(injectionVector[167]),
.p_desc343_p_O_DFFX1mul_24_1_(injectionVector[168]),
.p_desc344_p_O_DFFX1mul_24_1_(injectionVector[169]),
.p_desc345_p_O_DFFX1mul_24_1_(injectionVector[170]),
.p_desc346_p_O_DFFX1mul_24_1_(injectionVector[171]),
.p_desc347_p_O_DFFX1mul_24_1_(injectionVector[172]),
.p_desc348_p_O_DFFX1mul_24_1_(injectionVector[173]),
.p_desc349_p_O_DFFX1mul_24_1_(injectionVector[174]),
.p_desc350_p_O_DFFX1mul_24_1_(injectionVector[175]),
.p_desc351_p_O_DFFX1mul_24_1_(injectionVector[176]),
.p_desc352_p_O_DFFX1mul_24_1_(injectionVector[177]),
.p_desc353_p_O_DFFX1mul_24_1_(injectionVector[178]),
.p_desc354_p_O_DFFX1mul_24_1_(injectionVector[179]),
.p_desc355_p_O_DFFX1mul_24_1_(injectionVector[180]),
.p_desc356_p_O_DFFX1mul_24_1_(injectionVector[181]),
.p_desc357_p_O_DFFX1mul_24_1_(injectionVector[182]),
.p_desc358_p_O_DFFX1mul_24_1_(injectionVector[183]),
.p_desc359_p_O_DFFX1mul_24_1_(injectionVector[184]),
.p_desc360_p_O_DFFX1mul_24_1_(injectionVector[185]),
.p_desc361_p_O_DFFX1mul_24_1_(injectionVector[186]),
.p_desc362_p_O_DFFX1mul_24_1_(injectionVector[187]),
.p_desc363_p_O_DFFX1mul_24_1_(injectionVector[188]),
.p_desc364_p_O_DFFX1mul_24_1_(injectionVector[189]),
.p_desc365_p_O_DFFX1mul_24_1_(injectionVector[190]),
.p_desc366_p_O_DFFX1mul_24_1_(injectionVector[191]),
.p_desc367_p_O_DFFX1mul_24_1_(injectionVector[192]),
.p_desc368_p_O_DFFX1mul_24_1_(injectionVector[193]),
.p_desc369_p_O_DFFX1mul_24_1_(injectionVector[194]),
.p_desc370_p_O_DFFX1mul_24_1_(injectionVector[195]),
.p_desc371_p_O_DFFX1mul_24_1_(injectionVector[196]),
.p_desc372_p_O_DFFX1mul_24_1_(injectionVector[197]),
.p_desc373_p_O_DFFX1mul_24_1_(injectionVector[198]),
.p_desc374_p_O_DFFX1mul_24_1_(injectionVector[199]),
.p_desc375_p_O_DFFX1mul_24_1_(injectionVector[200]),
.p_desc376_p_O_DFFX1mul_24_1_(injectionVector[201]),
.p_desc377_p_O_DFFX1mul_24_1_(injectionVector[202]),
.p_desc378_p_O_DFFX1mul_24_1_(injectionVector[203]),
.p_desc379_p_O_DFFX1mul_24_1_(injectionVector[204]),
.p_desc380_p_O_DFFX1mul_24_1_(injectionVector[205]),
.p_desc381_p_O_DFFX1mul_24_1_(injectionVector[206]),
.p_desc382_p_O_DFFX1mul_24_1_(injectionVector[207]),
.p_desc383_p_O_DFFX1mul_24_1_(injectionVector[208]),
.p_desc384_p_O_DFFX1mul_24_1_(injectionVector[209]),
.p_desc385_p_O_DFFX1mul_24_1_(injectionVector[210]),
.p_desc386_p_O_DFFX1mul_24_1_(injectionVector[211]),
.p_desc387_p_O_DFFX1mul_24_1_(injectionVector[212]),
.p_desc388_p_O_DFFX1mul_24_1_(injectionVector[213]),
.p_desc389_p_O_DFFX1mul_24_1_(injectionVector[214]),
.p_desc390_p_O_DFFX1mul_24_1_(injectionVector[215]),
.p_desc391_p_O_DFFX1mul_24_1_(injectionVector[216]),
.p_desc392_p_O_DFFX1mul_24_1_(injectionVector[217]),
.p_desc393_p_O_DFFX1mul_24_1_(injectionVector[218]),
.p_desc394_p_O_DFFX1mul_24_1_(injectionVector[219]),
.p_desc395_p_O_DFFX1mul_24_1_(injectionVector[220]),
.p_desc396_p_O_DFFX1mul_24_1_(injectionVector[221]),
.p_desc397_p_O_DFFX1mul_24_1_(injectionVector[222]),
.p_desc398_p_O_DFFX1mul_24_1_(injectionVector[223]),
.p_desc399_p_O_DFFX1mul_24_1_(injectionVector[224]),
.p_desc400_p_O_DFFX1mul_24_1_(injectionVector[225]),
.p_desc401_p_O_DFFX1mul_24_1_(injectionVector[226]),
.p_desc402_p_O_DFFX1mul_24_1_(injectionVector[227]),
.p_desc403_p_O_DFFX1mul_24_1_(injectionVector[228]),
.p_desc404_p_O_DFFX1mul_24_1_(injectionVector[229]),
.p_desc405_p_O_DFFX1mul_24_1_(injectionVector[230]),
.p_desc406_p_O_DFFX1mul_24_1_(injectionVector[231]),
.p_desc407_p_O_DFFX1mul_24_1_(injectionVector[232]),
.p_desc408_p_O_DFFX1mul_24_1_(injectionVector[233]),
.p_desc409_p_O_DFFX1mul_24_1_(injectionVector[234]),
.p_desc410_p_O_DFFX1mul_24_1_(injectionVector[235]),
.p_desc411_p_O_DFFX1mul_24_1_(injectionVector[236]),
.p_desc412_p_O_DFFX1mul_24_1_(injectionVector[237]),
.p_desc413_p_O_DFFX1mul_24_1_(injectionVector[238]),
.p_desc414_p_O_DFFX1mul_24_1_(injectionVector[239]),
.p_desc415_p_O_DFFX1mul_24_1_(injectionVector[240]),
.p_desc416_p_O_DFFX1mul_24_1_(injectionVector[241]),
.p_desc417_p_O_DFFX1mul_24_1_(injectionVector[242]),
.p_desc418_p_O_DFFX1mul_24_1_(injectionVector[243]),
.p_desc419_p_O_DFFX1mul_24_1_(injectionVector[244]),
.p_desc420_p_O_DFFX1mul_24_1_(injectionVector[245]),
.p_desc421_p_O_DFFX1mul_24_1_(injectionVector[246]),
.p_desc422_p_O_DFFX1mul_24_1_(injectionVector[247]),
.p_desc423_p_O_DFFX1mul_24_1_(injectionVector[248]),
.p_desc424_p_O_DFFX1mul_24_1_(injectionVector[249]),
.p_desc425_p_O_DFFX1mul_24_1_(injectionVector[250]),
.p_desc426_p_O_DFFX1mul_24_1_(injectionVector[251]),
.p_desc427_p_O_DFFX1mul_24_1_(injectionVector[252]),
.p_desc428_p_O_DFFX1mul_24_1_(injectionVector[253]),
.p_desc429_p_O_DFFX1mul_24_1_(injectionVector[254]),
.p_desc430_p_O_DFFX1mul_24_1_(injectionVector[255]),
.p_desc431_p_O_DFFX1mul_24_1_(injectionVector[256]),
.p_desc432_p_O_DFFX1mul_24_1_(injectionVector[257]),
.p_desc433_p_O_DFFX1mul_24_1_(injectionVector[258]),
.p_desc434_p_O_DFFX1mul_24_1_(injectionVector[259]),
.p_desc435_p_O_DFFX1mul_24_1_(injectionVector[260]),
.p_desc436_p_O_DFFX1mul_24_1_(injectionVector[261]),
.p_desc437_p_O_DFFX1mul_24_1_(injectionVector[262]),
.p_desc438_p_O_DFFX1mul_24_1_(injectionVector[263]),
.p_desc439_p_O_DFFX1mul_24_1_(injectionVector[264]),
.p_desc440_p_O_DFFX1mul_24_1_(injectionVector[265]),
.p_desc441_p_O_DFFX1mul_24_1_(injectionVector[266]),
.p_desc442_p_O_DFFX1mul_24_1_(injectionVector[267]),
.p_desc443_p_O_DFFX1mul_24_1_(injectionVector[268]),
.p_desc444_p_O_DFFX1mul_24_1_(injectionVector[269]),
.p_desc445_p_O_DFFX1mul_24_1_(injectionVector[270]),
.p_desc446_p_O_DFFX1mul_24_1_(injectionVector[271]),
.p_desc447_p_O_DFFX1mul_24_1_(injectionVector[272]),
.p_desc448_p_O_DFFX1mul_24_1_(injectionVector[273]),
.p_desc449_p_O_DFFX1mul_24_1_(injectionVector[274]),
.p_desc450_p_O_DFFX1mul_24_1_(injectionVector[275]),
.p_desc451_p_O_DFFX1mul_24_1_(injectionVector[276]),
.p_desc452_p_O_DFFX1mul_24_1_(injectionVector[277]),
.p_desc453_p_O_DFFX1mul_24_1_(injectionVector[278]),
.p_desc454_p_O_DFFX1mul_24_1_(injectionVector[279]),
.p_desc455_p_O_DFFX1mul_24_1_(injectionVector[280]),
.p_desc456_p_O_DFFX1mul_24_1_(injectionVector[281]),
.p_desc457_p_O_DFFX1mul_24_1_(injectionVector[282]),
.p_desc458_p_O_DFFX1mul_24_1_(injectionVector[283]),
.p_desc459_p_O_DFFX1mul_24_1_(injectionVector[284]),
.p_desc460_p_O_DFFX1mul_24_1_(injectionVector[285]),
.p_desc461_p_O_DFFX1mul_24_1_(injectionVector[286]),
.p_desc462_p_O_DFFX1mul_24_1_(injectionVector[287]),
.p_desc463_p_O_DFFX1mul_24_1_(injectionVector[288]),
.p_desc464_p_O_DFFX1mul_24_1_(injectionVector[289]),
.p_desc465_p_O_DFFX1mul_24_1_(injectionVector[290]),
.p_desc466_p_O_DFFX1mul_24_1_(injectionVector[291]),
.p_desc467_p_O_DFFX1mul_24_1_(injectionVector[292]),
.p_desc468_p_O_DFFX1mul_24_1_(injectionVector[293]),
.p_desc469_p_O_DFFX1mul_24_1_(injectionVector[294]),
.p_desc470_p_O_DFFX1mul_24_1_(injectionVector[295]),
.p_desc471_p_O_DFFX1mul_24_1_(injectionVector[296]),
.p_desc472_p_O_DFFX1mul_24_1_(injectionVector[297]),
.p_desc473_p_O_DFFX1mul_24_1_(injectionVector[298]),
.p_desc474_p_O_DFFX1mul_24_1_(injectionVector[299]),
.p_desc475_p_O_DFFX1mul_24_1_(injectionVector[300]),
.p_desc476_p_O_DFFX1mul_24_1_(injectionVector[301]),
.p_desc477_p_O_DFFX1mul_24_1_(injectionVector[302]),
.p_desc478_p_O_DFFX1mul_24_1_(injectionVector[303]),
.p_desc479_p_O_DFFX1mul_24_1_(injectionVector[304]),
.p_desc480_p_O_DFFX1mul_24_1_(injectionVector[305]),
.p_desc481_p_O_DFFX1mul_24_1_(injectionVector[306]),
.p_desc482_p_O_DFFX1mul_24_1_(injectionVector[307]),
.p_desc483_p_O_DFFX1mul_24_1_(injectionVector[308]),
.p_desc484_p_O_DFFX1mul_24_1_(injectionVector[309]),
.p_desc485_p_O_DFFX1mul_24_1_(injectionVector[310]),
.p_desc486_p_O_DFFX1mul_24_1_(injectionVector[311]),
.p_desc487_p_O_DFFX1mul_24_1_(injectionVector[312]),
.p_desc488_p_O_DFFX1mul_24_1_(injectionVector[313]),
.p_desc489_p_O_DFFX1mul_24_1_(injectionVector[314]),
.p_desc490_p_O_DFFX1mul_24_1_(injectionVector[315]),
.p_desc491_p_O_DFFX1mul_24_1_(injectionVector[316]),
.p_desc492_p_O_DFFX1mul_24_1_(injectionVector[317]),
.p_desc493_p_O_DFFX1mul_24_1_(injectionVector[318]),
.p_desc494_p_O_DFFX1mul_24_1_(injectionVector[319]),
.p_desc495_p_O_DFFX1mul_24_1_(injectionVector[320]),
.p_desc496_p_O_DFFX1mul_24_1_(injectionVector[321]),
.p_desc497_p_O_DFFX1mul_24_1_(injectionVector[322]),
.p_desc498_p_O_DFFX1mul_24_1_(injectionVector[323]),
.p_desc499_p_O_DFFX1mul_24_1_(injectionVector[324]),
.p_desc500_p_O_DFFX1mul_24_1_(injectionVector[325]),
.p_desc501_p_O_DFFX1mul_24_1_(injectionVector[326]),
.p_desc502_p_O_DFFX1mul_24_1_(injectionVector[327]),
.p_desc503_p_O_DFFX1mul_24_1_(injectionVector[328]),
.p_desc504_p_O_DFFX1mul_24_1_(injectionVector[329]),
.p_desc505_p_O_DFFX1mul_24_1_(injectionVector[330]),
.p_desc506_p_O_DFFX1mul_24_1_(injectionVector[331]),
.p_desc507_p_O_DFFX1mul_24_1_(injectionVector[332]),
.p_desc508_p_O_DFFX1mul_24_1_(injectionVector[333]),
.p_desc509_p_O_DFFX1mul_24_1_(injectionVector[334]),
.p_desc510_p_O_DFFX1mul_24_1_(injectionVector[335]),
.p_desc511_p_O_DFFX1mul_24_1_(injectionVector[336]),
.p_desc512_p_O_DFFX1mul_24_1_(injectionVector[337]),
.p_desc513_p_O_DFFX1mul_24_1_(injectionVector[338]),
.p_desc514_p_O_DFFX1mul_24_1_(injectionVector[339]),
.p_desc515_p_O_DFFX1mul_24_1_(injectionVector[340]),
.p_desc516_p_O_DFFX1mul_24_1_(injectionVector[341]),
.p_desc517_p_O_DFFX1mul_24_1_(injectionVector[342]),
.p_desc518_p_O_DFFX1mul_24_1_(injectionVector[343]),
.p_desc519_p_O_DFFX1mul_24_1_(injectionVector[344]),
.p_desc520_p_O_DFFX1mul_24_1_(injectionVector[345]),
.p_desc521_p_O_DFFX1mul_24_1_(injectionVector[346]),
.p_desc522_p_O_DFFX1mul_24_1_(injectionVector[347]),
.p_desc523_p_O_DFFX1mul_24_1_(injectionVector[348]),
.p_desc524_p_O_DFFX1mul_24_1_(injectionVector[349]),
.p_desc525_p_O_DFFX1mul_24_1_(injectionVector[350]),
.p_desc526_p_O_DFFX1mul_24_1_(injectionVector[351]),
.p_desc527_p_O_DFFX1mul_24_1_(injectionVector[352]),
.p_desc528_p_O_DFFX1mul_24_1_(injectionVector[353]),
.p_desc678_p_O_DFFX1post_norm_mul_1_(injectionVector[354]),
.p_desc679_p_O_DFFX1post_norm_mul_1_(injectionVector[355]),
.p_desc680_p_O_DFFX1post_norm_mul_1_(injectionVector[356]),
.p_desc681_p_O_DFFX1post_norm_mul_1_(injectionVector[357]),
.p_desc682_p_O_DFFX1post_norm_mul_1_(injectionVector[358]),
.p_desc683_p_O_DFFX1post_norm_mul_1_(injectionVector[359]),
.p_desc684_p_O_DFFX1post_norm_mul_1_(injectionVector[360]),
.p_desc685_p_O_DFFX1post_norm_mul_1_(injectionVector[361]),
.p_desc686_p_O_DFFX1post_norm_mul_1_(injectionVector[362]),
.p_desc687_p_O_DFFX1post_norm_mul_1_(injectionVector[363]),
.p_desc688_p_O_DFFX1post_norm_mul_1_(injectionVector[364]),
.p_desc689_p_O_DFFX1post_norm_mul_1_(injectionVector[365]),
.p_desc690_p_O_DFFX1post_norm_mul_1_(injectionVector[366]),
.p_desc691_p_O_DFFX1post_norm_mul_1_(injectionVector[367]),
.p_desc692_p_O_DFFX1post_norm_mul_1_(injectionVector[368]),
.p_desc693_p_O_DFFX1post_norm_mul_1_(injectionVector[369]),
.p_desc694_p_O_DFFX1post_norm_mul_1_(injectionVector[370]),
.p_desc695_p_O_DFFX1post_norm_mul_1_(injectionVector[371]),
.p_desc696_p_O_DFFX1post_norm_mul_1_(injectionVector[372]),
.p_desc697_p_O_DFFX1post_norm_mul_1_(injectionVector[373]),
.p_desc698_p_O_DFFX1post_norm_mul_1_(injectionVector[374]),
.p_desc699_p_O_DFFX1post_norm_mul_1_(injectionVector[375]),
.p_desc700_p_O_DFFX1post_norm_mul_1_(injectionVector[376]),
.p_desc701_p_O_DFFX1post_norm_mul_1_(injectionVector[377]),
.p_desc702_p_O_DFFX1post_norm_mul_1_(injectionVector[378]),
.p_desc703_p_O_DFFX1post_norm_mul_1_(injectionVector[379]),
.p_desc704_p_O_DFFX1post_norm_mul_1_(injectionVector[380]),
.p_desc705_p_O_DFFX1post_norm_mul_1_(injectionVector[381]),
.p_desc706_p_O_DFFX1post_norm_mul_1_(injectionVector[382]),
.p_desc707_p_O_DFFX1post_norm_mul_1_(injectionVector[383]),
.p_desc708_p_O_DFFX1post_norm_mul_1_(injectionVector[384]),
.p_desc709_p_O_DFFX1post_norm_mul_1_(injectionVector[385]),
.p_desc710_p_O_DFFX1post_norm_mul_1_(injectionVector[386]),
.p_desc711_p_O_DFFX1post_norm_mul_1_(injectionVector[387]),
.p_desc712_p_O_DFFX1post_norm_mul_1_(injectionVector[388]),
.p_desc713_p_O_DFFX1post_norm_mul_1_(injectionVector[389]),
.p_desc714_p_O_DFFX1post_norm_mul_1_(injectionVector[390]),
.p_desc715_p_O_DFFX1post_norm_mul_1_(injectionVector[391]),
.p_desc716_p_O_DFFX1post_norm_mul_1_(injectionVector[392]),
.p_desc717_p_O_DFFX1post_norm_mul_1_(injectionVector[393]),
.p_desc718_p_O_DFFX1post_norm_mul_1_(injectionVector[394]),
.p_desc719_p_O_DFFX1post_norm_mul_1_(injectionVector[395]),
.p_desc720_p_O_DFFX1post_norm_mul_1_(injectionVector[396]),
.p_desc721_p_O_DFFX1post_norm_mul_1_(injectionVector[397]),
.p_desc722_p_O_DFFX1post_norm_mul_1_(injectionVector[398]),
.p_desc723_p_O_DFFX1post_norm_mul_1_(injectionVector[399]),
.p_desc724_p_O_DFFX1post_norm_mul_1_(injectionVector[400]),
.p_desc725_p_O_DFFX1post_norm_mul_1_(injectionVector[401]),
.p_desc726_p_O_DFFX1post_norm_mul_1_(injectionVector[402]),
.p_desc727_p_O_DFFX1post_norm_mul_1_(injectionVector[403]),
.p_desc728_p_O_DFFX1post_norm_mul_1_(injectionVector[404]),
.p_desc729_p_O_DFFX1post_norm_mul_1_(injectionVector[405]),
.p_desc730_p_O_DFFX1post_norm_mul_1_(injectionVector[406]),
.p_desc731_p_O_DFFX1post_norm_mul_1_(injectionVector[407]),
.p_desc732_p_O_DFFX1post_norm_mul_1_(injectionVector[408]),
.p_desc733_p_O_DFFX1post_norm_mul_1_(injectionVector[409]),
.p_desc734_p_O_DFFX1post_norm_mul_1_(injectionVector[410]),
.p_desc735_p_O_DFFX1post_norm_mul_1_(injectionVector[411]),
.p_desc736_p_O_DFFX1post_norm_mul_1_(injectionVector[412]),
.p_desc737_p_O_DFFX1post_norm_mul_1_(injectionVector[413]),
.p_desc738_p_O_DFFX1post_norm_mul_1_(injectionVector[414]),
.p_desc739_p_O_DFFX1post_norm_mul_1_(injectionVector[415]),
.p_desc740_p_O_DFFX1post_norm_mul_1_(injectionVector[416]),
.p_desc741_p_O_DFFX1post_norm_mul_1_(injectionVector[417]),
.p_desc742_p_O_DFFX1post_norm_mul_1_(injectionVector[418]),
.p_desc743_p_O_DFFX1post_norm_mul_1_(injectionVector[419]),
.p_desc744_p_O_DFFX1post_norm_mul_1_(injectionVector[420]),
.p_desc745_p_O_DFFX1post_norm_mul_1_(injectionVector[421]),
.p_desc746_p_O_DFFX1post_norm_mul_1_(injectionVector[422]),
.p_desc747_p_O_DFFX1post_norm_mul_1_(injectionVector[423]),
.p_desc748_p_O_DFFX1post_norm_mul_1_(injectionVector[424]),
.p_desc749_p_O_DFFX1post_norm_mul_1_(injectionVector[425]),
.p_desc750_p_O_DFFX1post_norm_mul_1_(injectionVector[426]),
.p_desc751_p_O_DFFX1post_norm_mul_1_(injectionVector[427]),
.p_desc752_p_O_DFFX1post_norm_mul_1_(injectionVector[428]),
.p_desc753_p_O_DFFX1post_norm_mul_1_(injectionVector[429]),
.p_desc754_p_O_DFFX1post_norm_mul_1_(injectionVector[430]),
.p_desc755_p_O_DFFX1post_norm_mul_1_(injectionVector[431]),
.p_desc756_p_O_DFFX1post_norm_mul_1_(injectionVector[432]),
.p_desc757_p_O_DFFX1post_norm_mul_1_(injectionVector[433]),
.p_desc758_p_O_DFFX1post_norm_mul_1_(injectionVector[434]),
.p_desc759_p_O_DFFX1post_norm_mul_1_(injectionVector[435]),
.p_desc760_p_O_DFFX1post_norm_mul_1_(injectionVector[436]),
.p_desc761_p_O_DFFX1post_norm_mul_1_(injectionVector[437]),
.p_desc762_p_O_DFFX1post_norm_mul_1_(injectionVector[438]),
.p_desc763_p_O_DFFX1post_norm_mul_1_(injectionVector[439]),
.p_desc764_p_O_DFFX1post_norm_mul_1_(injectionVector[440]),
.p_desc765_p_O_DFFX1post_norm_mul_1_(injectionVector[441]),
.p_desc766_p_O_DFFX1post_norm_mul_1_(injectionVector[442]),
.p_desc767_p_O_DFFX1post_norm_mul_1_(injectionVector[443]),
.p_desc768_p_O_DFFX1post_norm_mul_1_(injectionVector[444]),
.p_desc769_p_O_DFFX1post_norm_mul_1_(injectionVector[445]),
.p_desc770_p_O_DFFX1post_norm_mul_1_(injectionVector[446]),
.p_desc771_p_O_DFFX1post_norm_mul_1_(injectionVector[447]),
.p_desc772_p_O_DFFX1post_norm_mul_1_(injectionVector[448]),
.p_desc773_p_O_DFFX1post_norm_mul_1_(injectionVector[449]),
.p_desc774_p_O_DFFX1post_norm_mul_1_(injectionVector[450]),
.p_desc775_p_O_DFFX1post_norm_mul_1_(injectionVector[451]),
.p_desc776_p_O_DFFX1post_norm_mul_1_(injectionVector[452]),
.p_desc777_p_O_DFFX1post_norm_mul_1_(injectionVector[453]),
.p_desc778_p_O_DFFX1post_norm_mul_1_(injectionVector[454]),
.p_desc779_p_O_DFFX1post_norm_mul_1_(injectionVector[455]),
.p_desc780_p_O_DFFX1post_norm_mul_1_(injectionVector[456]),
.p_desc781_p_O_DFFX1post_norm_mul_1_(injectionVector[457]),
.p_desc782_p_O_DFFX1post_norm_mul_1_(injectionVector[458]),
.p_desc783_p_O_DFFX1post_norm_mul_1_(injectionVector[459]),
.p_desc784_p_O_DFFX1post_norm_mul_1_(injectionVector[460]),
.p_desc785_p_O_DFFX1post_norm_mul_1_(injectionVector[461]),
.p_desc786_p_O_DFFX1post_norm_mul_1_(injectionVector[462]),
.p_desc787_p_O_DFFX1post_norm_mul_1_(injectionVector[463]),
.p_desc788_p_O_DFFX1post_norm_mul_1_(injectionVector[464]),
.p_desc789_p_O_DFFX1post_norm_mul_1_(injectionVector[465]),
.p_desc790_p_O_DFFX1post_norm_mul_1_(injectionVector[466]),
.p_desc791_p_O_DFFX1post_norm_mul_1_(injectionVector[467]),
.p_desc792_p_O_DFFX1post_norm_mul_1_(injectionVector[468]),
.p_desc793_p_O_DFFX1post_norm_mul_1_(injectionVector[469]),
.p_desc794_p_O_DFFX1post_norm_mul_1_(injectionVector[470]),
.p_desc795_p_O_DFFX1post_norm_mul_1_(injectionVector[471]),
.p_desc796_p_O_DFFX1post_norm_mul_1_(injectionVector[472]),
.p_desc797_p_O_DFFX1post_norm_mul_1_(injectionVector[473]),
.p_desc798_p_O_DFFX1post_norm_mul_1_(injectionVector[474]),
.p_desc799_p_O_DFFX1post_norm_mul_1_(injectionVector[475]),
.p_desc800_p_O_DFFX1post_norm_mul_1_(injectionVector[476]),
.p_desc801_p_O_DFFX1post_norm_mul_1_(injectionVector[477]),
.p_desc802_p_O_DFFX1post_norm_mul_1_(injectionVector[478]),
.p_desc803_p_O_DFFX1post_norm_mul_1_(injectionVector[479]),
.p_desc804_p_O_DFFX1post_norm_mul_1_(injectionVector[480]),
.p_desc805_p_O_DFFX1post_norm_mul_1_(injectionVector[481]),
.p_desc806_p_O_DFFX1post_norm_mul_1_(injectionVector[482]),
.p_desc807_p_O_DFFX1post_norm_mul_1_(injectionVector[483]),
.p_desc808_p_O_DFFX1post_norm_mul_1_(injectionVector[484]),
.p_desc809_p_O_DFFX1post_norm_mul_1_(injectionVector[485]),
.p_desc810_p_O_DFFX1post_norm_mul_1_(injectionVector[486]),
.p_desc811_p_O_DFFX1post_norm_mul_1_(injectionVector[487]),
.p_desc812_p_O_DFFX1post_norm_mul_1_(injectionVector[488]),
.p_desc813_p_O_DFFX1post_norm_mul_1_(injectionVector[489]),
.p_s_sign_i_reg_p_O_DFFX1post_norm_mul_1_(injectionVector[490]),
.p_desc814_p_O_DFFX1post_norm_mul_1_(injectionVector[491]),
.p_desc815_p_O_DFFX1post_norm_mul_1_(injectionVector[492]),
.p_desc816_p_O_DFFX1post_norm_mul_1_(injectionVector[493]),
.p_desc817_p_O_DFFX1post_norm_mul_1_(injectionVector[494]),
.p_desc818_p_O_DFFX1post_norm_mul_1_(injectionVector[495]),
.p_desc819_p_O_DFFX1post_norm_mul_1_(injectionVector[496]),
.p_desc820_p_O_DFFX1post_norm_mul_1_(injectionVector[497]),
.p_desc821_p_O_DFFX1post_norm_mul_1_(injectionVector[498]),
.p_desc822_p_O_DFFX1post_norm_mul_1_(injectionVector[499]),
.p_desc823_p_O_DFFX1post_norm_mul_1_(injectionVector[500]),
.p_desc824_p_O_DFFX1post_norm_mul_1_(injectionVector[501]),
.p_desc825_p_O_DFFX1post_norm_mul_1_(injectionVector[502]),
.p_desc826_p_O_DFFX1post_norm_mul_1_(injectionVector[503]),
.p_desc827_p_O_DFFX1post_norm_mul_1_(injectionVector[504]),
.p_desc828_p_O_DFFX1post_norm_mul_1_(injectionVector[505]),
.p_desc829_p_O_DFFX1post_norm_mul_1_(injectionVector[506]),
.p_desc830_p_O_DFFX1post_norm_mul_1_(injectionVector[507]),
.p_desc831_p_O_DFFX1post_norm_mul_1_(injectionVector[508]),
.p_desc832_p_O_DFFX1post_norm_mul_1_(injectionVector[509]),
.p_desc833_p_O_DFFX1post_norm_mul_1_(injectionVector[510]),
.p_desc834_p_O_DFFX1post_norm_mul_1_(injectionVector[511]),
.p_desc835_p_O_DFFX1post_norm_mul_1_(injectionVector[512]),
.p_desc836_p_O_DFFX1post_norm_mul_1_(injectionVector[513]),
.p_desc837_p_O_DFFX1post_norm_mul_1_(injectionVector[514]),
.p_desc838_p_O_DFFX1post_norm_mul_1_(injectionVector[515]),
.p_desc839_p_O_DFFX1post_norm_mul_1_(injectionVector[516]),
.p_desc840_p_O_DFFX1post_norm_mul_1_(injectionVector[517]),
.p_desc841_p_O_DFFX1post_norm_mul_1_(injectionVector[518]),
.p_desc842_p_O_DFFX1post_norm_mul_1_(injectionVector[519]),
.p_desc843_p_O_DFFX1post_norm_mul_1_(injectionVector[520]),
.p_desc844_p_O_DFFX1post_norm_mul_1_(injectionVector[521]),
.p_desc845_p_O_DFFX1post_norm_mul_1_(injectionVector[522]),
.p_desc846_p_O_DFFX1post_norm_mul_1_(injectionVector[523]),
.p_desc847_p_O_DFFX1post_norm_mul_1_(injectionVector[524]),
.p_desc848_p_O_DFFX1post_norm_mul_1_(injectionVector[525]),
.p_desc849_p_O_DFFX1post_norm_mul_1_(injectionVector[526]),
.p_desc850_p_O_DFFX1post_norm_mul_1_(injectionVector[527]),
.p_desc851_p_O_DFFX1post_norm_mul_1_(injectionVector[528]),
.p_desc852_p_O_DFFX1post_norm_mul_1_(injectionVector[529]),
.p_desc853_p_O_DFFX1post_norm_mul_1_(injectionVector[530]),
.p_desc854_p_O_DFFX1post_norm_mul_1_(injectionVector[531]),
.p_desc855_p_O_DFFX1post_norm_mul_1_(injectionVector[532]),
.p_desc856_p_O_DFFX1post_norm_mul_1_(injectionVector[533]),
.p_desc857_p_O_DFFX1post_norm_mul_1_(injectionVector[534]),
.p_desc858_p_O_DFFX1post_norm_mul_1_(injectionVector[535]),
.p_desc859_p_O_DFFX1post_norm_mul_1_(injectionVector[536]),
.p_desc860_p_O_DFFX1post_norm_mul_1_(injectionVector[537]),
.p_desc861_p_O_DFFX1post_norm_mul_1_(injectionVector[538]),
.p_desc862_p_O_DFFX1post_norm_mul_1_(injectionVector[539]),
.p_desc863_p_O_DFFX1post_norm_mul_1_(injectionVector[540]),
.p_desc864_p_O_DFFX1post_norm_mul_1_(injectionVector[541]),
.p_desc865_p_O_DFFX1post_norm_mul_1_(injectionVector[542]),
.p_desc866_p_O_DFFX1post_norm_mul_1_(injectionVector[543]),
.p_desc867_p_O_DFFX1post_norm_mul_1_(injectionVector[544]),
.p_desc868_p_O_DFFX1post_norm_mul_1_(injectionVector[545]),
.p_desc869_p_O_DFFX1post_norm_mul_1_(injectionVector[546]),
.p_desc870_p_O_DFFX1post_norm_mul_1_(injectionVector[547]),
.p_desc871_p_O_DFFX1post_norm_mul_1_(injectionVector[548]),
.p_desc872_p_O_DFFX1post_norm_mul_1_(injectionVector[549]),
.p_desc873_p_O_DFFX1post_norm_mul_1_(injectionVector[550]),
.p_desc874_p_O_DFFX1post_norm_mul_1_(injectionVector[551]),
.p_desc875_p_O_DFFX1post_norm_mul_1_(injectionVector[552]),
.p_desc876_p_O_DFFX1post_norm_mul_1_(injectionVector[553]),
.p_desc877_p_O_DFFX1post_norm_mul_1_(injectionVector[554]),
.p_desc878_p_O_DFFX1post_norm_mul_1_(injectionVector[555]),
.p_desc879_p_O_DFFX1post_norm_mul_1_(injectionVector[556]),
.p_desc880_p_O_DFFX1post_norm_mul_1_(injectionVector[557]),
.p_desc881_p_O_DFFX1post_norm_mul_1_(injectionVector[558]),
.p_desc882_p_O_DFFX1post_norm_mul_1_(injectionVector[559]),
.p_desc883_p_O_DFFX1post_norm_mul_1_(injectionVector[560]),
.p_desc884_p_O_DFFX1post_norm_mul_1_(injectionVector[561]),
.p_desc885_p_O_DFFX1post_norm_mul_1_(injectionVector[562]),
.p_desc886_p_O_DFFX1post_norm_mul_1_(injectionVector[563]),
.p_desc887_p_O_DFFX1post_norm_mul_1_(injectionVector[564]),
.p_desc888_p_O_DFFX1post_norm_mul_1_(injectionVector[565]),
.p_desc889_p_O_DFFX1post_norm_mul_1_(injectionVector[566]),
.p_desc890_p_O_DFFX1post_norm_mul_1_(injectionVector[567]),
.p_desc891_p_O_DFFX1post_norm_mul_1_(injectionVector[568]),
.p_desc892_p_O_DFFX1post_norm_mul_1_(injectionVector[569]),
.p_desc893_p_O_DFFX1post_norm_mul_1_(injectionVector[570]),
.p_desc894_p_O_DFFX1post_norm_mul_1_(injectionVector[571]),
.p_desc895_p_O_DFFX1post_norm_mul_1_(injectionVector[572]),
.p_desc896_p_O_DFFX1post_norm_mul_1_(injectionVector[573]),
.p_desc897_p_O_DFFX1post_norm_mul_1_(injectionVector[574]),
.p_ine_o_reg_p_O_DFFX1post_norm_mul_1_(injectionVector[575]),
.p_desc898_p_O_DFFX1post_norm_mul_1_(injectionVector[576]),
.p_desc899_p_O_DFFX1post_norm_mul_1_(injectionVector[577]),
.p_desc900_p_O_DFFX1post_norm_mul_1_(injectionVector[578]),
.p_desc901_p_O_DFFX1post_norm_mul_1_(injectionVector[579]),
.p_desc902_p_O_DFFX1post_norm_mul_1_(injectionVector[580]),
.p_desc903_p_O_DFFX1post_norm_mul_1_(injectionVector[581]),
.p_desc904_p_O_DFFX1post_norm_mul_1_(injectionVector[582]),
.p_desc905_p_O_DFFX1post_norm_mul_1_(injectionVector[583]),
.p_desc906_p_O_DFFX1post_norm_mul_1_(injectionVector[584]),
.p_desc907_p_O_DFFX1post_norm_mul_1_(injectionVector[585]),
.p_desc908_p_O_DFFX1post_norm_mul_1_(injectionVector[586]),
.p_desc909_p_O_DFFX1post_norm_mul_1_(injectionVector[587]),
.p_desc910_p_O_DFFX1post_norm_mul_1_(injectionVector[588]),
.p_desc911_p_O_DFFX1post_norm_mul_1_(injectionVector[589]),
.p_desc912_p_O_DFFX1post_norm_mul_1_(injectionVector[590]),
.p_desc913_p_O_DFFX1post_norm_mul_1_(injectionVector[591]),
.p_desc914_p_O_DFFX1post_norm_mul_1_(injectionVector[592]),
.p_desc915_p_O_DFFX1post_norm_mul_1_(injectionVector[593]),
.p_desc916_p_O_DFFX1post_norm_mul_1_(injectionVector[594]),
.p_desc917_p_O_DFFX1post_norm_mul_1_(injectionVector[595]),
.p_desc918_p_O_DFFX1post_norm_mul_1_(injectionVector[596]),
.p_desc919_p_O_DFFX1post_norm_mul_1_(injectionVector[597]),
.p_desc920_p_O_DFFX1post_norm_mul_1_(injectionVector[598]),
.p_desc921_p_O_DFFX1post_norm_mul_1_(injectionVector[599]),
.p_desc922_p_O_DFFX1post_norm_mul_1_(injectionVector[600]),
.p_desc923_p_O_DFFX1post_norm_mul_1_(injectionVector[601]),
.p_desc924_p_O_DFFX1post_norm_mul_1_(injectionVector[602]),
.p_desc925_p_O_DFFX1post_norm_mul_1_(injectionVector[603]),
.p_desc926_p_O_DFFX1post_norm_mul_1_(injectionVector[604]),
.p_desc927_p_O_DFFX1post_norm_mul_1_(injectionVector[605]),
.p_desc928_p_O_DFFX1post_norm_mul_1_(injectionVector[606]),
.p_desc929_p_O_DFFX1post_norm_mul_1_(injectionVector[607]),
.p_desc930_p_O_DFFX1post_norm_mul_1_(injectionVector[608]),
.p_desc931_p_O_DFFX1post_norm_mul_1_(injectionVector[609]),
.p_desc932_p_O_DFFX1post_norm_mul_1_(injectionVector[610]),
.p_desc933_p_O_DFFX1post_norm_mul_1_(injectionVector[611]),
.p_desc934_p_O_DFFX1post_norm_mul_1_(injectionVector[612]),
.p_desc935_p_O_DFFX1post_norm_mul_1_(injectionVector[613]),
.p_desc936_p_O_DFFX1post_norm_mul_1_(injectionVector[614]),
.p_desc937_p_O_DFFX1post_norm_mul_1_(injectionVector[615]),
.p_desc938_p_O_DFFX1post_norm_mul_1_(injectionVector[616]),
.p_desc939_p_O_DFFX1post_norm_mul_1_(injectionVector[617]),
.p_desc940_p_O_DFFX1post_norm_mul_1_(injectionVector[618]),
.p_desc941_p_O_DFFX1post_norm_mul_1_(injectionVector[619]),
.p_desc942_p_O_DFFX1post_norm_mul_1_(injectionVector[620]),
.p_desc943_p_O_DFFX1post_norm_mul_1_(injectionVector[621]),
.p_desc944_p_O_DFFX1post_norm_mul_1_(injectionVector[622]),
.p_desc945_p_O_DFFX1post_norm_mul_1_(injectionVector[623]),
.p_desc946_p_O_DFFX1post_norm_mul_1_(injectionVector[624]),
.p_desc947_p_O_DFFX1post_norm_mul_1_(injectionVector[625]),
.p_desc948_p_O_DFFX1post_norm_mul_1_(injectionVector[626]),
.p_desc949_p_O_DFFX1post_norm_mul_1_(injectionVector[627]),
.p_desc950_p_O_DFFX1post_norm_mul_1_(injectionVector[628]),
.p_desc951_p_O_DFFX1post_norm_mul_1_(injectionVector[629]),
.p_desc952_p_O_DFFX1post_norm_mul_1_(injectionVector[630]));
endmodule