`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[439:0] injectionVector;
fpu_inj toplevel_instance (
.OPA0I(testVector [31:0]),
.OPB0I(testVector [63:32]),
.FPU0OP0I(testVector [66:64]),
.RMODE0I(testVector [68:67]),
.OUTPUT0O(resultVector [31:0]),
.CLK0I(clk),
.START0I(testVector[69]),
.READY0O(resultVector[32]),
.INE0O(resultVector[33]),
.OVERFLOW0O(resultVector[34]),
.UNDERFLOW0O(resultVector[35]),
.DIV0ZERO0O(resultVector[36]),
.INF0O(resultVector[37]),
.ZERO0O(resultVector[38]),
.QNAN0O(resultVector[39]),
.SNAN0O(resultVector[40]),
.p_desc953_p_O_DFFX1pre_norm_div_1_(injectionVector[0]),
.p_desc954_p_O_DFFX1pre_norm_div_1_(injectionVector[1]),
.p_desc955_p_O_DFFX1pre_norm_div_1_(injectionVector[2]),
.p_desc956_p_O_DFFX1pre_norm_div_1_(injectionVector[3]),
.p_desc957_p_O_DFFX1pre_norm_div_1_(injectionVector[4]),
.p_desc958_p_O_DFFX1pre_norm_div_1_(injectionVector[5]),
.p_desc959_p_O_DFFX1pre_norm_div_1_(injectionVector[6]),
.p_desc960_p_O_DFFX1pre_norm_div_1_(injectionVector[7]),
.p_desc961_p_O_DFFX1pre_norm_div_1_(injectionVector[8]),
.p_desc962_p_O_DFFX1pre_norm_div_1_(injectionVector[9]),
.p_desc963_p_O_DFFX1pre_norm_div_1_(injectionVector[10]),
.p_desc964_p_O_DFFX1pre_norm_div_1_(injectionVector[11]),
.p_desc965_p_O_DFFX1pre_norm_div_1_(injectionVector[12]),
.p_desc966_p_O_DFFX1pre_norm_div_1_(injectionVector[13]),
.p_desc967_p_O_DFFX1pre_norm_div_1_(injectionVector[14]),
.p_desc968_p_O_DFFX1pre_norm_div_1_(injectionVector[15]),
.p_desc969_p_O_DFFX1pre_norm_div_1_(injectionVector[16]),
.p_desc970_p_O_DFFX1pre_norm_div_1_(injectionVector[17]),
.p_desc971_p_O_DFFX1pre_norm_div_1_(injectionVector[18]),
.p_desc972_p_O_DFFX1pre_norm_div_1_(injectionVector[19]),
.p_desc973_p_O_DFFX1pre_norm_div_1_(injectionVector[20]),
.p_desc974_p_O_DFFX1pre_norm_div_1_(injectionVector[21]),
.p_desc975_p_O_DFFX1pre_norm_div_1_(injectionVector[22]),
.p_desc976_p_O_DFFX1pre_norm_div_1_(injectionVector[23]),
.p_desc977_p_O_DFFX1pre_norm_div_1_(injectionVector[24]),
.p_desc978_p_O_DFFX1pre_norm_div_1_(injectionVector[25]),
.p_desc979_p_O_DFFX1pre_norm_div_1_(injectionVector[26]),
.p_desc980_p_O_DFFX1pre_norm_div_1_(injectionVector[27]),
.p_desc981_p_O_DFFX1pre_norm_div_1_(injectionVector[28]),
.p_desc982_p_O_DFFX1pre_norm_div_1_(injectionVector[29]),
.p_desc983_p_O_DFFX1pre_norm_div_1_(injectionVector[30]),
.p_desc984_p_O_DFFX1pre_norm_div_1_(injectionVector[31]),
.p_desc985_p_O_DFFX1pre_norm_div_1_(injectionVector[32]),
.p_desc986_p_O_DFFX1pre_norm_div_1_(injectionVector[33]),
.p_desc987_p_O_DFFX1pre_norm_div_1_(injectionVector[34]),
.p_desc988_p_O_DFFX1pre_norm_div_1_(injectionVector[35]),
.p_desc989_p_O_DFFX1serial_div_1_(injectionVector[36]),
.p_desc990_p_O_DFFX1serial_div_1_(injectionVector[37]),
.p_desc991_p_O_DFFX1serial_div_1_(injectionVector[38]),
.p_desc992_p_O_DFFX1serial_div_1_(injectionVector[39]),
.p_desc993_p_O_DFFX1serial_div_1_(injectionVector[40]),
.p_desc994_p_O_DFFX1serial_div_1_(injectionVector[41]),
.p_desc995_p_O_DFFX1serial_div_1_(injectionVector[42]),
.p_desc996_p_O_DFFX1serial_div_1_(injectionVector[43]),
.p_desc997_p_O_DFFX1serial_div_1_(injectionVector[44]),
.p_desc998_p_O_DFFX1serial_div_1_(injectionVector[45]),
.p_desc999_p_O_DFFX1serial_div_1_(injectionVector[46]),
.p_desc1000_p_O_DFFX1serial_div_1_(injectionVector[47]),
.p_desc1001_p_O_DFFX1serial_div_1_(injectionVector[48]),
.p_desc1002_p_O_DFFX1serial_div_1_(injectionVector[49]),
.p_desc1003_p_O_DFFX1serial_div_1_(injectionVector[50]),
.p_desc1004_p_O_DFFX1serial_div_1_(injectionVector[51]),
.p_desc1005_p_O_DFFX1serial_div_1_(injectionVector[52]),
.p_desc1006_p_O_DFFX1serial_div_1_(injectionVector[53]),
.p_desc1007_p_O_DFFX1serial_div_1_(injectionVector[54]),
.p_desc1008_p_O_DFFX1serial_div_1_(injectionVector[55]),
.p_desc1009_p_O_DFFX1serial_div_1_(injectionVector[56]),
.p_desc1010_p_O_DFFX1serial_div_1_(injectionVector[57]),
.p_desc1011_p_O_DFFX1serial_div_1_(injectionVector[58]),
.p_desc1012_p_O_DFFX1serial_div_1_(injectionVector[59]),
.p_desc1013_p_O_DFFX1serial_div_1_(injectionVector[60]),
.p_desc1014_p_O_DFFX1serial_div_1_(injectionVector[61]),
.p_desc1015_p_O_DFFX1serial_div_1_(injectionVector[62]),
.p_desc1016_p_O_DFFX1serial_div_1_(injectionVector[63]),
.p_desc1017_p_O_DFFX1serial_div_1_(injectionVector[64]),
.p_desc1018_p_O_DFFX1serial_div_1_(injectionVector[65]),
.p_desc1019_p_O_DFFX1serial_div_1_(injectionVector[66]),
.p_desc1020_p_O_DFFX1serial_div_1_(injectionVector[67]),
.p_desc1021_p_O_DFFX1serial_div_1_(injectionVector[68]),
.p_desc1022_p_O_DFFX1serial_div_1_(injectionVector[69]),
.p_desc1023_p_O_DFFX1serial_div_1_(injectionVector[70]),
.p_desc1024_p_O_DFFX1serial_div_1_(injectionVector[71]),
.p_desc1025_p_O_DFFX1serial_div_1_(injectionVector[72]),
.p_desc1026_p_O_DFFX1serial_div_1_(injectionVector[73]),
.p_desc1027_p_O_DFFX1serial_div_1_(injectionVector[74]),
.p_desc1028_p_O_DFFX1serial_div_1_(injectionVector[75]),
.p_desc1029_p_O_DFFX1serial_div_1_(injectionVector[76]),
.p_desc1030_p_O_DFFX1serial_div_1_(injectionVector[77]),
.p_desc1031_p_O_DFFX1serial_div_1_(injectionVector[78]),
.p_desc1032_p_O_DFFX1serial_div_1_(injectionVector[79]),
.p_desc1033_p_O_DFFX1serial_div_1_(injectionVector[80]),
.p_desc1034_p_O_DFFX1serial_div_1_(injectionVector[81]),
.p_desc1035_p_O_DFFX1serial_div_1_(injectionVector[82]),
.p_desc1036_p_O_DFFX1serial_div_1_(injectionVector[83]),
.p_desc1037_p_O_DFFX1serial_div_1_(injectionVector[84]),
.p_desc1038_p_O_DFFX1serial_div_1_(injectionVector[85]),
.p_desc1039_p_O_DFFX1serial_div_1_(injectionVector[86]),
.p_desc1040_p_O_DFFX1serial_div_1_(injectionVector[87]),
.p_desc1041_p_O_DFFX1serial_div_1_(injectionVector[88]),
.p_desc1042_p_O_DFFX1serial_div_1_(injectionVector[89]),
.p_desc1043_p_O_DFFX1serial_div_1_(injectionVector[90]),
.p_desc1044_p_O_DFFX1serial_div_1_(injectionVector[91]),
.p_desc1045_p_O_DFFX1serial_div_1_(injectionVector[92]),
.p_desc1046_p_O_DFFX1serial_div_1_(injectionVector[93]),
.p_desc1047_p_O_DFFX1serial_div_1_(injectionVector[94]),
.p_desc1048_p_O_DFFX1serial_div_1_(injectionVector[95]),
.p_desc1049_p_O_DFFX1serial_div_1_(injectionVector[96]),
.p_desc1050_p_O_DFFX1serial_div_1_(injectionVector[97]),
.p_desc1051_p_O_DFFX1serial_div_1_(injectionVector[98]),
.p_desc1052_p_O_DFFX1serial_div_1_(injectionVector[99]),
.p_desc1053_p_O_DFFX1serial_div_1_(injectionVector[100]),
.p_desc1054_p_O_DFFX1serial_div_1_(injectionVector[101]),
.p_desc1055_p_O_DFFX1serial_div_1_(injectionVector[102]),
.p_desc1056_p_O_DFFX1serial_div_1_(injectionVector[103]),
.p_desc1057_p_O_DFFX1serial_div_1_(injectionVector[104]),
.p_desc1058_p_O_DFFX1serial_div_1_(injectionVector[105]),
.p_desc1059_p_O_DFFX1serial_div_1_(injectionVector[106]),
.p_desc1060_p_O_DFFX1serial_div_1_(injectionVector[107]),
.p_desc1061_p_O_DFFX1serial_div_1_(injectionVector[108]),
.p_desc1062_p_O_DFFX1serial_div_1_(injectionVector[109]),
.p_desc1063_p_O_DFFX1serial_div_1_(injectionVector[110]),
.p_desc1064_p_O_DFFX1serial_div_1_(injectionVector[111]),
.p_desc1065_p_O_DFFX1serial_div_1_(injectionVector[112]),
.p_s_start_i_reg_p_O_DFFX1serial_div_1_(injectionVector[113]),
.p_desc1066_p_O_DFFX1serial_div_1_(injectionVector[114]),
.p_s_state_reg_p_O_DFFX1serial_div_1_(injectionVector[115]),
.p_s_ready_o_reg_p_O_DFFX1serial_div_1_(injectionVector[116]),
.p_desc1067_p_O_DFFX1serial_div_1_(injectionVector[117]),
.p_desc1068_p_O_DFFX1serial_div_1_(injectionVector[118]),
.p_desc1069_p_O_DFFX1serial_div_1_(injectionVector[119]),
.p_desc1070_p_O_DFFX1serial_div_1_(injectionVector[120]),
.p_desc1071_p_O_DFFX1serial_div_1_(injectionVector[121]),
.p_desc1072_p_O_DFFX1serial_div_1_(injectionVector[122]),
.p_desc1073_p_O_DFFX1serial_div_1_(injectionVector[123]),
.p_desc1074_p_O_DFFX1serial_div_1_(injectionVector[124]),
.p_desc1075_p_O_DFFX1serial_div_1_(injectionVector[125]),
.p_desc1076_p_O_DFFX1serial_div_1_(injectionVector[126]),
.p_desc1077_p_O_DFFX1serial_div_1_(injectionVector[127]),
.p_desc1078_p_O_DFFX1serial_div_1_(injectionVector[128]),
.p_desc1079_p_O_DFFX1serial_div_1_(injectionVector[129]),
.p_desc1080_p_O_DFFX1serial_div_1_(injectionVector[130]),
.p_desc1081_p_O_DFFX1serial_div_1_(injectionVector[131]),
.p_desc1082_p_O_DFFX1serial_div_1_(injectionVector[132]),
.p_desc1083_p_O_DFFX1serial_div_1_(injectionVector[133]),
.p_desc1084_p_O_DFFX1serial_div_1_(injectionVector[134]),
.p_desc1085_p_O_DFFX1serial_div_1_(injectionVector[135]),
.p_desc1086_p_O_DFFX1serial_div_1_(injectionVector[136]),
.p_desc1087_p_O_DFFX1serial_div_1_(injectionVector[137]),
.p_desc1088_p_O_DFFX1serial_div_1_(injectionVector[138]),
.p_desc1089_p_O_DFFX1serial_div_1_(injectionVector[139]),
.p_desc1090_p_O_DFFX1serial_div_1_(injectionVector[140]),
.p_desc1091_p_O_DFFX1serial_div_1_(injectionVector[141]),
.p_desc1092_p_O_DFFX1serial_div_1_(injectionVector[142]),
.p_desc1093_p_O_DFFX1serial_div_1_(injectionVector[143]),
.p_desc1094_p_O_DFFX1serial_div_1_(injectionVector[144]),
.p_desc1095_p_O_DFFX1serial_div_1_(injectionVector[145]),
.p_desc1096_p_O_DFFX1serial_div_1_(injectionVector[146]),
.p_desc1097_p_O_DFFX1serial_div_1_(injectionVector[147]),
.p_desc1098_p_O_DFFX1serial_div_1_(injectionVector[148]),
.p_desc1099_p_O_DFFX1serial_div_1_(injectionVector[149]),
.p_desc1100_p_O_DFFX1serial_div_1_(injectionVector[150]),
.p_desc1101_p_O_DFFX1serial_div_1_(injectionVector[151]),
.p_desc1102_p_O_DFFX1serial_div_1_(injectionVector[152]),
.p_desc1103_p_O_DFFX1serial_div_1_(injectionVector[153]),
.p_desc1104_p_O_DFFX1serial_div_1_(injectionVector[154]),
.p_desc1105_p_O_DFFX1serial_div_1_(injectionVector[155]),
.p_desc1106_p_O_DFFX1serial_div_1_(injectionVector[156]),
.p_desc1107_p_O_DFFX1serial_div_1_(injectionVector[157]),
.p_desc1108_p_O_DFFX1serial_div_1_(injectionVector[158]),
.p_desc1109_p_O_DFFX1serial_div_1_(injectionVector[159]),
.p_desc1110_p_O_DFFX1serial_div_1_(injectionVector[160]),
.p_desc1111_p_O_DFFX1serial_div_1_(injectionVector[161]),
.p_desc1112_p_O_DFFX1serial_div_1_(injectionVector[162]),
.p_desc1113_p_O_DFFX1serial_div_1_(injectionVector[163]),
.p_desc1114_p_O_DFFX1serial_div_1_(injectionVector[164]),
.p_desc1115_p_O_DFFX1serial_div_1_(injectionVector[165]),
.p_desc1116_p_O_DFFX1serial_div_1_(injectionVector[166]),
.p_desc1117_p_O_DFFX1serial_div_1_(injectionVector[167]),
.p_desc1118_p_O_DFFX1serial_div_1_(injectionVector[168]),
.p_desc1119_p_O_DFFX1serial_div_1_(injectionVector[169]),
.p_desc1120_p_O_DFFX1serial_div_1_(injectionVector[170]),
.p_desc1121_p_O_DFFX1serial_div_1_(injectionVector[171]),
.p_desc1122_p_O_DFFX1serial_div_1_(injectionVector[172]),
.p_desc1123_p_O_DFFX1serial_div_1_(injectionVector[173]),
.p_desc1124_p_O_DFFX1serial_div_1_(injectionVector[174]),
.p_desc1125_p_O_DFFX1serial_div_1_(injectionVector[175]),
.p_desc1126_p_O_DFFX1serial_div_1_(injectionVector[176]),
.p_desc1127_p_O_DFFX1serial_div_1_(injectionVector[177]),
.p_desc1128_p_O_DFFX1serial_div_1_(injectionVector[178]),
.p_desc1129_p_O_DFFX1serial_div_1_(injectionVector[179]),
.p_desc1130_p_O_DFFX1serial_div_1_(injectionVector[180]),
.p_desc1131_p_O_DFFX1serial_div_1_(injectionVector[181]),
.p_desc1132_p_O_DFFX1serial_div_1_(injectionVector[182]),
.p_desc1133_p_O_DFFX1serial_div_1_(injectionVector[183]),
.p_desc1134_p_O_DFFX1serial_div_1_(injectionVector[184]),
.p_desc1135_p_O_DFFX1serial_div_1_(injectionVector[185]),
.p_desc1136_p_O_DFFX1serial_div_1_(injectionVector[186]),
.p_desc1137_p_O_DFFX1serial_div_1_(injectionVector[187]),
.p_desc1138_p_O_DFFX1serial_div_1_(injectionVector[188]),
.p_desc1139_p_O_DFFX1serial_div_1_(injectionVector[189]),
.p_desc1140_p_O_DFFX1serial_div_1_(injectionVector[190]),
.p_desc1141_p_O_DFFX1serial_div_1_(injectionVector[191]),
.p_desc1142_p_O_DFFX1serial_div_1_(injectionVector[192]),
.p_desc1143_p_O_DFFX1serial_div_1_(injectionVector[193]),
.p_desc1144_p_O_DFFX1serial_div_1_(injectionVector[194]),
.p_desc1145_p_O_DFFX1serial_div_1_(injectionVector[195]),
.p_desc1146_p_O_DFFX1serial_div_1_(injectionVector[196]),
.p_desc1147_p_O_DFFX1serial_div_1_(injectionVector[197]),
.p_desc1148_p_O_DFFX1serial_div_1_(injectionVector[198]),
.p_desc1149_p_O_DFFX1serial_div_1_(injectionVector[199]),
.p_desc1150_p_O_DFFX1serial_div_1_(injectionVector[200]),
.p_desc1151_p_O_DFFX1post_norm_div_1_(injectionVector[201]),
.p_desc1152_p_O_DFFX1post_norm_div_1_(injectionVector[202]),
.p_desc1153_p_O_DFFX1post_norm_div_1_(injectionVector[203]),
.p_desc1154_p_O_DFFX1post_norm_div_1_(injectionVector[204]),
.p_desc1155_p_O_DFFX1post_norm_div_1_(injectionVector[205]),
.p_desc1156_p_O_DFFX1post_norm_div_1_(injectionVector[206]),
.p_desc1157_p_O_DFFX1post_norm_div_1_(injectionVector[207]),
.p_desc1158_p_O_DFFX1post_norm_div_1_(injectionVector[208]),
.p_desc1159_p_O_DFFX1post_norm_div_1_(injectionVector[209]),
.p_desc1160_p_O_DFFX1post_norm_div_1_(injectionVector[210]),
.p_desc1161_p_O_DFFX1post_norm_div_1_(injectionVector[211]),
.p_desc1162_p_O_DFFX1post_norm_div_1_(injectionVector[212]),
.p_desc1163_p_O_DFFX1post_norm_div_1_(injectionVector[213]),
.p_desc1164_p_O_DFFX1post_norm_div_1_(injectionVector[214]),
.p_desc1165_p_O_DFFX1post_norm_div_1_(injectionVector[215]),
.p_desc1166_p_O_DFFX1post_norm_div_1_(injectionVector[216]),
.p_desc1167_p_O_DFFX1post_norm_div_1_(injectionVector[217]),
.p_desc1168_p_O_DFFX1post_norm_div_1_(injectionVector[218]),
.p_desc1169_p_O_DFFX1post_norm_div_1_(injectionVector[219]),
.p_desc1170_p_O_DFFX1post_norm_div_1_(injectionVector[220]),
.p_desc1171_p_O_DFFX1post_norm_div_1_(injectionVector[221]),
.p_desc1172_p_O_DFFX1post_norm_div_1_(injectionVector[222]),
.p_desc1173_p_O_DFFX1post_norm_div_1_(injectionVector[223]),
.p_desc1174_p_O_DFFX1post_norm_div_1_(injectionVector[224]),
.p_desc1175_p_O_DFFX1post_norm_div_1_(injectionVector[225]),
.p_desc1176_p_O_DFFX1post_norm_div_1_(injectionVector[226]),
.p_desc1177_p_O_DFFX1post_norm_div_1_(injectionVector[227]),
.p_desc1178_p_O_DFFX1post_norm_div_1_(injectionVector[228]),
.p_desc1179_p_O_DFFX1post_norm_div_1_(injectionVector[229]),
.p_desc1180_p_O_DFFX1post_norm_div_1_(injectionVector[230]),
.p_desc1181_p_O_DFFX1post_norm_div_1_(injectionVector[231]),
.p_desc1182_p_O_DFFX1post_norm_div_1_(injectionVector[232]),
.p_desc1183_p_O_DFFX1post_norm_div_1_(injectionVector[233]),
.p_desc1184_p_O_DFFX1post_norm_div_1_(injectionVector[234]),
.p_desc1185_p_O_DFFX1post_norm_div_1_(injectionVector[235]),
.p_desc1186_p_O_DFFX1post_norm_div_1_(injectionVector[236]),
.p_desc1187_p_O_DFFX1post_norm_div_1_(injectionVector[237]),
.p_desc1188_p_O_DFFX1post_norm_div_1_(injectionVector[238]),
.p_desc1189_p_O_DFFX1post_norm_div_1_(injectionVector[239]),
.p_desc1190_p_O_DFFX1post_norm_div_1_(injectionVector[240]),
.p_desc1191_p_O_DFFX1post_norm_div_1_(injectionVector[241]),
.p_desc1192_p_O_DFFX1post_norm_div_1_(injectionVector[242]),
.p_desc1193_p_O_DFFX1post_norm_div_1_(injectionVector[243]),
.p_desc1194_p_O_DFFX1post_norm_div_1_(injectionVector[244]),
.p_desc1195_p_O_DFFX1post_norm_div_1_(injectionVector[245]),
.p_desc1196_p_O_DFFX1post_norm_div_1_(injectionVector[246]),
.p_desc1197_p_O_DFFX1post_norm_div_1_(injectionVector[247]),
.p_desc1198_p_O_DFFX1post_norm_div_1_(injectionVector[248]),
.p_desc1199_p_O_DFFX1post_norm_div_1_(injectionVector[249]),
.p_desc1200_p_O_DFFX1post_norm_div_1_(injectionVector[250]),
.p_desc1201_p_O_DFFX1post_norm_div_1_(injectionVector[251]),
.p_desc1202_p_O_DFFX1post_norm_div_1_(injectionVector[252]),
.p_desc1203_p_O_DFFX1post_norm_div_1_(injectionVector[253]),
.p_desc1204_p_O_DFFX1post_norm_div_1_(injectionVector[254]),
.p_desc1205_p_O_DFFX1post_norm_div_1_(injectionVector[255]),
.p_desc1206_p_O_DFFX1post_norm_div_1_(injectionVector[256]),
.p_desc1207_p_O_DFFX1post_norm_div_1_(injectionVector[257]),
.p_desc1208_p_O_DFFX1post_norm_div_1_(injectionVector[258]),
.p_desc1209_p_O_DFFX1post_norm_div_1_(injectionVector[259]),
.p_desc1210_p_O_DFFX1post_norm_div_1_(injectionVector[260]),
.p_desc1211_p_O_DFFX1post_norm_div_1_(injectionVector[261]),
.p_desc1212_p_O_DFFX1post_norm_div_1_(injectionVector[262]),
.p_desc1213_p_O_DFFX1post_norm_div_1_(injectionVector[263]),
.p_desc1214_p_O_DFFX1post_norm_div_1_(injectionVector[264]),
.p_desc1215_p_O_DFFX1post_norm_div_1_(injectionVector[265]),
.p_desc1216_p_O_DFFX1post_norm_div_1_(injectionVector[266]),
.p_desc1217_p_O_DFFX1post_norm_div_1_(injectionVector[267]),
.p_desc1218_p_O_DFFX1post_norm_div_1_(injectionVector[268]),
.p_desc1219_p_O_DFFX1post_norm_div_1_(injectionVector[269]),
.p_desc1220_p_O_DFFX1post_norm_div_1_(injectionVector[270]),
.p_desc1221_p_O_DFFX1post_norm_div_1_(injectionVector[271]),
.p_desc1222_p_O_DFFX1post_norm_div_1_(injectionVector[272]),
.p_desc1223_p_O_DFFX1post_norm_div_1_(injectionVector[273]),
.p_desc1224_p_O_DFFX1post_norm_div_1_(injectionVector[274]),
.p_desc1225_p_O_DFFX1post_norm_div_1_(injectionVector[275]),
.p_desc1226_p_O_DFFX1post_norm_div_1_(injectionVector[276]),
.p_desc1227_p_O_DFFX1post_norm_div_1_(injectionVector[277]),
.p_desc1228_p_O_DFFX1post_norm_div_1_(injectionVector[278]),
.p_desc1229_p_O_DFFX1post_norm_div_1_(injectionVector[279]),
.p_desc1230_p_O_DFFX1post_norm_div_1_(injectionVector[280]),
.p_desc1231_p_O_DFFX1post_norm_div_1_(injectionVector[281]),
.p_desc1232_p_O_DFFX1post_norm_div_1_(injectionVector[282]),
.p_desc1233_p_O_DFFX1post_norm_div_1_(injectionVector[283]),
.p_desc1234_p_O_DFFX1post_norm_div_1_(injectionVector[284]),
.p_desc1235_p_O_DFFX1post_norm_div_1_(injectionVector[285]),
.p_desc1236_p_O_DFFX1post_norm_div_1_(injectionVector[286]),
.p_desc1237_p_O_DFFX1post_norm_div_1_(injectionVector[287]),
.p_desc1238_p_O_DFFX1post_norm_div_1_(injectionVector[288]),
.p_desc1239_p_O_DFFX1post_norm_div_1_(injectionVector[289]),
.p_desc1240_p_O_DFFX1post_norm_div_1_(injectionVector[290]),
.p_desc1241_p_O_DFFX1post_norm_div_1_(injectionVector[291]),
.p_desc1242_p_O_DFFX1post_norm_div_1_(injectionVector[292]),
.p_desc1243_p_O_DFFX1post_norm_div_1_(injectionVector[293]),
.p_desc1244_p_O_DFFX1post_norm_div_1_(injectionVector[294]),
.p_desc1245_p_O_DFFX1post_norm_div_1_(injectionVector[295]),
.p_desc1246_p_O_DFFX1post_norm_div_1_(injectionVector[296]),
.p_desc1247_p_O_DFFX1post_norm_div_1_(injectionVector[297]),
.p_desc1248_p_O_DFFX1post_norm_div_1_(injectionVector[298]),
.p_desc1249_p_O_DFFX1post_norm_div_1_(injectionVector[299]),
.p_desc1250_p_O_DFFX1post_norm_div_1_(injectionVector[300]),
.p_desc1251_p_O_DFFX1post_norm_div_1_(injectionVector[301]),
.p_desc1252_p_O_DFFX1post_norm_div_1_(injectionVector[302]),
.p_desc1253_p_O_DFFX1post_norm_div_1_(injectionVector[303]),
.p_desc1254_p_O_DFFX1post_norm_div_1_(injectionVector[304]),
.p_desc1255_p_O_DFFX1post_norm_div_1_(injectionVector[305]),
.p_desc1256_p_O_DFFX1post_norm_div_1_(injectionVector[306]),
.p_desc1257_p_O_DFFX1post_norm_div_1_(injectionVector[307]),
.p_desc1258_p_O_DFFX1post_norm_div_1_(injectionVector[308]),
.p_desc1259_p_O_DFFX1post_norm_div_1_(injectionVector[309]),
.p_desc1260_p_O_DFFX1post_norm_div_1_(injectionVector[310]),
.p_desc1261_p_O_DFFX1post_norm_div_1_(injectionVector[311]),
.p_desc1262_p_O_DFFX1post_norm_div_1_(injectionVector[312]),
.p_desc1263_p_O_DFFX1post_norm_div_1_(injectionVector[313]),
.p_desc1264_p_O_DFFX1post_norm_div_1_(injectionVector[314]),
.p_desc1265_p_O_DFFX1post_norm_div_1_(injectionVector[315]),
.p_desc1266_p_O_DFFX1post_norm_div_1_(injectionVector[316]),
.p_desc1267_p_O_DFFX1post_norm_div_1_(injectionVector[317]),
.p_desc1268_p_O_DFFX1post_norm_div_1_(injectionVector[318]),
.p_desc1269_p_O_DFFX1post_norm_div_1_(injectionVector[319]),
.p_desc1270_p_O_DFFX1post_norm_div_1_(injectionVector[320]),
.p_desc1271_p_O_DFFX1post_norm_div_1_(injectionVector[321]),
.p_desc1272_p_O_DFFX1post_norm_div_1_(injectionVector[322]),
.p_desc1273_p_O_DFFX1post_norm_div_1_(injectionVector[323]),
.p_desc1274_p_O_DFFX1post_norm_div_1_(injectionVector[324]),
.p_desc1275_p_O_DFFX1post_norm_div_1_(injectionVector[325]),
.p_desc1276_p_O_DFFX1post_norm_div_1_(injectionVector[326]),
.p_desc1277_p_O_DFFX1post_norm_div_1_(injectionVector[327]),
.p_desc1278_p_O_DFFX1post_norm_div_1_(injectionVector[328]),
.p_desc1279_p_O_DFFX1post_norm_div_1_(injectionVector[329]),
.p_desc1280_p_O_DFFX1post_norm_div_1_(injectionVector[330]),
.p_desc1281_p_O_DFFX1post_norm_div_1_(injectionVector[331]),
.p_desc1282_p_O_DFFX1post_norm_div_1_(injectionVector[332]),
.p_desc1283_p_O_DFFX1post_norm_div_1_(injectionVector[333]),
.p_desc1284_p_O_DFFX1post_norm_div_1_(injectionVector[334]),
.p_desc1285_p_O_DFFX1post_norm_div_1_(injectionVector[335]),
.p_desc1286_p_O_DFFX1post_norm_div_1_(injectionVector[336]),
.p_desc1287_p_O_DFFX1post_norm_div_1_(injectionVector[337]),
.p_desc1288_p_O_DFFX1post_norm_div_1_(injectionVector[338]),
.p_desc1289_p_O_DFFX1post_norm_div_1_(injectionVector[339]),
.p_desc1290_p_O_DFFX1post_norm_div_1_(injectionVector[340]),
.p_desc1291_p_O_DFFX1post_norm_div_1_(injectionVector[341]),
.p_desc1292_p_O_DFFX1post_norm_div_1_(injectionVector[342]),
.p_s_sign_i_reg_p_O_DFFX1post_norm_div_1_(injectionVector[343]),
.p_desc1293_p_O_DFFX1post_norm_div_1_(injectionVector[344]),
.p_desc1294_p_O_DFFX1post_norm_div_1_(injectionVector[345]),
.p_desc1295_p_O_DFFX1post_norm_div_1_(injectionVector[346]),
.p_desc1299_p_O_DFFX1post_norm_div_1_(injectionVector[347]),
.p_desc1300_p_O_DFFX1post_norm_div_1_(injectionVector[348]),
.p_desc1304_p_O_DFFX1post_norm_div_1_(injectionVector[349]),
.p_desc1305_p_O_DFFX1post_norm_div_1_(injectionVector[350]),
.p_desc1306_p_O_DFFX1post_norm_div_1_(injectionVector[351]),
.p_desc1307_p_O_DFFX1post_norm_div_1_(injectionVector[352]),
.p_desc1308_p_O_DFFX1post_norm_div_1_(injectionVector[353]),
.p_desc1309_p_O_DFFX1post_norm_div_1_(injectionVector[354]),
.p_desc1310_p_O_DFFX1post_norm_div_1_(injectionVector[355]),
.p_desc1311_p_O_DFFX1post_norm_div_1_(injectionVector[356]),
.p_desc1312_p_O_DFFX1post_norm_div_1_(injectionVector[357]),
.p_desc1313_p_O_DFFX1post_norm_div_1_(injectionVector[358]),
.p_desc1314_p_O_DFFX1post_norm_div_1_(injectionVector[359]),
.p_desc1315_p_O_DFFX1post_norm_div_1_(injectionVector[360]),
.p_desc1316_p_O_DFFX1post_norm_div_1_(injectionVector[361]),
.p_desc1317_p_O_DFFX1post_norm_div_1_(injectionVector[362]),
.p_desc1318_p_O_DFFX1post_norm_div_1_(injectionVector[363]),
.p_desc1319_p_O_DFFX1post_norm_div_1_(injectionVector[364]),
.p_desc1320_p_O_DFFX1post_norm_div_1_(injectionVector[365]),
.p_desc1321_p_O_DFFX1post_norm_div_1_(injectionVector[366]),
.p_desc1322_p_O_DFFX1post_norm_div_1_(injectionVector[367]),
.p_desc1323_p_O_DFFX1post_norm_div_1_(injectionVector[368]),
.p_desc1324_p_O_DFFX1post_norm_div_1_(injectionVector[369]),
.p_desc1325_p_O_DFFX1post_norm_div_1_(injectionVector[370]),
.p_desc1326_p_O_DFFX1post_norm_div_1_(injectionVector[371]),
.p_desc1327_p_O_DFFX1post_norm_div_1_(injectionVector[372]),
.p_desc1328_p_O_DFFX1post_norm_div_1_(injectionVector[373]),
.p_desc1329_p_O_DFFX1post_norm_div_1_(injectionVector[374]),
.p_desc1330_p_O_DFFX1post_norm_div_1_(injectionVector[375]),
.p_desc1331_p_O_DFFX1post_norm_div_1_(injectionVector[376]),
.p_desc1332_p_O_DFFX1post_norm_div_1_(injectionVector[377]),
.p_desc1333_p_O_DFFX1post_norm_div_1_(injectionVector[378]),
.p_desc1334_p_O_DFFX1post_norm_div_1_(injectionVector[379]),
.p_desc1335_p_O_DFFX1post_norm_div_1_(injectionVector[380]),
.p_desc1336_p_O_DFFX1post_norm_div_1_(injectionVector[381]),
.p_desc1337_p_O_DFFX1post_norm_div_1_(injectionVector[382]),
.p_desc1338_p_O_DFFX1post_norm_div_1_(injectionVector[383]),
.p_desc1339_p_O_DFFX1post_norm_div_1_(injectionVector[384]),
.p_desc1340_p_O_DFFX1post_norm_div_1_(injectionVector[385]),
.p_desc1341_p_O_DFFX1post_norm_div_1_(injectionVector[386]),
.p_desc1342_p_O_DFFX1post_norm_div_1_(injectionVector[387]),
.p_desc1343_p_O_DFFX1post_norm_div_1_(injectionVector[388]),
.p_desc1344_p_O_DFFX1post_norm_div_1_(injectionVector[389]),
.p_desc1345_p_O_DFFX1post_norm_div_1_(injectionVector[390]),
.p_desc1346_p_O_DFFX1post_norm_div_1_(injectionVector[391]),
.p_desc1347_p_O_DFFX1post_norm_div_1_(injectionVector[392]),
.p_desc1348_p_O_DFFX1post_norm_div_1_(injectionVector[393]),
.p_desc1349_p_O_DFFX1post_norm_div_1_(injectionVector[394]),
.p_desc1350_p_O_DFFX1post_norm_div_1_(injectionVector[395]),
.p_desc1351_p_O_DFFX1post_norm_div_1_(injectionVector[396]),
.p_desc1352_p_O_DFFX1post_norm_div_1_(injectionVector[397]),
.p_desc1353_p_O_DFFX1post_norm_div_1_(injectionVector[398]),
.p_desc1354_p_O_DFFX1post_norm_div_1_(injectionVector[399]),
.p_desc1355_p_O_DFFX1post_norm_div_1_(injectionVector[400]),
.p_desc1356_p_O_DFFX1post_norm_div_1_(injectionVector[401]),
.p_desc1357_p_O_DFFX1post_norm_div_1_(injectionVector[402]),
.p_desc1358_p_O_DFFX1post_norm_div_1_(injectionVector[403]),
.p_desc1359_p_O_DFFX1post_norm_div_1_(injectionVector[404]),
.p_desc1360_p_O_DFFX1post_norm_div_1_(injectionVector[405]),
.p_desc1361_p_O_DFFX1post_norm_div_1_(injectionVector[406]),
.p_desc1362_p_O_DFFX1post_norm_div_1_(injectionVector[407]),
.p_desc1363_p_O_DFFX1post_norm_div_1_(injectionVector[408]),
.p_desc1364_p_O_DFFX1post_norm_div_1_(injectionVector[409]),
.p_desc1365_p_O_DFFX1post_norm_div_1_(injectionVector[410]),
.p_desc1366_p_O_DFFX1post_norm_div_1_(injectionVector[411]),
.p_desc1367_p_O_DFFX1post_norm_div_1_(injectionVector[412]),
.p_desc1368_p_O_DFFX1post_norm_div_1_(injectionVector[413]),
.p_desc1369_p_O_DFFX1post_norm_div_1_(injectionVector[414]),
.p_desc1370_p_O_DFFX1post_norm_div_1_(injectionVector[415]),
.p_ine_o_reg_p_O_DFFX1post_norm_div_1_(injectionVector[416]),
.p_desc1371_p_O_DFFX1post_norm_div_1_(injectionVector[417]),
.p_desc1379_p_O_DFFX1post_norm_div_1_(injectionVector[418]),
.p_desc1380_p_O_DFFX1post_norm_div_1_(injectionVector[419]),
.p_desc1381_p_O_DFFX1post_norm_div_1_(injectionVector[420]),
.p_desc1382_p_O_DFFX1post_norm_div_1_(injectionVector[421]),
.p_desc1383_p_O_DFFX1post_norm_div_1_(injectionVector[422]),
.p_desc1384_p_O_DFFX1post_norm_div_1_(injectionVector[423]),
.p_desc1385_p_O_DFFX1post_norm_div_1_(injectionVector[424]),
.p_desc1386_p_O_DFFX1post_norm_div_1_(injectionVector[425]),
.p_desc1387_p_O_DFFX1post_norm_div_1_(injectionVector[426]),
.p_desc1388_p_O_DFFX1post_norm_div_1_(injectionVector[427]),
.p_desc1389_p_O_DFFX1post_norm_div_1_(injectionVector[428]),
.p_desc1390_p_O_DFFX1post_norm_div_1_(injectionVector[429]),
.p_desc1391_p_O_DFFX1post_norm_div_1_(injectionVector[430]),
.p_desc1392_p_O_DFFX1post_norm_div_1_(injectionVector[431]),
.p_desc1393_p_O_DFFX1post_norm_div_1_(injectionVector[432]),
.p_desc1394_p_O_DFFX1post_norm_div_1_(injectionVector[433]),
.p_desc1395_p_O_DFFX1post_norm_div_1_(injectionVector[434]),
.p_desc1396_p_O_DFFX1post_norm_div_1_(injectionVector[435]),
.p_desc1397_p_O_DFFX1post_norm_div_1_(injectionVector[436]),
.p_desc1398_p_O_DFFX1post_norm_div_1_(injectionVector[437]),
.p_desc1399_p_O_DFFX1post_norm_div_1_(injectionVector[438]),
.p_desc1400_p_O_DFFX1post_norm_div_1_(injectionVector[439]));
endmodule