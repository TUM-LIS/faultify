module add_subZ0_add_r_inj (mult_out_r,out_inner_prod_r,un2_pre_out_10,un2_pre_out_9,un2_pre_out_7,un2_pre_out_6,un2_pre_out_5,un2_pre_out_4,un2_pre_out_3,un2_pre_out_2,un2_pre_out_1,acc_clear,un2_pre_out_s_11,N_26_i,N_20_i);
input [11:0] mult_out_r ;
input [11:0] out_inner_prod_r ;
output un2_pre_out_10 ;
output un2_pre_out_9 ;
output un2_pre_out_7 ;
output un2_pre_out_6 ;
output un2_pre_out_5 ;
output un2_pre_out_4 ;
output un2_pre_out_3 ;
output un2_pre_out_2 ;
output un2_pre_out_1 ;
input acc_clear ;
output un2_pre_out_s_11 ;
output N_26_i ;
output N_20_i ;
wire un2_pre_out_10 ;
wire un2_pre_out_9 ;
wire un2_pre_out_7 ;
wire un2_pre_out_6 ;
wire un2_pre_out_5 ;
wire un2_pre_out_4 ;
wire un2_pre_out_3 ;
wire un2_pre_out_2 ;
wire un2_pre_out_1 ;
wire acc_clear ;
wire un2_pre_out_s_11 ;
wire N_26_i ;
wire N_20_i ;
wire [8:0] un2_pre_out ;
wire VCC ;
wire un2_pre_out_axb_1 ;
wire un2_pre_out_axb_2 ;
wire un2_pre_out_axb_3 ;
wire un2_pre_out_axb_4 ;
wire un2_pre_out_axb_5 ;
wire un2_pre_out_axb_6 ;
wire un2_pre_out_axb_7 ;
wire un2_pre_out_axb_8 ;
wire un2_pre_out_axb_9 ;
wire un2_pre_out_axb_10 ;
wire un2_pre_out_axb_11 ;
wire un2_pre_out_cry_10 ;
wire un2_pre_out_cry_9 ;
wire un2_pre_out_cry_8 ;
wire un2_pre_out_cry_7 ;
wire un2_pre_out_cry_6 ;
wire un2_pre_out_cry_5 ;
wire un2_pre_out_cry_4 ;
wire un2_pre_out_cry_3 ;
wire un2_pre_out_cry_2 ;
wire un2_pre_out_cry_1 ;
wire un2_pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 un2_pre_out_axb_0(.I0(mult_out_r[0:0]),.I1(out_inner_prod_r[0:0]),.O(un2_pre_out[0:0]));
defparam un2_pre_out_axb_0.INIT=4'h6;
  LUT2 un2_pre_out_axb_1_cZ(.I0(mult_out_r[1:1]),.I1(out_inner_prod_r[1:1]),.O(un2_pre_out_axb_1));
defparam un2_pre_out_axb_1_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_2_cZ(.I0(mult_out_r[2:2]),.I1(out_inner_prod_r[2:2]),.O(un2_pre_out_axb_2));
defparam un2_pre_out_axb_2_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_3_cZ(.I0(mult_out_r[3:3]),.I1(out_inner_prod_r[3:3]),.O(un2_pre_out_axb_3));
defparam un2_pre_out_axb_3_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_4_cZ(.I0(mult_out_r[4:4]),.I1(out_inner_prod_r[4:4]),.O(un2_pre_out_axb_4));
defparam un2_pre_out_axb_4_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_5_cZ(.I0(mult_out_r[5:5]),.I1(out_inner_prod_r[5:5]),.O(un2_pre_out_axb_5));
defparam un2_pre_out_axb_5_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_6_cZ(.I0(mult_out_r[6:6]),.I1(out_inner_prod_r[6:6]),.O(un2_pre_out_axb_6));
defparam un2_pre_out_axb_6_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_7_cZ(.I0(mult_out_r[7:7]),.I1(out_inner_prod_r[7:7]),.O(un2_pre_out_axb_7));
defparam un2_pre_out_axb_7_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_8_cZ(.I0(mult_out_r[8:8]),.I1(out_inner_prod_r[8:8]),.O(un2_pre_out_axb_8));
defparam un2_pre_out_axb_8_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_9_cZ(.I0(mult_out_r[9:9]),.I1(out_inner_prod_r[9:9]),.O(un2_pre_out_axb_9));
defparam un2_pre_out_axb_9_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_10_cZ(.I0(mult_out_r[10:10]),.I1(out_inner_prod_r[10:10]),.O(un2_pre_out_axb_10));
defparam un2_pre_out_axb_10_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_11_cZ(.I0(mult_out_r[11:11]),.I1(out_inner_prod_r[11:11]),.O(un2_pre_out_axb_11));
defparam un2_pre_out_axb_11_cZ.INIT=4'h6;
  XORCY un2_pre_out_s_11_c(.LI(un2_pre_out_axb_11),.CI(un2_pre_out_cry_10),.O(un2_pre_out_s_11));
  XORCY un2_pre_out_s_10(.LI(un2_pre_out_axb_10),.CI(un2_pre_out_cry_9),.O(un2_pre_out_10));
  MUXCY_L un2_pre_out_cry_10_cZ(.DI(mult_out_r[10:10]),.CI(un2_pre_out_cry_9),.S(un2_pre_out_axb_10),.LO(un2_pre_out_cry_10));
  XORCY un2_pre_out_s_9(.LI(un2_pre_out_axb_9),.CI(un2_pre_out_cry_8),.O(un2_pre_out_9));
  MUXCY_L un2_pre_out_cry_9_cZ(.DI(mult_out_r[9:9]),.CI(un2_pre_out_cry_8),.S(un2_pre_out_axb_9),.LO(un2_pre_out_cry_9));
  XORCY un2_pre_out_s_8(.LI(un2_pre_out_axb_8),.CI(un2_pre_out_cry_7),.O(un2_pre_out[8:8]));
  MUXCY_L un2_pre_out_cry_8_cZ(.DI(mult_out_r[8:8]),.CI(un2_pre_out_cry_7),.S(un2_pre_out_axb_8),.LO(un2_pre_out_cry_8));
  XORCY un2_pre_out_s_7(.LI(un2_pre_out_axb_7),.CI(un2_pre_out_cry_6),.O(un2_pre_out_7));
  MUXCY_L un2_pre_out_cry_7_cZ(.DI(mult_out_r[7:7]),.CI(un2_pre_out_cry_6),.S(un2_pre_out_axb_7),.LO(un2_pre_out_cry_7));
  XORCY un2_pre_out_s_6(.LI(un2_pre_out_axb_6),.CI(un2_pre_out_cry_5),.O(un2_pre_out_6));
  MUXCY_L un2_pre_out_cry_6_cZ(.DI(mult_out_r[6:6]),.CI(un2_pre_out_cry_5),.S(un2_pre_out_axb_6),.LO(un2_pre_out_cry_6));
  XORCY un2_pre_out_s_5(.LI(un2_pre_out_axb_5),.CI(un2_pre_out_cry_4),.O(un2_pre_out_5));
  MUXCY_L un2_pre_out_cry_5_cZ(.DI(mult_out_r[5:5]),.CI(un2_pre_out_cry_4),.S(un2_pre_out_axb_5),.LO(un2_pre_out_cry_5));
  XORCY un2_pre_out_s_4(.LI(un2_pre_out_axb_4),.CI(un2_pre_out_cry_3),.O(un2_pre_out_4));
  MUXCY_L un2_pre_out_cry_4_cZ(.DI(mult_out_r[4:4]),.CI(un2_pre_out_cry_3),.S(un2_pre_out_axb_4),.LO(un2_pre_out_cry_4));
  XORCY un2_pre_out_s_3(.LI(un2_pre_out_axb_3),.CI(un2_pre_out_cry_2),.O(un2_pre_out_3));
  MUXCY_L un2_pre_out_cry_3_cZ(.DI(mult_out_r[3:3]),.CI(un2_pre_out_cry_2),.S(un2_pre_out_axb_3),.LO(un2_pre_out_cry_3));
  XORCY un2_pre_out_s_2(.LI(un2_pre_out_axb_2),.CI(un2_pre_out_cry_1),.O(un2_pre_out_2));
  MUXCY_L un2_pre_out_cry_2_cZ(.DI(mult_out_r[2:2]),.CI(un2_pre_out_cry_1),.S(un2_pre_out_axb_2),.LO(un2_pre_out_cry_2));
  XORCY un2_pre_out_s_1(.LI(un2_pre_out_axb_1),.CI(un2_pre_out_cry_0),.O(un2_pre_out_1));
  MUXCY_L un2_pre_out_cry_1_cZ(.DI(mult_out_r[1:1]),.CI(un2_pre_out_cry_0),.S(un2_pre_out_axb_1),.LO(un2_pre_out_cry_1));
  MUXCY_L un2_pre_out_cry_0_cZ(.DI(mult_out_r[0:0]),.CI(GND),.S(un2_pre_out[0:0]),.LO(un2_pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 un2_pre_out_s_8_RNIQ3111_o6(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out_s_11),.O(N_26_i));
defparam un2_pre_out_s_8_RNIQ3111_o6.INIT=16'h3220;
  LUT5 un2_pre_out_s_8_RNIQ3111_o5(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[8:8]),.I4(un2_pre_out_s_11),.O(N_20_i));
defparam un2_pre_out_s_8_RNIQ3111_o5.INIT=32'h33011300;
endmodule
module add_subZ0_add_r_1_inj (mult_out_i,out_inner_prod_i,un2_pre_out_10,un2_pre_out_9,un2_pre_out_8,un2_pre_out_7,un2_pre_out_6,un2_pre_out_5,un2_pre_out_4,un2_pre_out_3,un2_pre_out_2,un2_pre_out_1,un2_pre_out_s_11_0);
input [11:0] mult_out_i ;
input [11:0] out_inner_prod_i ;
output un2_pre_out_10 ;
output un2_pre_out_9 ;
output un2_pre_out_8 ;
output un2_pre_out_7 ;
output un2_pre_out_6 ;
output un2_pre_out_5 ;
output un2_pre_out_4 ;
output un2_pre_out_3 ;
output un2_pre_out_2 ;
output un2_pre_out_1 ;
output un2_pre_out_s_11_0 ;
wire un2_pre_out_10 ;
wire un2_pre_out_9 ;
wire un2_pre_out_8 ;
wire un2_pre_out_7 ;
wire un2_pre_out_6 ;
wire un2_pre_out_5 ;
wire un2_pre_out_4 ;
wire un2_pre_out_3 ;
wire un2_pre_out_2 ;
wire un2_pre_out_1 ;
wire un2_pre_out_s_11_0 ;
wire un2_pre_out ;
wire un2_pre_out_axb_1 ;
wire un2_pre_out_axb_2 ;
wire un2_pre_out_axb_3 ;
wire un2_pre_out_axb_4 ;
wire un2_pre_out_axb_5 ;
wire un2_pre_out_axb_6 ;
wire un2_pre_out_axb_7 ;
wire un2_pre_out_axb_8 ;
wire un2_pre_out_axb_9 ;
wire un2_pre_out_axb_10 ;
wire un2_pre_out_axb_11 ;
wire un2_pre_out_cry_10 ;
wire un2_pre_out_cry_9 ;
wire un2_pre_out_cry_8 ;
wire un2_pre_out_cry_7 ;
wire un2_pre_out_cry_6 ;
wire un2_pre_out_cry_5 ;
wire un2_pre_out_cry_4 ;
wire un2_pre_out_cry_3 ;
wire un2_pre_out_cry_2 ;
wire un2_pre_out_cry_1 ;
wire un2_pre_out_cry_0 ;
wire GND ;
wire VCC ;
// instances
  LUT2 un2_pre_out_axb_0(.I0(mult_out_i[0:0]),.I1(out_inner_prod_i[0:0]),.O(un2_pre_out));
defparam un2_pre_out_axb_0.INIT=4'h6;
  LUT2 un2_pre_out_axb_1_cZ(.I0(mult_out_i[1:1]),.I1(out_inner_prod_i[1:1]),.O(un2_pre_out_axb_1));
defparam un2_pre_out_axb_1_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_2_cZ(.I0(mult_out_i[2:2]),.I1(out_inner_prod_i[2:2]),.O(un2_pre_out_axb_2));
defparam un2_pre_out_axb_2_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_3_cZ(.I0(mult_out_i[3:3]),.I1(out_inner_prod_i[3:3]),.O(un2_pre_out_axb_3));
defparam un2_pre_out_axb_3_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_4_cZ(.I0(mult_out_i[4:4]),.I1(out_inner_prod_i[4:4]),.O(un2_pre_out_axb_4));
defparam un2_pre_out_axb_4_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_5_cZ(.I0(mult_out_i[5:5]),.I1(out_inner_prod_i[5:5]),.O(un2_pre_out_axb_5));
defparam un2_pre_out_axb_5_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_6_cZ(.I0(mult_out_i[6:6]),.I1(out_inner_prod_i[6:6]),.O(un2_pre_out_axb_6));
defparam un2_pre_out_axb_6_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_7_cZ(.I0(mult_out_i[7:7]),.I1(out_inner_prod_i[7:7]),.O(un2_pre_out_axb_7));
defparam un2_pre_out_axb_7_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_8_cZ(.I0(mult_out_i[8:8]),.I1(out_inner_prod_i[8:8]),.O(un2_pre_out_axb_8));
defparam un2_pre_out_axb_8_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_9_cZ(.I0(mult_out_i[9:9]),.I1(out_inner_prod_i[9:9]),.O(un2_pre_out_axb_9));
defparam un2_pre_out_axb_9_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_10_cZ(.I0(mult_out_i[10:10]),.I1(out_inner_prod_i[10:10]),.O(un2_pre_out_axb_10));
defparam un2_pre_out_axb_10_cZ.INIT=4'h6;
  LUT2 un2_pre_out_axb_11_cZ(.I0(mult_out_i[11:11]),.I1(out_inner_prod_i[11:11]),.O(un2_pre_out_axb_11));
defparam un2_pre_out_axb_11_cZ.INIT=4'h6;
  XORCY un2_pre_out_s_11(.LI(un2_pre_out_axb_11),.CI(un2_pre_out_cry_10),.O(un2_pre_out_s_11_0));
  XORCY un2_pre_out_s_10(.LI(un2_pre_out_axb_10),.CI(un2_pre_out_cry_9),.O(un2_pre_out_10));
  MUXCY_L un2_pre_out_cry_10_cZ(.DI(mult_out_i[10:10]),.CI(un2_pre_out_cry_9),.S(un2_pre_out_axb_10),.LO(un2_pre_out_cry_10));
  XORCY un2_pre_out_s_9(.LI(un2_pre_out_axb_9),.CI(un2_pre_out_cry_8),.O(un2_pre_out_9));
  MUXCY_L un2_pre_out_cry_9_cZ(.DI(mult_out_i[9:9]),.CI(un2_pre_out_cry_8),.S(un2_pre_out_axb_9),.LO(un2_pre_out_cry_9));
  XORCY un2_pre_out_s_8(.LI(un2_pre_out_axb_8),.CI(un2_pre_out_cry_7),.O(un2_pre_out_8));
  MUXCY_L un2_pre_out_cry_8_cZ(.DI(mult_out_i[8:8]),.CI(un2_pre_out_cry_7),.S(un2_pre_out_axb_8),.LO(un2_pre_out_cry_8));
  XORCY un2_pre_out_s_7(.LI(un2_pre_out_axb_7),.CI(un2_pre_out_cry_6),.O(un2_pre_out_7));
  MUXCY_L un2_pre_out_cry_7_cZ(.DI(mult_out_i[7:7]),.CI(un2_pre_out_cry_6),.S(un2_pre_out_axb_7),.LO(un2_pre_out_cry_7));
  XORCY un2_pre_out_s_6(.LI(un2_pre_out_axb_6),.CI(un2_pre_out_cry_5),.O(un2_pre_out_6));
  MUXCY_L un2_pre_out_cry_6_cZ(.DI(mult_out_i[6:6]),.CI(un2_pre_out_cry_5),.S(un2_pre_out_axb_6),.LO(un2_pre_out_cry_6));
  XORCY un2_pre_out_s_5(.LI(un2_pre_out_axb_5),.CI(un2_pre_out_cry_4),.O(un2_pre_out_5));
  MUXCY_L un2_pre_out_cry_5_cZ(.DI(mult_out_i[5:5]),.CI(un2_pre_out_cry_4),.S(un2_pre_out_axb_5),.LO(un2_pre_out_cry_5));
  XORCY un2_pre_out_s_4(.LI(un2_pre_out_axb_4),.CI(un2_pre_out_cry_3),.O(un2_pre_out_4));
  MUXCY_L un2_pre_out_cry_4_cZ(.DI(mult_out_i[4:4]),.CI(un2_pre_out_cry_3),.S(un2_pre_out_axb_4),.LO(un2_pre_out_cry_4));
  XORCY un2_pre_out_s_3(.LI(un2_pre_out_axb_3),.CI(un2_pre_out_cry_2),.O(un2_pre_out_3));
  MUXCY_L un2_pre_out_cry_3_cZ(.DI(mult_out_i[3:3]),.CI(un2_pre_out_cry_2),.S(un2_pre_out_axb_3),.LO(un2_pre_out_cry_3));
  XORCY un2_pre_out_s_2(.LI(un2_pre_out_axb_2),.CI(un2_pre_out_cry_1),.O(un2_pre_out_2));
  MUXCY_L un2_pre_out_cry_2_cZ(.DI(mult_out_i[2:2]),.CI(un2_pre_out_cry_1),.S(un2_pre_out_axb_2),.LO(un2_pre_out_cry_2));
  XORCY un2_pre_out_s_1(.LI(un2_pre_out_axb_1),.CI(un2_pre_out_cry_0),.O(un2_pre_out_1));
  MUXCY_L un2_pre_out_cry_1_cZ(.DI(mult_out_i[1:1]),.CI(un2_pre_out_cry_0),.S(un2_pre_out_axb_1),.LO(un2_pre_out_cry_1));
  MUXCY_L un2_pre_out_cry_0_cZ(.DI(mult_out_i[0:0]),.CI(GND),.S(un2_pre_out),.LO(un2_pre_out_cry_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module add_subZ1_inj (pre_out_r,in_a_r_reg,in_b_r_reg,mult2_out_0,P_uc_34_0,PATTERNDETECT_7,clk);
output [23:7] pre_out_r ;
input [11:0] in_a_r_reg ;
input [11:0] in_b_r_reg ;
input [23:0] mult2_out_0 ;
input [47:24] P_uc_34_0 ;
output PATTERNDETECT_7 ;
input clk ;
wire PATTERNDETECT_7 ;
wire clk ;
wire [29:0] ACOUT_7 ;
wire [17:0] BCOUT_7 ;
wire [3:0] CARRYOUT_7 ;
wire [6:0] un2_pre_out ;
wire [47:24] P_uc_7 ;
wire [47:0] PCOUT_7 ;
wire CARRYCASCOUT_7 ;
wire MULTSIGNOUT_7 ;
wire OVERFLOW_7 ;
wire PATTERNBDETECT_7 ;
wire UNDERFLOW_7 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc268(.ACOUT(ACOUT_7[29:0]),.BCOUT(BCOUT_7[17:0]),.CARRYCASCOUT(CARRYCASCOUT_7),.CARRYOUT(CARRYOUT_7[3:0]),.MULTSIGNOUT(MULTSIGNOUT_7),.OVERFLOW(OVERFLOW_7),.P({P_uc_7[47:24],pre_out_r[23:7],un2_pre_out[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_7),.PATTERNDETECT(PATTERNDETECT_7),.PCOUT(PCOUT_7[47:0]),.UNDERFLOW(UNDERFLOW_7),.A({in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(VCC),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_34_0[47:24],mult2_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc268.ACASCREG=0;
defparam desc268.ADREG=0;
defparam desc268.ALUMODEREG=0;
defparam desc268.AREG=0;
defparam desc268.AUTORESET_PATDET="NO_RESET";
defparam desc268.A_INPUT="DIRECT";
defparam desc268.BCASCREG=0;
defparam desc268.BREG=0;
defparam desc268.B_INPUT="DIRECT";
defparam desc268.CARRYINREG=0;
defparam desc268.CARRYINSELREG=0;
defparam desc268.CREG=1;
defparam desc268.DREG=0;
defparam desc268.INMODEREG=0;
defparam desc268.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc268.MREG=1;
defparam desc268.OPMODEREG=0;
defparam desc268.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc268.PREG=0;
defparam desc268.SEL_MASK="MASK";
defparam desc268.USE_DPORT="FALSE";
defparam desc268.USE_MULT="MULTIPLY";
defparam desc268.USE_PATTERN_DETECT="PATDET";
defparam desc268.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ1_1_inj (pre_out_i,vec_out_r_AQ_2,in_b_i_reg,mult4_out_0,P_uc_27_0,PATTERNDETECT_3,clk);
output [23:7] pre_out_i ;
input [11:0] vec_out_r_AQ_2 ;
input [11:0] in_b_i_reg ;
input [23:0] mult4_out_0 ;
input [47:24] P_uc_27_0 ;
output PATTERNDETECT_3 ;
input clk ;
wire PATTERNDETECT_3 ;
wire clk ;
wire [29:0] ACOUT_3 ;
wire [17:0] BCOUT_3 ;
wire [3:0] CARRYOUT_3 ;
wire [6:0] un2_pre_out ;
wire [47:24] P_uc_3 ;
wire [47:0] PCOUT_3 ;
wire CARRYCASCOUT_3 ;
wire MULTSIGNOUT_3 ;
wire OVERFLOW_3 ;
wire PATTERNBDETECT_3 ;
wire UNDERFLOW_3 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc480(.ACOUT(ACOUT_3[29:0]),.BCOUT(BCOUT_3[17:0]),.CARRYCASCOUT(CARRYCASCOUT_3),.CARRYOUT(CARRYOUT_3[3:0]),.MULTSIGNOUT(MULTSIGNOUT_3),.OVERFLOW(OVERFLOW_3),.P({P_uc_3[47:24],pre_out_i[23:7],un2_pre_out[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_3),.PATTERNDETECT(PATTERNDETECT_3),.PCOUT(PCOUT_3[47:0]),.UNDERFLOW(UNDERFLOW_3),.A({vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_27_0[47:24],mult4_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc480.ACASCREG=2;
defparam desc480.ADREG=0;
defparam desc480.ALUMODEREG=0;
defparam desc480.AREG=2;
defparam desc480.AUTORESET_PATDET="NO_RESET";
defparam desc480.A_INPUT="DIRECT";
defparam desc480.BCASCREG=1;
defparam desc480.BREG=1;
defparam desc480.B_INPUT="DIRECT";
defparam desc480.CARRYINREG=0;
defparam desc480.CARRYINSELREG=0;
defparam desc480.CREG=1;
defparam desc480.DREG=0;
defparam desc480.INMODEREG=0;
defparam desc480.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc480.MREG=0;
defparam desc480.OPMODEREG=0;
defparam desc480.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc480.PREG=0;
defparam desc480.SEL_MASK="MASK";
defparam desc480.USE_DPORT="FALSE";
defparam desc480.USE_MULT="MULTIPLY";
defparam desc480.USE_PATTERN_DETECT="PATDET";
defparam desc480.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ1_2_inj (pre_out_i,vec_out_r_AQ_1,in_b_i_reg,mult4_out_0,P_uc_23_0,PATTERNDETECT_1,clk);
output [23:7] pre_out_i ;
input [11:0] vec_out_r_AQ_1 ;
input [11:0] in_b_i_reg ;
input [23:0] mult4_out_0 ;
input [47:24] P_uc_23_0 ;
output PATTERNDETECT_1 ;
input clk ;
wire PATTERNDETECT_1 ;
wire clk ;
wire [29:0] ACOUT_1 ;
wire [17:0] BCOUT_1 ;
wire [3:0] CARRYOUT_1 ;
wire [6:0] un2_pre_out ;
wire [47:24] P_uc_1 ;
wire [47:0] PCOUT_1 ;
wire CARRYCASCOUT_1 ;
wire MULTSIGNOUT_1 ;
wire OVERFLOW_1 ;
wire PATTERNBDETECT_1 ;
wire UNDERFLOW_1 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc535(.ACOUT(ACOUT_1[29:0]),.BCOUT(BCOUT_1[17:0]),.CARRYCASCOUT(CARRYCASCOUT_1),.CARRYOUT(CARRYOUT_1[3:0]),.MULTSIGNOUT(MULTSIGNOUT_1),.OVERFLOW(OVERFLOW_1),.P({P_uc_1[47:24],pre_out_i[23:7],un2_pre_out[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_1),.PATTERNDETECT(PATTERNDETECT_1),.PCOUT(PCOUT_1[47:0]),.UNDERFLOW(UNDERFLOW_1),.A({vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_23_0[47:24],mult4_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc535.ACASCREG=2;
defparam desc535.ADREG=0;
defparam desc535.ALUMODEREG=0;
defparam desc535.AREG=2;
defparam desc535.AUTORESET_PATDET="NO_RESET";
defparam desc535.A_INPUT="DIRECT";
defparam desc535.BCASCREG=1;
defparam desc535.BREG=1;
defparam desc535.B_INPUT="DIRECT";
defparam desc535.CARRYINREG=0;
defparam desc535.CARRYINSELREG=0;
defparam desc535.CREG=1;
defparam desc535.DREG=0;
defparam desc535.INMODEREG=0;
defparam desc535.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc535.MREG=0;
defparam desc535.OPMODEREG=0;
defparam desc535.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc535.PREG=0;
defparam desc535.SEL_MASK="MASK";
defparam desc535.USE_DPORT="FALSE";
defparam desc535.USE_MULT="MULTIPLY";
defparam desc535.USE_PATTERN_DETECT="PATDET";
defparam desc535.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ1_3_inj (pre_out_i,vec_out_r_AQ_0,in_b_i_reg,mult4_out_0,P_uc_19_0,PATTERNDETECT,clk);
output [23:7] pre_out_i ;
input [11:0] vec_out_r_AQ_0 ;
input [11:0] in_b_i_reg ;
input [23:0] mult4_out_0 ;
input [47:24] P_uc_19_0 ;
output PATTERNDETECT ;
input clk ;
wire PATTERNDETECT ;
wire clk ;
wire [29:0] ACOUT ;
wire [17:0] BCOUT ;
wire [3:0] CARRYOUT ;
wire [6:0] un2_pre_out ;
wire [47:24] P_uc ;
wire [47:0] PCOUT ;
wire CARRYCASCOUT ;
wire MULTSIGNOUT ;
wire OVERFLOW ;
wire PATTERNBDETECT ;
wire UNDERFLOW ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc590(.ACOUT(ACOUT[29:0]),.BCOUT(BCOUT[17:0]),.CARRYCASCOUT(CARRYCASCOUT),.CARRYOUT(CARRYOUT[3:0]),.MULTSIGNOUT(MULTSIGNOUT),.OVERFLOW(OVERFLOW),.P({P_uc[47:24],pre_out_i[23:7],un2_pre_out[6:0]}),.PATTERNBDETECT(PATTERNBDETECT),.PATTERNDETECT(PATTERNDETECT),.PCOUT(PCOUT[47:0]),.UNDERFLOW(UNDERFLOW),.A({vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_19_0[47:24],mult4_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc590.ACASCREG=2;
defparam desc590.ADREG=0;
defparam desc590.ALUMODEREG=0;
defparam desc590.AREG=2;
defparam desc590.AUTORESET_PATDET="NO_RESET";
defparam desc590.A_INPUT="DIRECT";
defparam desc590.BCASCREG=1;
defparam desc590.BREG=1;
defparam desc590.B_INPUT="DIRECT";
defparam desc590.CARRYINREG=0;
defparam desc590.CARRYINSELREG=0;
defparam desc590.CREG=1;
defparam desc590.DREG=0;
defparam desc590.INMODEREG=0;
defparam desc590.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc590.MREG=0;
defparam desc590.OPMODEREG=0;
defparam desc590.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc590.PREG=0;
defparam desc590.SEL_MASK="MASK";
defparam desc590.USE_DPORT="FALSE";
defparam desc590.USE_MULT="MULTIPLY";
defparam desc590.USE_PATTERN_DETECT="PATDET";
defparam desc590.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ1_4_inj (pre_out_i,vec_out_r_AQ_3,in_b_i_reg,mult4_out_0,P_uc_31_0,PATTERNDETECT_5,clk);
output [23:7] pre_out_i ;
input [11:0] vec_out_r_AQ_3 ;
input [11:0] in_b_i_reg ;
input [23:0] mult4_out_0 ;
input [47:24] P_uc_31_0 ;
output PATTERNDETECT_5 ;
input clk ;
wire PATTERNDETECT_5 ;
wire clk ;
wire [29:0] ACOUT_5 ;
wire [17:0] BCOUT_5 ;
wire [3:0] CARRYOUT_5 ;
wire [6:0] un2_pre_out ;
wire [47:24] P_uc_5 ;
wire [47:0] PCOUT_5 ;
wire CARRYCASCOUT_5 ;
wire MULTSIGNOUT_5 ;
wire OVERFLOW_5 ;
wire PATTERNBDETECT_5 ;
wire UNDERFLOW_5 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc645(.ACOUT(ACOUT_5[29:0]),.BCOUT(BCOUT_5[17:0]),.CARRYCASCOUT(CARRYCASCOUT_5),.CARRYOUT(CARRYOUT_5[3:0]),.MULTSIGNOUT(MULTSIGNOUT_5),.OVERFLOW(OVERFLOW_5),.P({P_uc_5[47:24],pre_out_i[23:7],un2_pre_out[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_5),.PATTERNDETECT(PATTERNDETECT_5),.PCOUT(PCOUT_5[47:0]),.UNDERFLOW(UNDERFLOW_5),.A({vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_31_0[47:24],mult4_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc645.ACASCREG=2;
defparam desc645.ADREG=0;
defparam desc645.ALUMODEREG=0;
defparam desc645.AREG=2;
defparam desc645.AUTORESET_PATDET="NO_RESET";
defparam desc645.A_INPUT="DIRECT";
defparam desc645.BCASCREG=1;
defparam desc645.BREG=1;
defparam desc645.B_INPUT="DIRECT";
defparam desc645.CARRYINREG=0;
defparam desc645.CARRYINSELREG=0;
defparam desc645.CREG=1;
defparam desc645.DREG=0;
defparam desc645.INMODEREG=0;
defparam desc645.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc645.MREG=0;
defparam desc645.OPMODEREG=0;
defparam desc645.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc645.PREG=0;
defparam desc645.SEL_MASK="MASK";
defparam desc645.USE_DPORT="FALSE";
defparam desc645.USE_MULT="MULTIPLY";
defparam desc645.USE_PATTERN_DETECT="PATDET";
defparam desc645.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ2_inj (pre_out_i,in_a_i_reg,in_b_r_reg,mult3_out_0,P_uc_35_0,PATTERNDETECT_8,clk);
output [23:7] pre_out_i ;
input [11:0] in_a_i_reg ;
input [11:0] in_b_r_reg ;
input [23:0] mult3_out_0 ;
input [47:24] P_uc_35_0 ;
output PATTERNDETECT_8 ;
input clk ;
wire PATTERNDETECT_8 ;
wire clk ;
wire [29:0] ACOUT_8 ;
wire [17:0] BCOUT_8 ;
wire [3:0] CARRYOUT_8 ;
wire [6:0] output_Z ;
wire [47:24] P_uc_8 ;
wire [47:0] PCOUT_8 ;
wire CARRYCASCOUT_8 ;
wire MULTSIGNOUT_8 ;
wire OVERFLOW_8 ;
wire PATTERNBDETECT_8 ;
wire UNDERFLOW_8 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc269(.ACOUT(ACOUT_8[29:0]),.BCOUT(BCOUT_8[17:0]),.CARRYCASCOUT(CARRYCASCOUT_8),.CARRYOUT(CARRYOUT_8[3:0]),.MULTSIGNOUT(MULTSIGNOUT_8),.OVERFLOW(OVERFLOW_8),.P({P_uc_8[47:24],pre_out_i[23:7],output_Z[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_8),.PATTERNDETECT(PATTERNDETECT_8),.PCOUT(PCOUT_8[47:0]),.UNDERFLOW(UNDERFLOW_8),.A({in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,VCC,VCC}),.B({in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(VCC),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_35_0[47:24],mult3_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc269.ACASCREG=0;
defparam desc269.ADREG=0;
defparam desc269.ALUMODEREG=0;
defparam desc269.AREG=0;
defparam desc269.AUTORESET_PATDET="NO_RESET";
defparam desc269.A_INPUT="DIRECT";
defparam desc269.BCASCREG=0;
defparam desc269.BREG=0;
defparam desc269.B_INPUT="DIRECT";
defparam desc269.CARRYINREG=0;
defparam desc269.CARRYINSELREG=0;
defparam desc269.CREG=1;
defparam desc269.DREG=0;
defparam desc269.INMODEREG=0;
defparam desc269.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc269.MREG=1;
defparam desc269.OPMODEREG=0;
defparam desc269.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc269.PREG=0;
defparam desc269.SEL_MASK="MASK";
defparam desc269.USE_DPORT="FALSE";
defparam desc269.USE_MULT="MULTIPLY";
defparam desc269.USE_PATTERN_DETECT="PATDET";
defparam desc269.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ2_1_inj (pre_out_r,vec_out_i_AQ_2,in_b_i_reg,mult1_out_0,P_uc_24_0,PATTERNDETECT_4,clk);
output [23:7] pre_out_r ;
input [11:0] vec_out_i_AQ_2 ;
input [11:0] in_b_i_reg ;
input [23:0] mult1_out_0 ;
input [47:24] P_uc_24_0 ;
output PATTERNDETECT_4 ;
input clk ;
wire PATTERNDETECT_4 ;
wire clk ;
wire [29:0] ACOUT_4 ;
wire [17:0] BCOUT_4 ;
wire [3:0] CARRYOUT_4 ;
wire [6:0] output_Z ;
wire [47:24] P_uc_4 ;
wire [47:0] PCOUT_4 ;
wire CARRYCASCOUT_4 ;
wire MULTSIGNOUT_4 ;
wire OVERFLOW_4 ;
wire PATTERNBDETECT_4 ;
wire UNDERFLOW_4 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc479(.ACOUT(ACOUT_4[29:0]),.BCOUT(BCOUT_4[17:0]),.CARRYCASCOUT(CARRYCASCOUT_4),.CARRYOUT(CARRYOUT_4[3:0]),.MULTSIGNOUT(MULTSIGNOUT_4),.OVERFLOW(OVERFLOW_4),.P({P_uc_4[47:24],pre_out_r[23:7],output_Z[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_4),.PATTERNDETECT(PATTERNDETECT_4),.PCOUT(PCOUT_4[47:0]),.UNDERFLOW(UNDERFLOW_4),.A({vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,VCC,VCC}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_24_0[47:24],mult1_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc479.ACASCREG=2;
defparam desc479.ADREG=0;
defparam desc479.ALUMODEREG=0;
defparam desc479.AREG=2;
defparam desc479.AUTORESET_PATDET="NO_RESET";
defparam desc479.A_INPUT="DIRECT";
defparam desc479.BCASCREG=1;
defparam desc479.BREG=1;
defparam desc479.B_INPUT="DIRECT";
defparam desc479.CARRYINREG=0;
defparam desc479.CARRYINSELREG=0;
defparam desc479.CREG=1;
defparam desc479.DREG=0;
defparam desc479.INMODEREG=0;
defparam desc479.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc479.MREG=0;
defparam desc479.OPMODEREG=0;
defparam desc479.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc479.PREG=0;
defparam desc479.SEL_MASK="MASK";
defparam desc479.USE_DPORT="FALSE";
defparam desc479.USE_MULT="MULTIPLY";
defparam desc479.USE_PATTERN_DETECT="PATDET";
defparam desc479.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ2_2_inj (pre_out_r,vec_out_i_AQ_1,in_b_i_reg,mult1_out_0,P_uc_20_0,PATTERNDETECT_2,clk);
output [23:7] pre_out_r ;
input [11:0] vec_out_i_AQ_1 ;
input [11:0] in_b_i_reg ;
input [23:0] mult1_out_0 ;
input [47:24] P_uc_20_0 ;
output PATTERNDETECT_2 ;
input clk ;
wire PATTERNDETECT_2 ;
wire clk ;
wire [29:0] ACOUT_2 ;
wire [17:0] BCOUT_2 ;
wire [3:0] CARRYOUT_2 ;
wire [6:0] output_Z ;
wire [47:24] P_uc_2 ;
wire [47:0] PCOUT_2 ;
wire CARRYCASCOUT_2 ;
wire MULTSIGNOUT_2 ;
wire OVERFLOW_2 ;
wire PATTERNBDETECT_2 ;
wire UNDERFLOW_2 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc534(.ACOUT(ACOUT_2[29:0]),.BCOUT(BCOUT_2[17:0]),.CARRYCASCOUT(CARRYCASCOUT_2),.CARRYOUT(CARRYOUT_2[3:0]),.MULTSIGNOUT(MULTSIGNOUT_2),.OVERFLOW(OVERFLOW_2),.P({P_uc_2[47:24],pre_out_r[23:7],output_Z[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_2),.PATTERNDETECT(PATTERNDETECT_2),.PCOUT(PCOUT_2[47:0]),.UNDERFLOW(UNDERFLOW_2),.A({vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,VCC,VCC}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_20_0[47:24],mult1_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc534.ACASCREG=2;
defparam desc534.ADREG=0;
defparam desc534.ALUMODEREG=0;
defparam desc534.AREG=2;
defparam desc534.AUTORESET_PATDET="NO_RESET";
defparam desc534.A_INPUT="DIRECT";
defparam desc534.BCASCREG=1;
defparam desc534.BREG=1;
defparam desc534.B_INPUT="DIRECT";
defparam desc534.CARRYINREG=0;
defparam desc534.CARRYINSELREG=0;
defparam desc534.CREG=1;
defparam desc534.DREG=0;
defparam desc534.INMODEREG=0;
defparam desc534.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc534.MREG=0;
defparam desc534.OPMODEREG=0;
defparam desc534.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc534.PREG=0;
defparam desc534.SEL_MASK="MASK";
defparam desc534.USE_DPORT="FALSE";
defparam desc534.USE_MULT="MULTIPLY";
defparam desc534.USE_PATTERN_DETECT="PATDET";
defparam desc534.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ2_3_inj (pre_out_r,vec_out_i_AQ_0,in_b_i_reg,mult1_out_0,P_uc_16_0,PATTERNDETECT_0,clk);
output [23:7] pre_out_r ;
input [11:0] vec_out_i_AQ_0 ;
input [11:0] in_b_i_reg ;
input [23:0] mult1_out_0 ;
input [47:24] P_uc_16_0 ;
output PATTERNDETECT_0 ;
input clk ;
wire PATTERNDETECT_0 ;
wire clk ;
wire [29:0] ACOUT_0 ;
wire [17:0] BCOUT_0 ;
wire [3:0] CARRYOUT_0 ;
wire [6:0] output_Z ;
wire [47:24] P_uc_0 ;
wire [47:0] PCOUT_0 ;
wire CARRYCASCOUT_0 ;
wire MULTSIGNOUT_0 ;
wire OVERFLOW_0 ;
wire PATTERNBDETECT_0 ;
wire UNDERFLOW_0 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc589(.ACOUT(ACOUT_0[29:0]),.BCOUT(BCOUT_0[17:0]),.CARRYCASCOUT(CARRYCASCOUT_0),.CARRYOUT(CARRYOUT_0[3:0]),.MULTSIGNOUT(MULTSIGNOUT_0),.OVERFLOW(OVERFLOW_0),.P({P_uc_0[47:24],pre_out_r[23:7],output_Z[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_0),.PATTERNDETECT(PATTERNDETECT_0),.PCOUT(PCOUT_0[47:0]),.UNDERFLOW(UNDERFLOW_0),.A({vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,VCC,VCC}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_16_0[47:24],mult1_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc589.ACASCREG=2;
defparam desc589.ADREG=0;
defparam desc589.ALUMODEREG=0;
defparam desc589.AREG=2;
defparam desc589.AUTORESET_PATDET="NO_RESET";
defparam desc589.A_INPUT="DIRECT";
defparam desc589.BCASCREG=1;
defparam desc589.BREG=1;
defparam desc589.B_INPUT="DIRECT";
defparam desc589.CARRYINREG=0;
defparam desc589.CARRYINSELREG=0;
defparam desc589.CREG=1;
defparam desc589.DREG=0;
defparam desc589.INMODEREG=0;
defparam desc589.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc589.MREG=0;
defparam desc589.OPMODEREG=0;
defparam desc589.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc589.PREG=0;
defparam desc589.SEL_MASK="MASK";
defparam desc589.USE_DPORT="FALSE";
defparam desc589.USE_MULT="MULTIPLY";
defparam desc589.USE_PATTERN_DETECT="PATDET";
defparam desc589.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ2_4_inj (pre_out_r,vec_out_i_AQ_3,in_b_i_reg,mult1_out_0,P_uc_28_0,PATTERNDETECT_6,clk);
output [23:7] pre_out_r ;
input [11:0] vec_out_i_AQ_3 ;
input [11:0] in_b_i_reg ;
input [23:0] mult1_out_0 ;
input [47:24] P_uc_28_0 ;
output PATTERNDETECT_6 ;
input clk ;
wire PATTERNDETECT_6 ;
wire clk ;
wire [29:0] ACOUT_6 ;
wire [17:0] BCOUT_6 ;
wire [3:0] CARRYOUT_6 ;
wire [6:0] output_Z ;
wire [47:24] P_uc_6 ;
wire [47:0] PCOUT_6 ;
wire CARRYCASCOUT_6 ;
wire MULTSIGNOUT_6 ;
wire OVERFLOW_6 ;
wire PATTERNBDETECT_6 ;
wire UNDERFLOW_6 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc644(.ACOUT(ACOUT_6[29:0]),.BCOUT(BCOUT_6[17:0]),.CARRYCASCOUT(CARRYCASCOUT_6),.CARRYOUT(CARRYOUT_6[3:0]),.MULTSIGNOUT(MULTSIGNOUT_6),.OVERFLOW(OVERFLOW_6),.P({P_uc_6[47:24],pre_out_r[23:7],output_Z[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_6),.PATTERNDETECT(PATTERNDETECT_6),.PCOUT(PCOUT_6[47:0]),.UNDERFLOW(UNDERFLOW_6),.A({vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,VCC,VCC}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,VCC,GND,VCC,GND,VCC}),.PCIN({P_uc_28_0[47:24],mult1_out_0[23:0]}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc644.ACASCREG=2;
defparam desc644.ADREG=0;
defparam desc644.ALUMODEREG=0;
defparam desc644.AREG=2;
defparam desc644.AUTORESET_PATDET="NO_RESET";
defparam desc644.A_INPUT="DIRECT";
defparam desc644.BCASCREG=1;
defparam desc644.BREG=1;
defparam desc644.B_INPUT="DIRECT";
defparam desc644.CARRYINREG=0;
defparam desc644.CARRYINSELREG=0;
defparam desc644.CREG=1;
defparam desc644.DREG=0;
defparam desc644.INMODEREG=0;
defparam desc644.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc644.MREG=0;
defparam desc644.OPMODEREG=0;
defparam desc644.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc644.PREG=0;
defparam desc644.SEL_MASK="MASK";
defparam desc644.USE_DPORT="FALSE";
defparam desc644.USE_MULT="MULTIPLY";
defparam desc644.USE_PATTERN_DETECT="PATDET";
defparam desc644.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module add_subZ3_inj (pre_out_10,output_iv_0,output_iv_1,output_iv_9,output_iv_8,output_iv_6,output_iv_7,output_iv_2,output_iv_3,output_iv_4,out_r_vec_mult_0,in_a_r_reg_0,N_500);
output pre_out_10 ;
output output_iv_0 ;
output output_iv_1 ;
output output_iv_9 ;
output output_iv_8 ;
output output_iv_6 ;
output output_iv_7 ;
output output_iv_2 ;
output output_iv_3 ;
output output_iv_4 ;
input [11:0] out_r_vec_mult_0 ;
input [11:0] in_a_r_reg_0 ;
output N_500 ;
wire pre_out_10 ;
wire output_iv_0 ;
wire output_iv_1 ;
wire output_iv_9 ;
wire output_iv_8 ;
wire output_iv_6 ;
wire output_iv_7 ;
wire output_iv_2 ;
wire output_iv_3 ;
wire output_iv_4 ;
wire N_500 ;
wire [10:1] pre_out ;
wire pre_out_i ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 pre_out_axb_0(.I0(out_r_vec_mult_0[0:0]),.I1(in_a_r_reg_0[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_r_vec_mult_0[1:1]),.I1(in_a_r_reg_0[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_r_vec_mult_0[2:2]),.I1(in_a_r_reg_0[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_r_vec_mult_0[3:3]),.I1(in_a_r_reg_0[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_r_vec_mult_0[4:4]),.I1(in_a_r_reg_0[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_r_vec_mult_0[5:5]),.I1(in_a_r_reg_0[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_r_vec_mult_0[6:6]),.I1(in_a_r_reg_0[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_r_vec_mult_0[7:7]),.I1(in_a_r_reg_0[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_r_vec_mult_0[8:8]),.I1(in_a_r_reg_0[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_r_vec_mult_0[9:9]),.I1(in_a_r_reg_0[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_r_vec_mult_0[10:10]),.I1(in_a_r_reg_0[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT2 pre_out_axb_11_cZ(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out[10:10]));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_r_reg_0[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out[9:9]));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_r_reg_0[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out[8:8]));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_r_reg_0[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out[7:7]));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_r_reg_0[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_r_reg_0[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out[5:5]));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_r_reg_0[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_r_reg_0[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out[3:3]));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_r_reg_0[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out[2:2]));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_r_reg_0[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_r_reg_0[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_r_reg_0[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc711(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[5:5]),.I3(pre_out_10),.O(output_iv_4));
defparam desc711.INIT=16'h0D4F;
  LUT4 desc712(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[6:6]),.I3(pre_out_10),.O(N_500));
defparam desc712.INIT=16'h0D4F;
  LUT4 desc713(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[3:3]),.I3(pre_out_10),.O(output_iv_2));
defparam desc713.INIT=16'h0D4F;
  LUT4 desc714(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[4:4]),.I3(pre_out_10),.O(output_iv_3));
defparam desc714.INIT=16'h0D4F;
  LUT4 desc715(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[7:7]),.I3(pre_out_10),.O(output_iv_6));
defparam desc715.INIT=16'h0D4F;
  LUT4 desc716(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[8:8]),.I3(pre_out_10),.O(output_iv_7));
defparam desc716.INIT=16'h0D4F;
  LUT4 desc717(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[10:10]),.I3(pre_out_10),.O(output_iv_9));
defparam desc717.INIT=16'h0D4F;
  LUT4 desc718(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[9:9]),.I3(pre_out_10),.O(output_iv_8));
defparam desc718.INIT=16'h0D4F;
  LUT4 desc719(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[1:1]),.I3(pre_out_10),.O(output_iv_0));
defparam desc719.INIT=16'h0D4F;
  LUT4 desc720(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0[11:11]),.I2(pre_out[2:2]),.I3(pre_out_10),.O(output_iv_1));
defparam desc720.INIT=16'h0D4F;
endmodule
module add_subZ3_1_inj (pre_out_i_m_8,pre_out_i_m_4,pre_out_i_m_0,out_r_vec_mult_1,in_a_r_reg_1,pre_out_10,pre_out_9,pre_out_8,pre_out_6,pre_out_5,pre_out_4,pre_out_2,pre_out_1,pre_out_0,un5_output);
output pre_out_i_m_8 ;
output pre_out_i_m_4 ;
output pre_out_i_m_0 ;
input [11:0] out_r_vec_mult_1 ;
input [11:0] in_a_r_reg_1 ;
output pre_out_10 ;
output pre_out_9 ;
output pre_out_8 ;
output pre_out_6 ;
output pre_out_5 ;
output pre_out_4 ;
output pre_out_2 ;
output pre_out_1 ;
output pre_out_0 ;
output un5_output ;
wire pre_out_i_m_8 ;
wire pre_out_i_m_4 ;
wire pre_out_i_m_0 ;
wire pre_out_10 ;
wire pre_out_9 ;
wire pre_out_8 ;
wire pre_out_6 ;
wire pre_out_5 ;
wire pre_out_4 ;
wire pre_out_2 ;
wire pre_out_1 ;
wire pre_out_0 ;
wire un5_output ;
wire [8:4] pre_out ;
wire pre_out_i ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 pre_out_axb_0(.I0(out_r_vec_mult_1[0:0]),.I1(in_a_r_reg_1[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_r_vec_mult_1[1:1]),.I1(in_a_r_reg_1[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_r_vec_mult_1[2:2]),.I1(in_a_r_reg_1[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_r_vec_mult_1[3:3]),.I1(in_a_r_reg_1[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_r_vec_mult_1[4:4]),.I1(in_a_r_reg_1[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_r_vec_mult_1[5:5]),.I1(in_a_r_reg_1[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_r_vec_mult_1[6:6]),.I1(in_a_r_reg_1[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_r_vec_mult_1[7:7]),.I1(in_a_r_reg_1[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_r_vec_mult_1[8:8]),.I1(in_a_r_reg_1[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_r_vec_mult_1[9:9]),.I1(in_a_r_reg_1[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_r_vec_mult_1[10:10]),.I1(in_a_r_reg_1[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT2 pre_out_axb_11_cZ(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out_9));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_r_reg_1[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out_8));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_r_reg_1[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out[8:8]));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_r_reg_1[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out_6));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_r_reg_1[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out_5));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_r_reg_1[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out_4));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_r_reg_1[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_r_reg_1[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out_2));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_r_reg_1[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out_1));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_r_reg_1[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out_0));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_r_reg_1[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_r_reg_1[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 desc721(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(pre_out_10),.O(un5_output));
defparam desc721.INIT=8'hFB;
  LUT5 desc722(.I0(out_r_vec_mult_1[0:0]),.I1(in_a_r_reg_1[0:0]),.I2(out_r_vec_mult_1[11:11]),.I3(in_a_r_reg_1[11:11]),.I4(pre_out_10),.O(pre_out_i_m_0));
defparam desc722.INIT=32'h99099099;
  LUT4 pre_out_s_4_RNIDBUP_o6(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(pre_out[8:8]),.I3(pre_out_10),.O(pre_out_i_m_8));
defparam pre_out_s_4_RNIDBUP_o6.INIT=16'h0D0B;
  LUT4 pre_out_s_4_RNIDBUP_o5(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(pre_out[4:4]),.I3(pre_out_10),.O(pre_out_i_m_4));
defparam pre_out_s_4_RNIDBUP_o5.INIT=16'h0D0B;
endmodule
module add_subZ3_2_inj (out_r_vec_mult_2,in_a_r_reg_2,pre_out_i_m_6,pre_out_i_m_0,pre_out_10,pre_out_9,pre_out_8,pre_out_7,pre_out_6,pre_out_4,pre_out_3,pre_out_2,pre_out_1,pre_out_0,un5_output);
input [11:0] out_r_vec_mult_2 ;
input [11:0] in_a_r_reg_2 ;
output pre_out_i_m_6 ;
output pre_out_i_m_0 ;
output pre_out_10 ;
output pre_out_9 ;
output pre_out_8 ;
output pre_out_7 ;
output pre_out_6 ;
output pre_out_4 ;
output pre_out_3 ;
output pre_out_2 ;
output pre_out_1 ;
output pre_out_0 ;
output un5_output ;
wire pre_out_i_m_6 ;
wire pre_out_i_m_0 ;
wire pre_out_10 ;
wire pre_out_9 ;
wire pre_out_8 ;
wire pre_out_7 ;
wire pre_out_6 ;
wire pre_out_4 ;
wire pre_out_3 ;
wire pre_out_2 ;
wire pre_out_1 ;
wire pre_out_0 ;
wire un5_output ;
wire [6:6] pre_out ;
wire pre_out_i ;
wire GND ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
// instances
  LUT2 pre_out_axb_0(.I0(out_r_vec_mult_2[0:0]),.I1(in_a_r_reg_2[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_r_vec_mult_2[1:1]),.I1(in_a_r_reg_2[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_r_vec_mult_2[2:2]),.I1(in_a_r_reg_2[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_r_vec_mult_2[3:3]),.I1(in_a_r_reg_2[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_r_vec_mult_2[4:4]),.I1(in_a_r_reg_2[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_r_vec_mult_2[5:5]),.I1(in_a_r_reg_2[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_r_vec_mult_2[6:6]),.I1(in_a_r_reg_2[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_r_vec_mult_2[7:7]),.I1(in_a_r_reg_2[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_r_vec_mult_2[8:8]),.I1(in_a_r_reg_2[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_r_vec_mult_2[9:9]),.I1(in_a_r_reg_2[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_r_vec_mult_2[10:10]),.I1(in_a_r_reg_2[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT5 pre_out_s_11_RNI16U11(.I0(out_r_vec_mult_2[0:0]),.I1(in_a_r_reg_2[0:0]),.I2(out_r_vec_mult_2[11:11]),.I3(in_a_r_reg_2[11:11]),.I4(pre_out_10),.O(pre_out_i_m_0));
defparam pre_out_s_11_RNI16U11.INIT=32'h99099099;
  LUT2 pre_out_axb_11_cZ(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out_9));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_r_reg_2[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out_8));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_r_reg_2[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out_7));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_r_reg_2[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out_6));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_r_reg_2[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_r_reg_2[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out_4));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_r_reg_2[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out_3));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_r_reg_2[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out_2));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_r_reg_2[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out_1));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_r_reg_2[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out_0));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_r_reg_2[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_r_reg_2[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT4 pre_out_s_6_RNIRQ081_o6(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(pre_out[6:6]),.I3(pre_out_10),.O(pre_out_i_m_6));
defparam pre_out_s_6_RNIRQ081_o6.INIT=16'h0D0B;
  LUT3 pre_out_s_6_RNIRQ081_o5(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(pre_out_10),.O(un5_output));
defparam pre_out_s_6_RNIRQ081_o5.INIT=8'hFB;
endmodule
module add_subZ3_3_inj (out_r_vec_mult_3,in_a_r_reg_3,pre_out_i_m,pre_out_10,pre_out_9,pre_out_8,pre_out_7,pre_out_6,pre_out_5,pre_out_4,pre_out_3,pre_out_2,pre_out_1,un5_output);
input [11:0] out_r_vec_mult_3 ;
input [11:0] in_a_r_reg_3 ;
output [1:0] pre_out_i_m ;
output pre_out_10 ;
output pre_out_9 ;
output pre_out_8 ;
output pre_out_7 ;
output pre_out_6 ;
output pre_out_5 ;
output pre_out_4 ;
output pre_out_3 ;
output pre_out_2 ;
output pre_out_1 ;
output un5_output ;
wire pre_out_10 ;
wire pre_out_9 ;
wire pre_out_8 ;
wire pre_out_7 ;
wire pre_out_6 ;
wire pre_out_5 ;
wire pre_out_4 ;
wire pre_out_3 ;
wire pre_out_2 ;
wire pre_out_1 ;
wire un5_output ;
wire [1:1] pre_out ;
wire pre_out_i ;
wire GND ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
// instances
  LUT2 pre_out_axb_0(.I0(out_r_vec_mult_3[0:0]),.I1(in_a_r_reg_3[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_r_vec_mult_3[1:1]),.I1(in_a_r_reg_3[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_r_vec_mult_3[2:2]),.I1(in_a_r_reg_3[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_r_vec_mult_3[3:3]),.I1(in_a_r_reg_3[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_r_vec_mult_3[4:4]),.I1(in_a_r_reg_3[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_r_vec_mult_3[5:5]),.I1(in_a_r_reg_3[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_r_vec_mult_3[6:6]),.I1(in_a_r_reg_3[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_r_vec_mult_3[7:7]),.I1(in_a_r_reg_3[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_r_vec_mult_3[8:8]),.I1(in_a_r_reg_3[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_r_vec_mult_3[9:9]),.I1(in_a_r_reg_3[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_r_vec_mult_3[10:10]),.I1(in_a_r_reg_3[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT5 pre_out_s_11_RNI6TNU(.I0(out_r_vec_mult_3[0:0]),.I1(in_a_r_reg_3[0:0]),.I2(out_r_vec_mult_3[11:11]),.I3(in_a_r_reg_3[11:11]),.I4(pre_out_10),.O(pre_out_i_m[0:0]));
defparam pre_out_s_11_RNI6TNU.INIT=32'h99099099;
  LUT2 pre_out_axb_11_cZ(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out_9));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_r_reg_3[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out_8));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_r_reg_3[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out_7));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_r_reg_3[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out_6));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_r_reg_3[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out_5));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_r_reg_3[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out_4));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_r_reg_3[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out_3));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_r_reg_3[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out_2));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_r_reg_3[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out_1));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_r_reg_3[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_r_reg_3[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_r_reg_3[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT4 pre_out_s_1_RNIQIL91_o6(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(pre_out[1:1]),.I3(pre_out_10),.O(pre_out_i_m[1:1]));
defparam pre_out_s_1_RNIQIL91_o6.INIT=16'h0D0B;
  LUT3 pre_out_s_1_RNIQIL91_o5(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(pre_out_10),.O(un5_output));
defparam pre_out_s_1_RNIQIL91_o5.INIT=8'hFB;
endmodule
module add_subZ3_4_inj (pre_out_10,output_iv,out_i_vec_sub_0,out_i_vec_mult_0,in_a_i_reg_0);
output pre_out_10 ;
output [10:0] output_iv ;
output [11:11] out_i_vec_sub_0 ;
input [11:0] out_i_vec_mult_0 ;
input [11:0] in_a_i_reg_0 ;
wire pre_out_10 ;
wire [10:1] pre_out ;
wire pre_out_i ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 pre_out_axb_0(.I0(out_i_vec_mult_0[0:0]),.I1(in_a_i_reg_0[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_i_vec_mult_0[1:1]),.I1(in_a_i_reg_0[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_i_vec_mult_0[2:2]),.I1(in_a_i_reg_0[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_i_vec_mult_0[3:3]),.I1(in_a_i_reg_0[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_i_vec_mult_0[4:4]),.I1(in_a_i_reg_0[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_i_vec_mult_0[5:5]),.I1(in_a_i_reg_0[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_i_vec_mult_0[6:6]),.I1(in_a_i_reg_0[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_i_vec_mult_0[7:7]),.I1(in_a_i_reg_0[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_i_vec_mult_0[8:8]),.I1(in_a_i_reg_0[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_i_vec_mult_0[9:9]),.I1(in_a_i_reg_0[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_i_vec_mult_0[10:10]),.I1(in_a_i_reg_0[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT2 pre_out_axb_11_cZ(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out[10:10]));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_i_reg_0[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out[9:9]));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_i_reg_0[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out[8:8]));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_i_reg_0[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out[7:7]));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_i_reg_0[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_i_reg_0[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out[5:5]));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_i_reg_0[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_i_reg_0[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out[3:3]));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_i_reg_0[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out[2:2]));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_i_reg_0[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_i_reg_0[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_i_reg_0[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT5 desc723(.I0(out_i_vec_mult_0[0:0]),.I1(in_a_i_reg_0[0:0]),.I2(out_i_vec_mult_0[11:11]),.I3(in_a_i_reg_0[11:11]),.I4(pre_out_10),.O(output_iv[0:0]));
defparam desc723.INIT=32'h99099F99;
  LUT3 desc724(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out_10),.O(out_i_vec_sub_0[11:11]));
defparam desc724.INIT=8'hD4;
  LUT4 desc725(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[2:2]),.I3(pre_out_10),.O(output_iv[2:2]));
defparam desc725.INIT=16'h0D4F;
  LUT4 desc726(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[3:3]),.I3(pre_out_10),.O(output_iv[3:3]));
defparam desc726.INIT=16'h0D4F;
  LUT4 desc727(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[4:4]),.I3(pre_out_10),.O(output_iv[4:4]));
defparam desc727.INIT=16'h0D4F;
  LUT4 desc728(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[1:1]),.I3(pre_out_10),.O(output_iv[1:1]));
defparam desc728.INIT=16'h0D4F;
  LUT4 desc729(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[10:10]),.I3(pre_out_10),.O(output_iv[10:10]));
defparam desc729.INIT=16'h0D4F;
  LUT4 desc730(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[9:9]),.I3(pre_out_10),.O(output_iv[9:9]));
defparam desc730.INIT=16'h0D4F;
  LUT4 desc731(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[5:5]),.I3(pre_out_10),.O(output_iv[5:5]));
defparam desc731.INIT=16'h0D4F;
  LUT4 desc732(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[6:6]),.I3(pre_out_10),.O(output_iv[6:6]));
defparam desc732.INIT=16'h0D4F;
  LUT4 desc733(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[8:8]),.I3(pre_out_10),.O(output_iv[8:8]));
defparam desc733.INIT=16'h0D4F;
  LUT4 desc734(.I0(out_i_vec_mult_0[11:11]),.I1(in_a_i_reg_0[11:11]),.I2(pre_out[7:7]),.I3(pre_out_10),.O(output_iv[7:7]));
defparam desc734.INIT=16'h0D4F;
endmodule
module add_subZ3_5_inj (pre_out_i_m,out_i_vec_mult_1,in_a_i_reg_1,pre_out,un5_output);
output pre_out_i_m ;
input [11:0] out_i_vec_mult_1 ;
input [11:0] in_a_i_reg_1 ;
output [11:1] pre_out ;
output un5_output ;
wire un5_output ;
wire pre_out_i ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 pre_out_axb_0(.I0(out_i_vec_mult_1[0:0]),.I1(in_a_i_reg_1[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_i_vec_mult_1[1:1]),.I1(in_a_i_reg_1[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_i_vec_mult_1[2:2]),.I1(in_a_i_reg_1[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_i_vec_mult_1[3:3]),.I1(in_a_i_reg_1[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_i_vec_mult_1[4:4]),.I1(in_a_i_reg_1[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_i_vec_mult_1[5:5]),.I1(in_a_i_reg_1[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_i_vec_mult_1[6:6]),.I1(in_a_i_reg_1[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_i_vec_mult_1[7:7]),.I1(in_a_i_reg_1[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_i_vec_mult_1[8:8]),.I1(in_a_i_reg_1[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_i_vec_mult_1[9:9]),.I1(in_a_i_reg_1[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_i_vec_mult_1[10:10]),.I1(in_a_i_reg_1[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT2 pre_out_axb_11_cZ(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out[11:11]));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out[10:10]));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_i_reg_1[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out[9:9]));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_i_reg_1[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out[8:8]));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_i_reg_1[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out[7:7]));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_i_reg_1[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_i_reg_1[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out[5:5]));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_i_reg_1[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_i_reg_1[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out[3:3]));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_i_reg_1[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out[2:2]));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_i_reg_1[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_i_reg_1[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_i_reg_1[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 desc735(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(pre_out[11:11]),.O(un5_output));
defparam desc735.INIT=8'hFB;
  LUT5 desc736(.I0(out_i_vec_mult_1[0:0]),.I1(in_a_i_reg_1[0:0]),.I2(out_i_vec_mult_1[11:11]),.I3(in_a_i_reg_1[11:11]),.I4(pre_out[11:11]),.O(pre_out_i_m));
defparam desc736.INIT=32'h99099099;
endmodule
module add_subZ3_6_inj (pre_out_i_m,out_i_vec_mult_2,in_a_i_reg_2,pre_out,un5_output);
output pre_out_i_m ;
input [11:0] out_i_vec_mult_2 ;
input [11:0] in_a_i_reg_2 ;
output [11:1] pre_out ;
output un5_output ;
wire un5_output ;
wire pre_out_i ;
wire VCC ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
wire GND ;
// instances
  LUT2 pre_out_axb_0(.I0(out_i_vec_mult_2[0:0]),.I1(in_a_i_reg_2[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_i_vec_mult_2[1:1]),.I1(in_a_i_reg_2[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_i_vec_mult_2[2:2]),.I1(in_a_i_reg_2[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_i_vec_mult_2[3:3]),.I1(in_a_i_reg_2[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_i_vec_mult_2[4:4]),.I1(in_a_i_reg_2[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_i_vec_mult_2[5:5]),.I1(in_a_i_reg_2[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_i_vec_mult_2[6:6]),.I1(in_a_i_reg_2[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_i_vec_mult_2[7:7]),.I1(in_a_i_reg_2[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_i_vec_mult_2[8:8]),.I1(in_a_i_reg_2[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_i_vec_mult_2[9:9]),.I1(in_a_i_reg_2[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_i_vec_mult_2[10:10]),.I1(in_a_i_reg_2[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT2 pre_out_axb_11_cZ(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out[11:11]));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out[10:10]));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_i_reg_2[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out[9:9]));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_i_reg_2[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out[8:8]));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_i_reg_2[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out[7:7]));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_i_reg_2[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_i_reg_2[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out[5:5]));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_i_reg_2[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_i_reg_2[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out[3:3]));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_i_reg_2[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out[2:2]));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_i_reg_2[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_i_reg_2[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_i_reg_2[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 desc737(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(pre_out[11:11]),.O(un5_output));
defparam desc737.INIT=8'hFB;
  LUT5 desc738(.I0(out_i_vec_mult_2[0:0]),.I1(in_a_i_reg_2[0:0]),.I2(out_i_vec_mult_2[11:11]),.I3(in_a_i_reg_2[11:11]),.I4(pre_out[11:11]),.O(pre_out_i_m));
defparam desc738.INIT=32'h99099099;
endmodule
module add_subZ3_7_inj (out_i_vec_mult_3,in_a_i_reg_3,pre_out_i_m_1,pre_out_i_m_5,pre_out_i_m_2,pre_out_i_m_10,pre_out_i_m_9,pre_out_i_m_6,pre_out_i_m_7,pre_out_i_m_3,pre_out_i_m_4,pre_out_i_m_0,pre_out_10,pre_out_7,un5_output);
input [11:0] out_i_vec_mult_3 ;
input [11:0] in_a_i_reg_3 ;
output pre_out_i_m_1 ;
output pre_out_i_m_5 ;
output pre_out_i_m_2 ;
output pre_out_i_m_10 ;
output pre_out_i_m_9 ;
output pre_out_i_m_6 ;
output pre_out_i_m_7 ;
output pre_out_i_m_3 ;
output pre_out_i_m_4 ;
output pre_out_i_m_0 ;
output pre_out_10 ;
output pre_out_7 ;
output un5_output ;
wire pre_out_i_m_1 ;
wire pre_out_i_m_5 ;
wire pre_out_i_m_2 ;
wire pre_out_i_m_10 ;
wire pre_out_i_m_9 ;
wire pre_out_i_m_6 ;
wire pre_out_i_m_7 ;
wire pre_out_i_m_3 ;
wire pre_out_i_m_4 ;
wire pre_out_i_m_0 ;
wire pre_out_10 ;
wire pre_out_7 ;
wire un5_output ;
wire [10:1] pre_out ;
wire pre_out_i ;
wire VCC ;
wire GND ;
wire pre_out_axb_1 ;
wire pre_out_axb_2 ;
wire pre_out_axb_3 ;
wire pre_out_axb_4 ;
wire pre_out_axb_5 ;
wire pre_out_axb_6 ;
wire pre_out_axb_7 ;
wire pre_out_axb_8 ;
wire pre_out_axb_9 ;
wire pre_out_axb_10 ;
wire pre_out_axb_11 ;
wire pre_out_cry_10 ;
wire pre_out_cry_9 ;
wire pre_out_cry_8 ;
wire pre_out_cry_7 ;
wire pre_out_cry_6 ;
wire pre_out_cry_5 ;
wire pre_out_cry_4 ;
wire pre_out_cry_3 ;
wire pre_out_cry_2 ;
wire pre_out_cry_1 ;
wire pre_out_cry_0 ;
// instances
  LUT2 pre_out_axb_0(.I0(out_i_vec_mult_3[0:0]),.I1(in_a_i_reg_3[0:0]),.O(pre_out_i));
defparam pre_out_axb_0.INIT=4'h9;
  LUT2 pre_out_axb_1_cZ(.I0(out_i_vec_mult_3[1:1]),.I1(in_a_i_reg_3[1:1]),.O(pre_out_axb_1));
defparam pre_out_axb_1_cZ.INIT=4'h9;
  LUT2 pre_out_axb_2_cZ(.I0(out_i_vec_mult_3[2:2]),.I1(in_a_i_reg_3[2:2]),.O(pre_out_axb_2));
defparam pre_out_axb_2_cZ.INIT=4'h9;
  LUT2 pre_out_axb_3_cZ(.I0(out_i_vec_mult_3[3:3]),.I1(in_a_i_reg_3[3:3]),.O(pre_out_axb_3));
defparam pre_out_axb_3_cZ.INIT=4'h9;
  LUT2 pre_out_axb_4_cZ(.I0(out_i_vec_mult_3[4:4]),.I1(in_a_i_reg_3[4:4]),.O(pre_out_axb_4));
defparam pre_out_axb_4_cZ.INIT=4'h9;
  LUT2 pre_out_axb_5_cZ(.I0(out_i_vec_mult_3[5:5]),.I1(in_a_i_reg_3[5:5]),.O(pre_out_axb_5));
defparam pre_out_axb_5_cZ.INIT=4'h9;
  LUT2 pre_out_axb_6_cZ(.I0(out_i_vec_mult_3[6:6]),.I1(in_a_i_reg_3[6:6]),.O(pre_out_axb_6));
defparam pre_out_axb_6_cZ.INIT=4'h9;
  LUT2 pre_out_axb_7_cZ(.I0(out_i_vec_mult_3[7:7]),.I1(in_a_i_reg_3[7:7]),.O(pre_out_axb_7));
defparam pre_out_axb_7_cZ.INIT=4'h9;
  LUT2 pre_out_axb_8_cZ(.I0(out_i_vec_mult_3[8:8]),.I1(in_a_i_reg_3[8:8]),.O(pre_out_axb_8));
defparam pre_out_axb_8_cZ.INIT=4'h9;
  LUT2 pre_out_axb_9_cZ(.I0(out_i_vec_mult_3[9:9]),.I1(in_a_i_reg_3[9:9]),.O(pre_out_axb_9));
defparam pre_out_axb_9_cZ.INIT=4'h9;
  LUT2 pre_out_axb_10_cZ(.I0(out_i_vec_mult_3[10:10]),.I1(in_a_i_reg_3[10:10]),.O(pre_out_axb_10));
defparam pre_out_axb_10_cZ.INIT=4'h9;
  LUT5 pre_out_s_11_RNIPS481(.I0(out_i_vec_mult_3[0:0]),.I1(in_a_i_reg_3[0:0]),.I2(out_i_vec_mult_3[11:11]),.I3(in_a_i_reg_3[11:11]),.I4(pre_out_10),.O(pre_out_i_m_0));
defparam pre_out_s_11_RNIPS481.INIT=32'h99099099;
  LUT2 pre_out_axb_11_cZ(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.O(pre_out_axb_11));
defparam pre_out_axb_11_cZ.INIT=4'h9;
  XORCY pre_out_s_11(.LI(pre_out_axb_11),.CI(pre_out_cry_10),.O(pre_out_10));
  XORCY pre_out_s_10(.LI(pre_out_axb_10),.CI(pre_out_cry_9),.O(pre_out[10:10]));
  MUXCY_L pre_out_cry_10_cZ(.DI(in_a_i_reg_3[10:10]),.CI(pre_out_cry_9),.S(pre_out_axb_10),.LO(pre_out_cry_10));
  XORCY pre_out_s_9(.LI(pre_out_axb_9),.CI(pre_out_cry_8),.O(pre_out[9:9]));
  MUXCY_L pre_out_cry_9_cZ(.DI(in_a_i_reg_3[9:9]),.CI(pre_out_cry_8),.S(pre_out_axb_9),.LO(pre_out_cry_9));
  XORCY pre_out_s_8(.LI(pre_out_axb_8),.CI(pre_out_cry_7),.O(pre_out_7));
  MUXCY_L pre_out_cry_8_cZ(.DI(in_a_i_reg_3[8:8]),.CI(pre_out_cry_7),.S(pre_out_axb_8),.LO(pre_out_cry_8));
  XORCY pre_out_s_7(.LI(pre_out_axb_7),.CI(pre_out_cry_6),.O(pre_out[7:7]));
  MUXCY_L pre_out_cry_7_cZ(.DI(in_a_i_reg_3[7:7]),.CI(pre_out_cry_6),.S(pre_out_axb_7),.LO(pre_out_cry_7));
  XORCY pre_out_s_6(.LI(pre_out_axb_6),.CI(pre_out_cry_5),.O(pre_out[6:6]));
  MUXCY_L pre_out_cry_6_cZ(.DI(in_a_i_reg_3[6:6]),.CI(pre_out_cry_5),.S(pre_out_axb_6),.LO(pre_out_cry_6));
  XORCY pre_out_s_5(.LI(pre_out_axb_5),.CI(pre_out_cry_4),.O(pre_out[5:5]));
  MUXCY_L pre_out_cry_5_cZ(.DI(in_a_i_reg_3[5:5]),.CI(pre_out_cry_4),.S(pre_out_axb_5),.LO(pre_out_cry_5));
  XORCY pre_out_s_4(.LI(pre_out_axb_4),.CI(pre_out_cry_3),.O(pre_out[4:4]));
  MUXCY_L pre_out_cry_4_cZ(.DI(in_a_i_reg_3[4:4]),.CI(pre_out_cry_3),.S(pre_out_axb_4),.LO(pre_out_cry_4));
  XORCY pre_out_s_3(.LI(pre_out_axb_3),.CI(pre_out_cry_2),.O(pre_out[3:3]));
  MUXCY_L pre_out_cry_3_cZ(.DI(in_a_i_reg_3[3:3]),.CI(pre_out_cry_2),.S(pre_out_axb_3),.LO(pre_out_cry_3));
  XORCY pre_out_s_2(.LI(pre_out_axb_2),.CI(pre_out_cry_1),.O(pre_out[2:2]));
  MUXCY_L pre_out_cry_2_cZ(.DI(in_a_i_reg_3[2:2]),.CI(pre_out_cry_1),.S(pre_out_axb_2),.LO(pre_out_cry_2));
  XORCY pre_out_s_1(.LI(pre_out_axb_1),.CI(pre_out_cry_0),.O(pre_out[1:1]));
  MUXCY_L pre_out_cry_1_cZ(.DI(in_a_i_reg_3[1:1]),.CI(pre_out_cry_0),.S(pre_out_axb_1),.LO(pre_out_cry_1));
  MUXCY_L pre_out_cry_0_cZ(.DI(in_a_i_reg_3[0:0]),.CI(VCC),.S(pre_out_i),.LO(pre_out_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 pre_out_s_3_RNI5JVQ1_o6(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[3:3]),.I3(pre_out_10),.O(pre_out_i_m_3));
defparam pre_out_s_3_RNI5JVQ1_o6.INIT=16'h0D0B;
  LUT4 pre_out_s_3_RNI5JVQ1_o5(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[4:4]),.I3(pre_out_10),.O(pre_out_i_m_4));
defparam pre_out_s_3_RNI5JVQ1_o5.INIT=16'h0D0B;
  LUT4 pre_out_s_6_RNIBJVQ1_o6(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[6:6]),.I3(pre_out_10),.O(pre_out_i_m_6));
defparam pre_out_s_6_RNIBJVQ1_o6.INIT=16'h0D0B;
  LUT4 pre_out_s_6_RNIBJVQ1_o5(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[7:7]),.I3(pre_out_10),.O(pre_out_i_m_7));
defparam pre_out_s_6_RNIBJVQ1_o5.INIT=16'h0D0B;
  LUT4 pre_out_s_9_RNIOUVQ1_o6(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[10:10]),.I3(pre_out_10),.O(pre_out_i_m_10));
defparam pre_out_s_9_RNIOUVQ1_o6.INIT=16'h0D0B;
  LUT4 pre_out_s_9_RNIOUVQ1_o5(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[9:9]),.I3(pre_out_10),.O(pre_out_i_m_9));
defparam pre_out_s_9_RNIOUVQ1_o5.INIT=16'h0D0B;
  LUT4 pre_out_s_2_RNINIFC1_o6(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[2:2]),.I3(pre_out_10),.O(pre_out_i_m_2));
defparam pre_out_s_2_RNINIFC1_o6.INIT=16'h0D0B;
  LUT3 pre_out_s_2_RNINIFC1_o5(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out_10),.O(un5_output));
defparam pre_out_s_2_RNINIFC1_o5.INIT=8'hFB;
  LUT4 pre_out_s_1_RNI4JVQ1_o6(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[1:1]),.I3(pre_out_10),.O(pre_out_i_m_1));
defparam pre_out_s_1_RNI4JVQ1_o6.INIT=16'h0D0B;
  LUT4 pre_out_s_1_RNI4JVQ1_o5(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(pre_out[5:5]),.I3(pre_out_10),.O(pre_out_i_m_5));
defparam pre_out_s_1_RNI4JVQ1_o5.INIT=16'h0D0B;
endmodule
module complex_mult_pipe_prod_inj (mult_out_r,mult_out_i,in_a_r_reg,in_b_r_reg,in_a_i_reg,in_b_i_reg,clk);
output [11:0] mult_out_r ;
output [11:0] mult_out_i ;
input [11:0] in_a_r_reg ;
input [11:0] in_b_r_reg ;
input [11:0] in_a_i_reg ;
input [11:0] in_b_i_reg ;
input clk ;
wire clk ;
wire [23:7] pre_out_i ;
wire [23:7] pre_out_r ;
wire [23:23] mult2_out ;
wire [23:23] mult1_out ;
wire [23:23] mult3_out ;
wire [23:23] mult4_out ;
wire [11:11] pos_out_r ;
wire [11:11] pos_out_i ;
wire [10:0] un7_rnd_out_r ;
wire [10:0] pos_out_r_iv_i ;
wire [10:0] un5_rnd_out_i ;
wire [10:0] pos_out_i_iv_i ;
wire [23:0] mult2_out_0 ;
wire [47:24] P_uc_34_0 ;
wire [23:0] mult3_out_0 ;
wire [47:24] P_uc_35_0 ;
wire un5_rnd_out_i_axb_1 ;
wire un5_rnd_out_i_axb_2 ;
wire un5_rnd_out_i_axb_3 ;
wire un5_rnd_out_i_axb_4 ;
wire un5_rnd_out_i_axb_5 ;
wire un5_rnd_out_i_axb_6 ;
wire un5_rnd_out_i_axb_7 ;
wire un5_rnd_out_i_axb_8 ;
wire un5_rnd_out_i_axb_9 ;
wire un5_rnd_out_i_axb_10 ;
wire un5_rnd_out_i_axb_11 ;
wire un7_rnd_out_r_axb_1 ;
wire un7_rnd_out_r_axb_2 ;
wire un7_rnd_out_r_axb_3 ;
wire un7_rnd_out_r_axb_4 ;
wire un7_rnd_out_r_axb_5 ;
wire un7_rnd_out_r_axb_6 ;
wire un7_rnd_out_r_axb_7 ;
wire un7_rnd_out_r_axb_8 ;
wire un7_rnd_out_r_axb_9 ;
wire un7_rnd_out_r_axb_10 ;
wire un7_rnd_out_r_axb_11 ;
wire un7_rnd_out_r_axb_12 ;
wire un5_rnd_out_i_axb_12 ;
wire un4_rnd_sat_out_i_3 ;
wire un5_rnd_sat_out_r_3 ;
wire un1_pos_out_r_3 ;
wire un1_pos_out_i_3 ;
wire PATTERNDETECT_7 ;
wire un7_rnd_out_r_s_12 ;
wire PATTERNDETECT_8 ;
wire un5_rnd_out_i_s_12 ;
wire un7_rnd_out_r_cry_11 ;
wire un7_rnd_out_r_cry_10 ;
wire GND ;
wire un7_rnd_out_r_cry_9 ;
wire un7_rnd_out_r_cry_8 ;
wire un7_rnd_out_r_cry_7 ;
wire un7_rnd_out_r_cry_6 ;
wire un7_rnd_out_r_cry_5 ;
wire un7_rnd_out_r_cry_4 ;
wire un7_rnd_out_r_cry_3 ;
wire un7_rnd_out_r_cry_2 ;
wire un7_rnd_out_r_cry_1 ;
wire un5_rnd_out_i_cry_11 ;
wire un5_rnd_out_i_cry_10 ;
wire un5_rnd_out_i_cry_9 ;
wire un5_rnd_out_i_cry_8 ;
wire un5_rnd_out_i_cry_7 ;
wire un5_rnd_out_i_cry_6 ;
wire un5_rnd_out_i_cry_5 ;
wire un5_rnd_out_i_cry_4 ;
wire un5_rnd_out_i_cry_3 ;
wire un5_rnd_out_i_cry_2 ;
wire un5_rnd_out_i_cry_1 ;
wire VCC ;
// instances
  LUT1 un5_rnd_out_i_axb_1_cZ(.I0(pre_out_i[8:8]),.O(un5_rnd_out_i_axb_1));
defparam un5_rnd_out_i_axb_1_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_2_cZ(.I0(pre_out_i[9:9]),.O(un5_rnd_out_i_axb_2));
defparam un5_rnd_out_i_axb_2_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_3_cZ(.I0(pre_out_i[10:10]),.O(un5_rnd_out_i_axb_3));
defparam un5_rnd_out_i_axb_3_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_4_cZ(.I0(pre_out_i[11:11]),.O(un5_rnd_out_i_axb_4));
defparam un5_rnd_out_i_axb_4_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_5_cZ(.I0(pre_out_i[12:12]),.O(un5_rnd_out_i_axb_5));
defparam un5_rnd_out_i_axb_5_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_6_cZ(.I0(pre_out_i[13:13]),.O(un5_rnd_out_i_axb_6));
defparam un5_rnd_out_i_axb_6_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_7_cZ(.I0(pre_out_i[14:14]),.O(un5_rnd_out_i_axb_7));
defparam un5_rnd_out_i_axb_7_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_8_cZ(.I0(pre_out_i[15:15]),.O(un5_rnd_out_i_axb_8));
defparam un5_rnd_out_i_axb_8_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_9_cZ(.I0(pre_out_i[16:16]),.O(un5_rnd_out_i_axb_9));
defparam un5_rnd_out_i_axb_9_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_10_cZ(.I0(pre_out_i[17:17]),.O(un5_rnd_out_i_axb_10));
defparam un5_rnd_out_i_axb_10_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_11_cZ(.I0(pre_out_i[18:18]),.O(un5_rnd_out_i_axb_11));
defparam un5_rnd_out_i_axb_11_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_1_cZ(.I0(pre_out_r[8:8]),.O(un7_rnd_out_r_axb_1));
defparam un7_rnd_out_r_axb_1_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_2_cZ(.I0(pre_out_r[9:9]),.O(un7_rnd_out_r_axb_2));
defparam un7_rnd_out_r_axb_2_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_3_cZ(.I0(pre_out_r[10:10]),.O(un7_rnd_out_r_axb_3));
defparam un7_rnd_out_r_axb_3_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_4_cZ(.I0(pre_out_r[11:11]),.O(un7_rnd_out_r_axb_4));
defparam un7_rnd_out_r_axb_4_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_5_cZ(.I0(pre_out_r[12:12]),.O(un7_rnd_out_r_axb_5));
defparam un7_rnd_out_r_axb_5_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_6_cZ(.I0(pre_out_r[13:13]),.O(un7_rnd_out_r_axb_6));
defparam un7_rnd_out_r_axb_6_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_7_cZ(.I0(pre_out_r[14:14]),.O(un7_rnd_out_r_axb_7));
defparam un7_rnd_out_r_axb_7_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_8_cZ(.I0(pre_out_r[15:15]),.O(un7_rnd_out_r_axb_8));
defparam un7_rnd_out_r_axb_8_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_9_cZ(.I0(pre_out_r[16:16]),.O(un7_rnd_out_r_axb_9));
defparam un7_rnd_out_r_axb_9_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_10_cZ(.I0(pre_out_r[17:17]),.O(un7_rnd_out_r_axb_10));
defparam un7_rnd_out_r_axb_10_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_11_cZ(.I0(pre_out_r[18:18]),.O(un7_rnd_out_r_axb_11));
defparam un7_rnd_out_r_axb_11_cZ.INIT=2'h2;
  LUT1 un7_rnd_out_r_axb_12_cZ(.I0(pre_out_r[19:19]),.O(un7_rnd_out_r_axb_12));
defparam un7_rnd_out_r_axb_12_cZ.INIT=2'h2;
  LUT1 un5_rnd_out_i_axb_12_cZ(.I0(pre_out_i[19:19]),.O(un5_rnd_out_i_axb_12));
defparam un5_rnd_out_i_axb_12_cZ.INIT=2'h2;
  LUT4 un4_rnd_sat_out_i_3_cZ(.I0(pre_out_i[20:20]),.I1(pre_out_i[21:21]),.I2(pre_out_i[22:22]),.I3(pre_out_i[19:19]),.O(un4_rnd_sat_out_i_3));
defparam un4_rnd_sat_out_i_3_cZ.INIT=16'h8000;
  LUT4 un5_rnd_sat_out_r_3_cZ(.I0(pre_out_r[20:20]),.I1(pre_out_r[21:21]),.I2(pre_out_r[22:22]),.I3(pre_out_r[19:19]),.O(un5_rnd_sat_out_r_3));
defparam un5_rnd_sat_out_r_3_cZ.INIT=16'h8000;
  LUT3 un1_pos_out_r(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.O(un1_pos_out_r_3));
defparam un1_pos_out_r.INIT=8'h08;
  LUT3 un1_pos_out_i(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.O(un1_pos_out_i_3));
defparam un1_pos_out_i.INIT=8'h02;
  LUT6_L desc270(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r_s_12),.LO(pos_out_r[11:11]));
defparam desc270.INIT=64'hE7E0E7E00000E0E0;
  LUT6_L desc271(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i_s_12),.LO(pos_out_i[11:11]));
defparam desc271.INIT=64'hBDB0BDB00000B0B0;
  LUT6_L desc272(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(un7_rnd_out_r[0:0]),.I4(PATTERNDETECT_7),.I5(un5_rnd_sat_out_r_3),.LO(pos_out_r_iv_i[0:0]));
defparam desc272.INIT=64'hFF18FF1F1F181F1F;
  LUT6_L desc273(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[1:1]),.LO(pos_out_r_iv_i[1:1]));
defparam desc273.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc274(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[2:2]),.LO(pos_out_r_iv_i[2:2]));
defparam desc274.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc275(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[3:3]),.LO(pos_out_r_iv_i[3:3]));
defparam desc275.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc276(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[4:4]),.LO(pos_out_r_iv_i[4:4]));
defparam desc276.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc277(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[5:5]),.LO(pos_out_r_iv_i[5:5]));
defparam desc277.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc278(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[6:6]),.LO(pos_out_r_iv_i[6:6]));
defparam desc278.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc279(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[7:7]),.LO(pos_out_r_iv_i[7:7]));
defparam desc279.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc280(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[8:8]),.LO(pos_out_r_iv_i[8:8]));
defparam desc280.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc281(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[9:9]),.LO(pos_out_r_iv_i[9:9]));
defparam desc281.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc282(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_7),.I4(un5_rnd_sat_out_r_3),.I5(un7_rnd_out_r[10:10]),.LO(pos_out_r_iv_i[10:10]));
defparam desc282.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc283(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(un5_rnd_out_i[0:0]),.I4(PATTERNDETECT_8),.I5(un4_rnd_sat_out_i_3),.LO(pos_out_i_iv_i[0:0]));
defparam desc283.INIT=64'hFF42FF4F4F424F4F;
  LUT6_L desc284(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[1:1]),.LO(pos_out_i_iv_i[1:1]));
defparam desc284.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc285(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[2:2]),.LO(pos_out_i_iv_i[2:2]));
defparam desc285.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc286(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[3:3]),.LO(pos_out_i_iv_i[3:3]));
defparam desc286.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc287(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[4:4]),.LO(pos_out_i_iv_i[4:4]));
defparam desc287.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc288(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[5:5]),.LO(pos_out_i_iv_i[5:5]));
defparam desc288.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc289(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[6:6]),.LO(pos_out_i_iv_i[6:6]));
defparam desc289.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc290(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[7:7]),.LO(pos_out_i_iv_i[7:7]));
defparam desc290.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc291(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[8:8]),.LO(pos_out_i_iv_i[8:8]));
defparam desc291.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc292(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[9:9]),.LO(pos_out_i_iv_i[9:9]));
defparam desc292.INIT=64'hFFFF4F4F424F424F;
  LUT6_L desc293(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_8),.I4(un4_rnd_sat_out_i_3),.I5(un5_rnd_out_i[10:10]),.LO(pos_out_i_iv_i[10:10]));
defparam desc293.INIT=64'hFFFF4F4F424F424F;
  XORCY un7_rnd_out_r_s_12_cZ(.LI(un7_rnd_out_r_axb_12),.CI(un7_rnd_out_r_cry_11),.O(un7_rnd_out_r_s_12));
  XORCY un7_rnd_out_r_s_11(.LI(un7_rnd_out_r_axb_11),.CI(un7_rnd_out_r_cry_10),.O(un7_rnd_out_r[10:10]));
  MUXCY_L un7_rnd_out_r_cry_11_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_10),.S(un7_rnd_out_r_axb_11),.LO(un7_rnd_out_r_cry_11));
  XORCY un7_rnd_out_r_s_10(.LI(un7_rnd_out_r_axb_10),.CI(un7_rnd_out_r_cry_9),.O(un7_rnd_out_r[9:9]));
  MUXCY_L un7_rnd_out_r_cry_10_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_9),.S(un7_rnd_out_r_axb_10),.LO(un7_rnd_out_r_cry_10));
  XORCY un7_rnd_out_r_s_9(.LI(un7_rnd_out_r_axb_9),.CI(un7_rnd_out_r_cry_8),.O(un7_rnd_out_r[8:8]));
  MUXCY_L un7_rnd_out_r_cry_9_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_8),.S(un7_rnd_out_r_axb_9),.LO(un7_rnd_out_r_cry_9));
  XORCY un7_rnd_out_r_s_8(.LI(un7_rnd_out_r_axb_8),.CI(un7_rnd_out_r_cry_7),.O(un7_rnd_out_r[7:7]));
  MUXCY_L un7_rnd_out_r_cry_8_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_7),.S(un7_rnd_out_r_axb_8),.LO(un7_rnd_out_r_cry_8));
  XORCY un7_rnd_out_r_s_7(.LI(un7_rnd_out_r_axb_7),.CI(un7_rnd_out_r_cry_6),.O(un7_rnd_out_r[6:6]));
  MUXCY_L un7_rnd_out_r_cry_7_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_6),.S(un7_rnd_out_r_axb_7),.LO(un7_rnd_out_r_cry_7));
  XORCY un7_rnd_out_r_s_6(.LI(un7_rnd_out_r_axb_6),.CI(un7_rnd_out_r_cry_5),.O(un7_rnd_out_r[5:5]));
  MUXCY_L un7_rnd_out_r_cry_6_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_5),.S(un7_rnd_out_r_axb_6),.LO(un7_rnd_out_r_cry_6));
  XORCY un7_rnd_out_r_s_5(.LI(un7_rnd_out_r_axb_5),.CI(un7_rnd_out_r_cry_4),.O(un7_rnd_out_r[4:4]));
  MUXCY_L un7_rnd_out_r_cry_5_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_4),.S(un7_rnd_out_r_axb_5),.LO(un7_rnd_out_r_cry_5));
  XORCY un7_rnd_out_r_s_4(.LI(un7_rnd_out_r_axb_4),.CI(un7_rnd_out_r_cry_3),.O(un7_rnd_out_r[3:3]));
  MUXCY_L un7_rnd_out_r_cry_4_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_3),.S(un7_rnd_out_r_axb_4),.LO(un7_rnd_out_r_cry_4));
  XORCY un7_rnd_out_r_s_3(.LI(un7_rnd_out_r_axb_3),.CI(un7_rnd_out_r_cry_2),.O(un7_rnd_out_r[2:2]));
  MUXCY_L un7_rnd_out_r_cry_3_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_2),.S(un7_rnd_out_r_axb_3),.LO(un7_rnd_out_r_cry_3));
  XORCY un7_rnd_out_r_s_2(.LI(un7_rnd_out_r_axb_2),.CI(un7_rnd_out_r_cry_1),.O(un7_rnd_out_r[1:1]));
  MUXCY_L un7_rnd_out_r_cry_2_cZ(.DI(GND),.CI(un7_rnd_out_r_cry_1),.S(un7_rnd_out_r_axb_2),.LO(un7_rnd_out_r_cry_2));
  XORCY un7_rnd_out_r_s_1(.LI(un7_rnd_out_r_axb_1),.CI(pre_out_r[7:7]),.O(un7_rnd_out_r[0:0]));
  MUXCY_L un7_rnd_out_r_cry_1_cZ(.DI(GND),.CI(pre_out_r[7:7]),.S(un7_rnd_out_r_axb_1),.LO(un7_rnd_out_r_cry_1));
  XORCY un5_rnd_out_i_s_12_cZ(.LI(un5_rnd_out_i_axb_12),.CI(un5_rnd_out_i_cry_11),.O(un5_rnd_out_i_s_12));
  XORCY un5_rnd_out_i_s_11(.LI(un5_rnd_out_i_axb_11),.CI(un5_rnd_out_i_cry_10),.O(un5_rnd_out_i[10:10]));
  MUXCY_L un5_rnd_out_i_cry_11_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_10),.S(un5_rnd_out_i_axb_11),.LO(un5_rnd_out_i_cry_11));
  XORCY un5_rnd_out_i_s_10(.LI(un5_rnd_out_i_axb_10),.CI(un5_rnd_out_i_cry_9),.O(un5_rnd_out_i[9:9]));
  MUXCY_L un5_rnd_out_i_cry_10_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_9),.S(un5_rnd_out_i_axb_10),.LO(un5_rnd_out_i_cry_10));
  XORCY un5_rnd_out_i_s_9(.LI(un5_rnd_out_i_axb_9),.CI(un5_rnd_out_i_cry_8),.O(un5_rnd_out_i[8:8]));
  MUXCY_L un5_rnd_out_i_cry_9_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_8),.S(un5_rnd_out_i_axb_9),.LO(un5_rnd_out_i_cry_9));
  XORCY un5_rnd_out_i_s_8(.LI(un5_rnd_out_i_axb_8),.CI(un5_rnd_out_i_cry_7),.O(un5_rnd_out_i[7:7]));
  MUXCY_L un5_rnd_out_i_cry_8_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_7),.S(un5_rnd_out_i_axb_8),.LO(un5_rnd_out_i_cry_8));
  XORCY un5_rnd_out_i_s_7(.LI(un5_rnd_out_i_axb_7),.CI(un5_rnd_out_i_cry_6),.O(un5_rnd_out_i[6:6]));
  MUXCY_L un5_rnd_out_i_cry_7_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_6),.S(un5_rnd_out_i_axb_7),.LO(un5_rnd_out_i_cry_7));
  XORCY un5_rnd_out_i_s_6(.LI(un5_rnd_out_i_axb_6),.CI(un5_rnd_out_i_cry_5),.O(un5_rnd_out_i[5:5]));
  MUXCY_L un5_rnd_out_i_cry_6_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_5),.S(un5_rnd_out_i_axb_6),.LO(un5_rnd_out_i_cry_6));
  XORCY un5_rnd_out_i_s_5(.LI(un5_rnd_out_i_axb_5),.CI(un5_rnd_out_i_cry_4),.O(un5_rnd_out_i[4:4]));
  MUXCY_L un5_rnd_out_i_cry_5_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_4),.S(un5_rnd_out_i_axb_5),.LO(un5_rnd_out_i_cry_5));
  XORCY un5_rnd_out_i_s_4(.LI(un5_rnd_out_i_axb_4),.CI(un5_rnd_out_i_cry_3),.O(un5_rnd_out_i[3:3]));
  MUXCY_L un5_rnd_out_i_cry_4_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_3),.S(un5_rnd_out_i_axb_4),.LO(un5_rnd_out_i_cry_4));
  XORCY un5_rnd_out_i_s_3(.LI(un5_rnd_out_i_axb_3),.CI(un5_rnd_out_i_cry_2),.O(un5_rnd_out_i[2:2]));
  MUXCY_L un5_rnd_out_i_cry_3_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_2),.S(un5_rnd_out_i_axb_3),.LO(un5_rnd_out_i_cry_3));
  XORCY un5_rnd_out_i_s_2(.LI(un5_rnd_out_i_axb_2),.CI(un5_rnd_out_i_cry_1),.O(un5_rnd_out_i[1:1]));
  MUXCY_L un5_rnd_out_i_cry_2_cZ(.DI(GND),.CI(un5_rnd_out_i_cry_1),.S(un5_rnd_out_i_axb_2),.LO(un5_rnd_out_i_cry_2));
  XORCY un5_rnd_out_i_s_1(.LI(un5_rnd_out_i_axb_1),.CI(pre_out_i[7:7]),.O(un5_rnd_out_i[0:0]));
  MUXCY_L un5_rnd_out_i_cry_1_cZ(.DI(GND),.CI(pre_out_i[7:7]),.S(un5_rnd_out_i_axb_1),.LO(un5_rnd_out_i_cry_1));
  FDR desc294(.Q(mult_out_r[0:0]),.D(pos_out_r_iv_i[0:0]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc295(.Q(mult_out_r[1:1]),.D(pos_out_r_iv_i[1:1]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc296(.Q(mult_out_r[2:2]),.D(pos_out_r_iv_i[2:2]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc297(.Q(mult_out_r[3:3]),.D(pos_out_r_iv_i[3:3]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc298(.Q(mult_out_r[4:4]),.D(pos_out_r_iv_i[4:4]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc299(.Q(mult_out_r[5:5]),.D(pos_out_r_iv_i[5:5]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc300(.Q(mult_out_r[6:6]),.D(pos_out_r_iv_i[6:6]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc301(.Q(mult_out_r[7:7]),.D(pos_out_r_iv_i[7:7]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc302(.Q(mult_out_r[8:8]),.D(pos_out_r_iv_i[8:8]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc303(.Q(mult_out_r[9:9]),.D(pos_out_r_iv_i[9:9]),.C(clk),.R(un1_pos_out_r_3));
  FDR desc304(.Q(mult_out_r[10:10]),.D(pos_out_r_iv_i[10:10]),.C(clk),.R(un1_pos_out_r_3));
  FDS desc305(.Q(mult_out_r[11:11]),.D(pos_out_r[11:11]),.C(clk),.S(un1_pos_out_r_3));
  FDR desc306(.Q(mult_out_i[0:0]),.D(pos_out_i_iv_i[0:0]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc307(.Q(mult_out_i[1:1]),.D(pos_out_i_iv_i[1:1]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc308(.Q(mult_out_i[2:2]),.D(pos_out_i_iv_i[2:2]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc309(.Q(mult_out_i[3:3]),.D(pos_out_i_iv_i[3:3]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc310(.Q(mult_out_i[4:4]),.D(pos_out_i_iv_i[4:4]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc311(.Q(mult_out_i[5:5]),.D(pos_out_i_iv_i[5:5]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc312(.Q(mult_out_i[6:6]),.D(pos_out_i_iv_i[6:6]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc313(.Q(mult_out_i[7:7]),.D(pos_out_i_iv_i[7:7]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc314(.Q(mult_out_i[8:8]),.D(pos_out_i_iv_i[8:8]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc315(.Q(mult_out_i[9:9]),.D(pos_out_i_iv_i[9:9]),.C(clk),.R(un1_pos_out_i_3));
  FDR desc316(.Q(mult_out_i[10:10]),.D(pos_out_i_iv_i[10:10]),.C(clk),.R(un1_pos_out_i_3));
  FDS desc317(.Q(mult_out_i[11:11]),.D(pos_out_i[11:11]),.C(clk),.S(un1_pos_out_i_3));
  mult_pipe_inj mult1(.mult1_out(mult1_out[23:23]),.in_a_r_reg(in_a_r_reg[11:0]),.in_b_r_reg(in_b_r_reg[11:0]),.clk(clk));
  mult_pipe_1_inj mult2(.mult2_out_23(mult2_out[23:23]),.mult2_out_0(mult2_out_0[23:0]),.P_uc_34_0(P_uc_34_0[47:24]),.in_a_i_reg(in_a_i_reg[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk));
  mult_pipe_2_inj mult3(.mult3_out_23(mult3_out[23:23]),.mult3_out_0(mult3_out_0[23:0]),.P_uc_35_0(P_uc_35_0[47:24]),.in_a_r_reg(in_a_r_reg[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk));
  mult_pipe_3_inj mult4(.mult4_out(mult4_out[23:23]),.in_a_i_reg(in_a_i_reg[11:0]),.in_b_r_reg(in_b_r_reg[11:0]),.clk(clk));
  add_subZ1_inj add(.pre_out_r(pre_out_r[23:7]),.in_a_r_reg(in_a_r_reg[11:0]),.in_b_r_reg(in_b_r_reg[11:0]),.mult2_out_0(mult2_out_0[23:0]),.P_uc_34_0(P_uc_34_0[47:24]),.PATTERNDETECT_7(PATTERNDETECT_7),.clk(clk));
  add_subZ2_inj sub(.pre_out_i(pre_out_i[23:7]),.in_a_i_reg(in_a_i_reg[11:0]),.in_b_r_reg(in_b_r_reg[11:0]),.mult3_out_0(mult3_out_0[23:0]),.P_uc_35_0(P_uc_35_0[47:24]),.PATTERNDETECT_8(PATTERNDETECT_8),.clk(clk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module desc481_inj (out_i_vec_mult_2,out_r_vec_mult_2,out_inner_prod_r,vec_out_r_AQ_2,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,vec_out_i_AQ_2,out_inner_prod_i,in_b_i_reg,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output [11:0] out_i_vec_mult_2 ;
output [11:0] out_r_vec_mult_2 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_2 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input [11:0] vec_out_i_AQ_2 ;
input [11:0] out_inner_prod_i ;
input [11:0] in_b_i_reg ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [23:7] pre_out_r ;
wire [23:7] pre_out_i ;
wire [23:23] mult2_out ;
wire [23:23] mult1_out ;
wire [23:23] mult3_out ;
wire [23:23] mult4_out ;
wire [11:11] pos_out_r ;
wire [11:11] pos_out_i ;
wire [10:0] un1_rnd_out_i ;
wire [10:0] pos_out_i_iv_i ;
wire [10:0] un2_rnd_out_r ;
wire [10:0] pos_out_r_iv_i ;
wire [23:0] mult1_out_0 ;
wire [47:24] P_uc_24_0 ;
wire [23:0] mult4_out_0 ;
wire [47:24] P_uc_27_0 ;
wire un2_rnd_out_r_axb_1 ;
wire un2_rnd_out_r_axb_2 ;
wire un2_rnd_out_r_axb_3 ;
wire un2_rnd_out_r_axb_4 ;
wire un2_rnd_out_r_axb_5 ;
wire un2_rnd_out_r_axb_6 ;
wire un2_rnd_out_r_axb_7 ;
wire un2_rnd_out_r_axb_8 ;
wire un2_rnd_out_r_axb_9 ;
wire un2_rnd_out_r_axb_10 ;
wire un2_rnd_out_r_axb_11 ;
wire un1_rnd_out_i_axb_1 ;
wire un1_rnd_out_i_axb_2 ;
wire un1_rnd_out_i_axb_3 ;
wire un1_rnd_out_i_axb_4 ;
wire un1_rnd_out_i_axb_5 ;
wire un1_rnd_out_i_axb_6 ;
wire un1_rnd_out_i_axb_7 ;
wire un1_rnd_out_i_axb_8 ;
wire un1_rnd_out_i_axb_9 ;
wire un1_rnd_out_i_axb_10 ;
wire un1_rnd_out_i_axb_11 ;
wire un1_rnd_out_i_axb_12 ;
wire un2_rnd_out_r_axb_12 ;
wire un5_rnd_sat_out_r_3 ;
wire un4_rnd_sat_out_i_3 ;
wire un1_pos_out_r ;
wire un1_pos_out_i ;
wire PATTERNDETECT_4 ;
wire un2_rnd_out_r_s_12 ;
wire PATTERNDETECT_3 ;
wire un1_rnd_out_i_s_12 ;
wire un1_rnd_out_i_cry_11 ;
wire un1_rnd_out_i_cry_10 ;
wire GND ;
wire un1_rnd_out_i_cry_9 ;
wire un1_rnd_out_i_cry_8 ;
wire un1_rnd_out_i_cry_7 ;
wire un1_rnd_out_i_cry_6 ;
wire un1_rnd_out_i_cry_5 ;
wire un1_rnd_out_i_cry_4 ;
wire un1_rnd_out_i_cry_3 ;
wire un1_rnd_out_i_cry_2 ;
wire un1_rnd_out_i_cry_1 ;
wire un2_rnd_out_r_cry_11 ;
wire un2_rnd_out_r_cry_10 ;
wire un2_rnd_out_r_cry_9 ;
wire un2_rnd_out_r_cry_8 ;
wire un2_rnd_out_r_cry_7 ;
wire un2_rnd_out_r_cry_6 ;
wire un2_rnd_out_r_cry_5 ;
wire un2_rnd_out_r_cry_4 ;
wire un2_rnd_out_r_cry_3 ;
wire un2_rnd_out_r_cry_2 ;
wire un2_rnd_out_r_cry_1 ;
wire VCC ;
// instances
  LUT1 un2_rnd_out_r_axb_1_cZ(.I0(pre_out_r[8:8]),.O(un2_rnd_out_r_axb_1));
defparam un2_rnd_out_r_axb_1_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_2_cZ(.I0(pre_out_r[9:9]),.O(un2_rnd_out_r_axb_2));
defparam un2_rnd_out_r_axb_2_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_3_cZ(.I0(pre_out_r[10:10]),.O(un2_rnd_out_r_axb_3));
defparam un2_rnd_out_r_axb_3_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_4_cZ(.I0(pre_out_r[11:11]),.O(un2_rnd_out_r_axb_4));
defparam un2_rnd_out_r_axb_4_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_5_cZ(.I0(pre_out_r[12:12]),.O(un2_rnd_out_r_axb_5));
defparam un2_rnd_out_r_axb_5_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_6_cZ(.I0(pre_out_r[13:13]),.O(un2_rnd_out_r_axb_6));
defparam un2_rnd_out_r_axb_6_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_7_cZ(.I0(pre_out_r[14:14]),.O(un2_rnd_out_r_axb_7));
defparam un2_rnd_out_r_axb_7_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_8_cZ(.I0(pre_out_r[15:15]),.O(un2_rnd_out_r_axb_8));
defparam un2_rnd_out_r_axb_8_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_9_cZ(.I0(pre_out_r[16:16]),.O(un2_rnd_out_r_axb_9));
defparam un2_rnd_out_r_axb_9_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_10_cZ(.I0(pre_out_r[17:17]),.O(un2_rnd_out_r_axb_10));
defparam un2_rnd_out_r_axb_10_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_11_cZ(.I0(pre_out_r[18:18]),.O(un2_rnd_out_r_axb_11));
defparam un2_rnd_out_r_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_1_cZ(.I0(pre_out_i[8:8]),.O(un1_rnd_out_i_axb_1));
defparam un1_rnd_out_i_axb_1_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_2_cZ(.I0(pre_out_i[9:9]),.O(un1_rnd_out_i_axb_2));
defparam un1_rnd_out_i_axb_2_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_3_cZ(.I0(pre_out_i[10:10]),.O(un1_rnd_out_i_axb_3));
defparam un1_rnd_out_i_axb_3_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_4_cZ(.I0(pre_out_i[11:11]),.O(un1_rnd_out_i_axb_4));
defparam un1_rnd_out_i_axb_4_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_5_cZ(.I0(pre_out_i[12:12]),.O(un1_rnd_out_i_axb_5));
defparam un1_rnd_out_i_axb_5_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_6_cZ(.I0(pre_out_i[13:13]),.O(un1_rnd_out_i_axb_6));
defparam un1_rnd_out_i_axb_6_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_7_cZ(.I0(pre_out_i[14:14]),.O(un1_rnd_out_i_axb_7));
defparam un1_rnd_out_i_axb_7_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_8_cZ(.I0(pre_out_i[15:15]),.O(un1_rnd_out_i_axb_8));
defparam un1_rnd_out_i_axb_8_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_9_cZ(.I0(pre_out_i[16:16]),.O(un1_rnd_out_i_axb_9));
defparam un1_rnd_out_i_axb_9_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_10_cZ(.I0(pre_out_i[17:17]),.O(un1_rnd_out_i_axb_10));
defparam un1_rnd_out_i_axb_10_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_11_cZ(.I0(pre_out_i[18:18]),.O(un1_rnd_out_i_axb_11));
defparam un1_rnd_out_i_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_12_cZ(.I0(pre_out_i[19:19]),.O(un1_rnd_out_i_axb_12));
defparam un1_rnd_out_i_axb_12_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_12_cZ(.I0(pre_out_r[19:19]),.O(un2_rnd_out_r_axb_12));
defparam un2_rnd_out_r_axb_12_cZ.INIT=2'h2;
  LUT4 un5_rnd_sat_out_r_3_cZ(.I0(pre_out_r[20:20]),.I1(pre_out_r[21:21]),.I2(pre_out_r[22:22]),.I3(pre_out_r[19:19]),.O(un5_rnd_sat_out_r_3));
defparam un5_rnd_sat_out_r_3_cZ.INIT=16'h8000;
  LUT4 un4_rnd_sat_out_i_3_cZ(.I0(pre_out_i[20:20]),.I1(pre_out_i[21:21]),.I2(pre_out_i[22:22]),.I3(pre_out_i[19:19]),.O(un4_rnd_sat_out_i_3));
defparam un4_rnd_sat_out_i_3_cZ.INIT=16'h8000;
  LUT3 un1_pos_out_r_cZ(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.O(un1_pos_out_r));
defparam un1_pos_out_r_cZ.INIT=8'h04;
  LUT3 un1_pos_out_i_cZ(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.O(un1_pos_out_i));
defparam un1_pos_out_i_cZ.INIT=8'h08;
  LUT6_L desc482(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r_s_12),.LO(pos_out_r[11:11]));
defparam desc482.INIT=64'hDBD0DBD00000D0D0;
  LUT6_L desc483(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i_s_12),.LO(pos_out_i[11:11]));
defparam desc483.INIT=64'hE7E0E7E00000E0E0;
  LUT6_L desc484(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[10:10]),.LO(pos_out_i_iv_i[10:10]));
defparam desc484.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc485(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[9:9]),.LO(pos_out_i_iv_i[9:9]));
defparam desc485.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc486(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[8:8]),.LO(pos_out_i_iv_i[8:8]));
defparam desc486.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc487(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[7:7]),.LO(pos_out_i_iv_i[7:7]));
defparam desc487.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc488(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[6:6]),.LO(pos_out_i_iv_i[6:6]));
defparam desc488.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc489(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[5:5]),.LO(pos_out_i_iv_i[5:5]));
defparam desc489.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc490(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[4:4]),.LO(pos_out_i_iv_i[4:4]));
defparam desc490.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc491(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[3:3]),.LO(pos_out_i_iv_i[3:3]));
defparam desc491.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc492(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[2:2]),.LO(pos_out_i_iv_i[2:2]));
defparam desc492.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc493(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_3),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[1:1]),.LO(pos_out_i_iv_i[1:1]));
defparam desc493.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc494(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(un1_rnd_out_i[0:0]),.I4(PATTERNDETECT_3),.I5(un4_rnd_sat_out_i_3),.LO(pos_out_i_iv_i[0:0]));
defparam desc494.INIT=64'hFF18FF1F1F181F1F;
  LUT6_L desc495(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[10:10]),.LO(pos_out_r_iv_i[10:10]));
defparam desc495.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc496(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[9:9]),.LO(pos_out_r_iv_i[9:9]));
defparam desc496.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc497(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[8:8]),.LO(pos_out_r_iv_i[8:8]));
defparam desc497.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc498(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[7:7]),.LO(pos_out_r_iv_i[7:7]));
defparam desc498.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc499(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[6:6]),.LO(pos_out_r_iv_i[6:6]));
defparam desc499.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc500(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[5:5]),.LO(pos_out_r_iv_i[5:5]));
defparam desc500.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc501(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[4:4]),.LO(pos_out_r_iv_i[4:4]));
defparam desc501.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc502(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[3:3]),.LO(pos_out_r_iv_i[3:3]));
defparam desc502.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc503(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[2:2]),.LO(pos_out_r_iv_i[2:2]));
defparam desc503.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc504(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_4),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[1:1]),.LO(pos_out_r_iv_i[1:1]));
defparam desc504.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc505(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(un2_rnd_out_r[0:0]),.I4(PATTERNDETECT_4),.I5(un5_rnd_sat_out_r_3),.LO(pos_out_r_iv_i[0:0]));
defparam desc505.INIT=64'hFF24FF2F2F242F2F;
  XORCY un1_rnd_out_i_s_12_cZ(.LI(un1_rnd_out_i_axb_12),.CI(un1_rnd_out_i_cry_11),.O(un1_rnd_out_i_s_12));
  XORCY un1_rnd_out_i_s_11(.LI(un1_rnd_out_i_axb_11),.CI(un1_rnd_out_i_cry_10),.O(un1_rnd_out_i[10:10]));
  MUXCY_L un1_rnd_out_i_cry_11_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_10),.S(un1_rnd_out_i_axb_11),.LO(un1_rnd_out_i_cry_11));
  XORCY un1_rnd_out_i_s_10(.LI(un1_rnd_out_i_axb_10),.CI(un1_rnd_out_i_cry_9),.O(un1_rnd_out_i[9:9]));
  MUXCY_L un1_rnd_out_i_cry_10_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_9),.S(un1_rnd_out_i_axb_10),.LO(un1_rnd_out_i_cry_10));
  XORCY un1_rnd_out_i_s_9(.LI(un1_rnd_out_i_axb_9),.CI(un1_rnd_out_i_cry_8),.O(un1_rnd_out_i[8:8]));
  MUXCY_L un1_rnd_out_i_cry_9_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_8),.S(un1_rnd_out_i_axb_9),.LO(un1_rnd_out_i_cry_9));
  XORCY un1_rnd_out_i_s_8(.LI(un1_rnd_out_i_axb_8),.CI(un1_rnd_out_i_cry_7),.O(un1_rnd_out_i[7:7]));
  MUXCY_L un1_rnd_out_i_cry_8_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_7),.S(un1_rnd_out_i_axb_8),.LO(un1_rnd_out_i_cry_8));
  XORCY un1_rnd_out_i_s_7(.LI(un1_rnd_out_i_axb_7),.CI(un1_rnd_out_i_cry_6),.O(un1_rnd_out_i[6:6]));
  MUXCY_L un1_rnd_out_i_cry_7_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_6),.S(un1_rnd_out_i_axb_7),.LO(un1_rnd_out_i_cry_7));
  XORCY un1_rnd_out_i_s_6(.LI(un1_rnd_out_i_axb_6),.CI(un1_rnd_out_i_cry_5),.O(un1_rnd_out_i[5:5]));
  MUXCY_L un1_rnd_out_i_cry_6_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_5),.S(un1_rnd_out_i_axb_6),.LO(un1_rnd_out_i_cry_6));
  XORCY un1_rnd_out_i_s_5(.LI(un1_rnd_out_i_axb_5),.CI(un1_rnd_out_i_cry_4),.O(un1_rnd_out_i[4:4]));
  MUXCY_L un1_rnd_out_i_cry_5_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_4),.S(un1_rnd_out_i_axb_5),.LO(un1_rnd_out_i_cry_5));
  XORCY un1_rnd_out_i_s_4(.LI(un1_rnd_out_i_axb_4),.CI(un1_rnd_out_i_cry_3),.O(un1_rnd_out_i[3:3]));
  MUXCY_L un1_rnd_out_i_cry_4_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_3),.S(un1_rnd_out_i_axb_4),.LO(un1_rnd_out_i_cry_4));
  XORCY un1_rnd_out_i_s_3(.LI(un1_rnd_out_i_axb_3),.CI(un1_rnd_out_i_cry_2),.O(un1_rnd_out_i[2:2]));
  MUXCY_L un1_rnd_out_i_cry_3_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_2),.S(un1_rnd_out_i_axb_3),.LO(un1_rnd_out_i_cry_3));
  XORCY un1_rnd_out_i_s_2(.LI(un1_rnd_out_i_axb_2),.CI(un1_rnd_out_i_cry_1),.O(un1_rnd_out_i[1:1]));
  MUXCY_L un1_rnd_out_i_cry_2_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_1),.S(un1_rnd_out_i_axb_2),.LO(un1_rnd_out_i_cry_2));
  XORCY un1_rnd_out_i_s_1(.LI(un1_rnd_out_i_axb_1),.CI(pre_out_i[7:7]),.O(un1_rnd_out_i[0:0]));
  MUXCY_L un1_rnd_out_i_cry_1_cZ(.DI(GND),.CI(pre_out_i[7:7]),.S(un1_rnd_out_i_axb_1),.LO(un1_rnd_out_i_cry_1));
  XORCY un2_rnd_out_r_s_12_cZ(.LI(un2_rnd_out_r_axb_12),.CI(un2_rnd_out_r_cry_11),.O(un2_rnd_out_r_s_12));
  XORCY un2_rnd_out_r_s_11(.LI(un2_rnd_out_r_axb_11),.CI(un2_rnd_out_r_cry_10),.O(un2_rnd_out_r[10:10]));
  MUXCY_L un2_rnd_out_r_cry_11_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_10),.S(un2_rnd_out_r_axb_11),.LO(un2_rnd_out_r_cry_11));
  XORCY un2_rnd_out_r_s_10(.LI(un2_rnd_out_r_axb_10),.CI(un2_rnd_out_r_cry_9),.O(un2_rnd_out_r[9:9]));
  MUXCY_L un2_rnd_out_r_cry_10_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_9),.S(un2_rnd_out_r_axb_10),.LO(un2_rnd_out_r_cry_10));
  XORCY un2_rnd_out_r_s_9(.LI(un2_rnd_out_r_axb_9),.CI(un2_rnd_out_r_cry_8),.O(un2_rnd_out_r[8:8]));
  MUXCY_L un2_rnd_out_r_cry_9_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_8),.S(un2_rnd_out_r_axb_9),.LO(un2_rnd_out_r_cry_9));
  XORCY un2_rnd_out_r_s_8(.LI(un2_rnd_out_r_axb_8),.CI(un2_rnd_out_r_cry_7),.O(un2_rnd_out_r[7:7]));
  MUXCY_L un2_rnd_out_r_cry_8_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_7),.S(un2_rnd_out_r_axb_8),.LO(un2_rnd_out_r_cry_8));
  XORCY un2_rnd_out_r_s_7(.LI(un2_rnd_out_r_axb_7),.CI(un2_rnd_out_r_cry_6),.O(un2_rnd_out_r[6:6]));
  MUXCY_L un2_rnd_out_r_cry_7_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_6),.S(un2_rnd_out_r_axb_7),.LO(un2_rnd_out_r_cry_7));
  XORCY un2_rnd_out_r_s_6(.LI(un2_rnd_out_r_axb_6),.CI(un2_rnd_out_r_cry_5),.O(un2_rnd_out_r[5:5]));
  MUXCY_L un2_rnd_out_r_cry_6_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_5),.S(un2_rnd_out_r_axb_6),.LO(un2_rnd_out_r_cry_6));
  XORCY un2_rnd_out_r_s_5(.LI(un2_rnd_out_r_axb_5),.CI(un2_rnd_out_r_cry_4),.O(un2_rnd_out_r[4:4]));
  MUXCY_L un2_rnd_out_r_cry_5_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_4),.S(un2_rnd_out_r_axb_5),.LO(un2_rnd_out_r_cry_5));
  XORCY un2_rnd_out_r_s_4(.LI(un2_rnd_out_r_axb_4),.CI(un2_rnd_out_r_cry_3),.O(un2_rnd_out_r[3:3]));
  MUXCY_L un2_rnd_out_r_cry_4_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_3),.S(un2_rnd_out_r_axb_4),.LO(un2_rnd_out_r_cry_4));
  XORCY un2_rnd_out_r_s_3(.LI(un2_rnd_out_r_axb_3),.CI(un2_rnd_out_r_cry_2),.O(un2_rnd_out_r[2:2]));
  MUXCY_L un2_rnd_out_r_cry_3_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_2),.S(un2_rnd_out_r_axb_3),.LO(un2_rnd_out_r_cry_3));
  XORCY un2_rnd_out_r_s_2(.LI(un2_rnd_out_r_axb_2),.CI(un2_rnd_out_r_cry_1),.O(un2_rnd_out_r[1:1]));
  MUXCY_L un2_rnd_out_r_cry_2_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_1),.S(un2_rnd_out_r_axb_2),.LO(un2_rnd_out_r_cry_2));
  XORCY un2_rnd_out_r_s_1(.LI(un2_rnd_out_r_axb_1),.CI(pre_out_r[7:7]),.O(un2_rnd_out_r[0:0]));
  MUXCY_L un2_rnd_out_r_cry_1_cZ(.DI(GND),.CI(pre_out_r[7:7]),.S(un2_rnd_out_r_axb_1),.LO(un2_rnd_out_r_cry_1));
  FDS desc506(.Q(out_i_vec_mult_2[11:11]),.D(pos_out_i[11:11]),.C(clk),.S(un1_pos_out_i));
  FDR desc507(.Q(out_i_vec_mult_2[10:10]),.D(pos_out_i_iv_i[10:10]),.C(clk),.R(un1_pos_out_i));
  FDR desc508(.Q(out_i_vec_mult_2[9:9]),.D(pos_out_i_iv_i[9:9]),.C(clk),.R(un1_pos_out_i));
  FDR desc509(.Q(out_i_vec_mult_2[8:8]),.D(pos_out_i_iv_i[8:8]),.C(clk),.R(un1_pos_out_i));
  FDR desc510(.Q(out_i_vec_mult_2[7:7]),.D(pos_out_i_iv_i[7:7]),.C(clk),.R(un1_pos_out_i));
  FDR desc511(.Q(out_i_vec_mult_2[6:6]),.D(pos_out_i_iv_i[6:6]),.C(clk),.R(un1_pos_out_i));
  FDR desc512(.Q(out_i_vec_mult_2[5:5]),.D(pos_out_i_iv_i[5:5]),.C(clk),.R(un1_pos_out_i));
  FDR desc513(.Q(out_i_vec_mult_2[4:4]),.D(pos_out_i_iv_i[4:4]),.C(clk),.R(un1_pos_out_i));
  FDR desc514(.Q(out_i_vec_mult_2[3:3]),.D(pos_out_i_iv_i[3:3]),.C(clk),.R(un1_pos_out_i));
  FDR desc515(.Q(out_i_vec_mult_2[2:2]),.D(pos_out_i_iv_i[2:2]),.C(clk),.R(un1_pos_out_i));
  FDR desc516(.Q(out_i_vec_mult_2[1:1]),.D(pos_out_i_iv_i[1:1]),.C(clk),.R(un1_pos_out_i));
  FDR desc517(.Q(out_i_vec_mult_2[0:0]),.D(pos_out_i_iv_i[0:0]),.C(clk),.R(un1_pos_out_i));
  FDS desc518(.Q(out_r_vec_mult_2[11:11]),.D(pos_out_r[11:11]),.C(clk),.S(un1_pos_out_r));
  FDR desc519(.Q(out_r_vec_mult_2[10:10]),.D(pos_out_r_iv_i[10:10]),.C(clk),.R(un1_pos_out_r));
  FDR desc520(.Q(out_r_vec_mult_2[9:9]),.D(pos_out_r_iv_i[9:9]),.C(clk),.R(un1_pos_out_r));
  FDR desc521(.Q(out_r_vec_mult_2[8:8]),.D(pos_out_r_iv_i[8:8]),.C(clk),.R(un1_pos_out_r));
  FDR desc522(.Q(out_r_vec_mult_2[7:7]),.D(pos_out_r_iv_i[7:7]),.C(clk),.R(un1_pos_out_r));
  FDR desc523(.Q(out_r_vec_mult_2[6:6]),.D(pos_out_r_iv_i[6:6]),.C(clk),.R(un1_pos_out_r));
  FDR desc524(.Q(out_r_vec_mult_2[5:5]),.D(pos_out_r_iv_i[5:5]),.C(clk),.R(un1_pos_out_r));
  FDR desc525(.Q(out_r_vec_mult_2[4:4]),.D(pos_out_r_iv_i[4:4]),.C(clk),.R(un1_pos_out_r));
  FDR desc526(.Q(out_r_vec_mult_2[3:3]),.D(pos_out_r_iv_i[3:3]),.C(clk),.R(un1_pos_out_r));
  FDR desc527(.Q(out_r_vec_mult_2[2:2]),.D(pos_out_r_iv_i[2:2]),.C(clk),.R(un1_pos_out_r));
  FDR desc528(.Q(out_r_vec_mult_2[1:1]),.D(pos_out_r_iv_i[1:1]),.C(clk),.R(un1_pos_out_r));
  FDR desc529(.Q(out_r_vec_mult_2[0:0]),.D(pos_out_r_iv_i[0:0]),.C(clk),.R(un1_pos_out_r));
  mult_pipe_4_inj mult1(.mult1_out_23(mult1_out[23:23]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_24_0(P_uc_24_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  mult_pipe_5_inj mult2(.mult2_out_23(mult2_out[23:23]),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_6_inj mult3(.mult3_out_23(mult3_out[23:23]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_7_inj mult4(.mult4_out_23(mult4_out[23:23]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_27_0(P_uc_27_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  add_subZ2_1_inj sub(.pre_out_r(pre_out_r[23:7]),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_24_0(P_uc_24_0[47:24]),.PATTERNDETECT_4(PATTERNDETECT_4),.clk(clk));
  add_subZ1_1_inj add(.pre_out_i(pre_out_i[23:7]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_27_0(P_uc_27_0[47:24]),.PATTERNDETECT_3(PATTERNDETECT_3),.clk(clk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module desc536_inj (out_i_vec_mult_1,out_r_vec_mult_1,out_inner_prod_r,vec_out_r_AQ_1,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,vec_out_i_AQ_1,out_inner_prod_i,in_b_i_reg,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output [11:0] out_i_vec_mult_1 ;
output [11:0] out_r_vec_mult_1 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_1 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input [11:0] vec_out_i_AQ_1 ;
input [11:0] out_inner_prod_i ;
input [11:0] in_b_i_reg ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [23:7] pre_out_r ;
wire [23:7] pre_out_i ;
wire [23:23] mult2_out ;
wire [23:23] mult1_out ;
wire [23:23] mult3_out ;
wire [23:23] mult4_out ;
wire [11:11] pos_out_r ;
wire [11:11] pos_out_i ;
wire [10:0] un1_rnd_out_i ;
wire [10:0] pos_out_i_iv_i ;
wire [10:0] un2_rnd_out_r ;
wire [10:0] pos_out_r_iv_i ;
wire [23:0] mult1_out_0 ;
wire [47:24] P_uc_20_0 ;
wire [23:0] mult4_out_0 ;
wire [47:24] P_uc_23_0 ;
wire un2_rnd_out_r_axb_1 ;
wire un2_rnd_out_r_axb_2 ;
wire un2_rnd_out_r_axb_3 ;
wire un2_rnd_out_r_axb_4 ;
wire un2_rnd_out_r_axb_5 ;
wire un2_rnd_out_r_axb_6 ;
wire un2_rnd_out_r_axb_7 ;
wire un2_rnd_out_r_axb_8 ;
wire un2_rnd_out_r_axb_9 ;
wire un2_rnd_out_r_axb_10 ;
wire un2_rnd_out_r_axb_11 ;
wire un1_rnd_out_i_axb_1 ;
wire un1_rnd_out_i_axb_2 ;
wire un1_rnd_out_i_axb_3 ;
wire un1_rnd_out_i_axb_4 ;
wire un1_rnd_out_i_axb_5 ;
wire un1_rnd_out_i_axb_6 ;
wire un1_rnd_out_i_axb_7 ;
wire un1_rnd_out_i_axb_8 ;
wire un1_rnd_out_i_axb_9 ;
wire un1_rnd_out_i_axb_10 ;
wire un1_rnd_out_i_axb_11 ;
wire un1_rnd_out_i_axb_12 ;
wire un2_rnd_out_r_axb_12 ;
wire un4_rnd_sat_out_i_3 ;
wire un5_rnd_sat_out_r_3 ;
wire un1_pos_out_r_0 ;
wire un1_pos_out_i_0 ;
wire PATTERNDETECT_2 ;
wire un2_rnd_out_r_s_12_2 ;
wire PATTERNDETECT_1 ;
wire un1_rnd_out_i_s_12_2 ;
wire un1_rnd_out_i_cry_11 ;
wire un1_rnd_out_i_cry_10 ;
wire GND ;
wire un1_rnd_out_i_cry_9 ;
wire un1_rnd_out_i_cry_8 ;
wire un1_rnd_out_i_cry_7 ;
wire un1_rnd_out_i_cry_6 ;
wire un1_rnd_out_i_cry_5 ;
wire un1_rnd_out_i_cry_4 ;
wire un1_rnd_out_i_cry_3 ;
wire un1_rnd_out_i_cry_2 ;
wire un1_rnd_out_i_cry_1 ;
wire un2_rnd_out_r_cry_11 ;
wire un2_rnd_out_r_cry_10 ;
wire un2_rnd_out_r_cry_9 ;
wire un2_rnd_out_r_cry_8 ;
wire un2_rnd_out_r_cry_7 ;
wire un2_rnd_out_r_cry_6 ;
wire un2_rnd_out_r_cry_5 ;
wire un2_rnd_out_r_cry_4 ;
wire un2_rnd_out_r_cry_3 ;
wire un2_rnd_out_r_cry_2 ;
wire un2_rnd_out_r_cry_1 ;
wire VCC ;
// instances
  LUT1 un2_rnd_out_r_axb_1_cZ(.I0(pre_out_r[8:8]),.O(un2_rnd_out_r_axb_1));
defparam un2_rnd_out_r_axb_1_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_2_cZ(.I0(pre_out_r[9:9]),.O(un2_rnd_out_r_axb_2));
defparam un2_rnd_out_r_axb_2_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_3_cZ(.I0(pre_out_r[10:10]),.O(un2_rnd_out_r_axb_3));
defparam un2_rnd_out_r_axb_3_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_4_cZ(.I0(pre_out_r[11:11]),.O(un2_rnd_out_r_axb_4));
defparam un2_rnd_out_r_axb_4_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_5_cZ(.I0(pre_out_r[12:12]),.O(un2_rnd_out_r_axb_5));
defparam un2_rnd_out_r_axb_5_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_6_cZ(.I0(pre_out_r[13:13]),.O(un2_rnd_out_r_axb_6));
defparam un2_rnd_out_r_axb_6_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_7_cZ(.I0(pre_out_r[14:14]),.O(un2_rnd_out_r_axb_7));
defparam un2_rnd_out_r_axb_7_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_8_cZ(.I0(pre_out_r[15:15]),.O(un2_rnd_out_r_axb_8));
defparam un2_rnd_out_r_axb_8_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_9_cZ(.I0(pre_out_r[16:16]),.O(un2_rnd_out_r_axb_9));
defparam un2_rnd_out_r_axb_9_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_10_cZ(.I0(pre_out_r[17:17]),.O(un2_rnd_out_r_axb_10));
defparam un2_rnd_out_r_axb_10_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_11_cZ(.I0(pre_out_r[18:18]),.O(un2_rnd_out_r_axb_11));
defparam un2_rnd_out_r_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_1_cZ(.I0(pre_out_i[8:8]),.O(un1_rnd_out_i_axb_1));
defparam un1_rnd_out_i_axb_1_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_2_cZ(.I0(pre_out_i[9:9]),.O(un1_rnd_out_i_axb_2));
defparam un1_rnd_out_i_axb_2_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_3_cZ(.I0(pre_out_i[10:10]),.O(un1_rnd_out_i_axb_3));
defparam un1_rnd_out_i_axb_3_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_4_cZ(.I0(pre_out_i[11:11]),.O(un1_rnd_out_i_axb_4));
defparam un1_rnd_out_i_axb_4_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_5_cZ(.I0(pre_out_i[12:12]),.O(un1_rnd_out_i_axb_5));
defparam un1_rnd_out_i_axb_5_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_6_cZ(.I0(pre_out_i[13:13]),.O(un1_rnd_out_i_axb_6));
defparam un1_rnd_out_i_axb_6_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_7_cZ(.I0(pre_out_i[14:14]),.O(un1_rnd_out_i_axb_7));
defparam un1_rnd_out_i_axb_7_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_8_cZ(.I0(pre_out_i[15:15]),.O(un1_rnd_out_i_axb_8));
defparam un1_rnd_out_i_axb_8_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_9_cZ(.I0(pre_out_i[16:16]),.O(un1_rnd_out_i_axb_9));
defparam un1_rnd_out_i_axb_9_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_10_cZ(.I0(pre_out_i[17:17]),.O(un1_rnd_out_i_axb_10));
defparam un1_rnd_out_i_axb_10_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_11_cZ(.I0(pre_out_i[18:18]),.O(un1_rnd_out_i_axb_11));
defparam un1_rnd_out_i_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_12_cZ(.I0(pre_out_i[19:19]),.O(un1_rnd_out_i_axb_12));
defparam un1_rnd_out_i_axb_12_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_12_cZ(.I0(pre_out_r[19:19]),.O(un2_rnd_out_r_axb_12));
defparam un2_rnd_out_r_axb_12_cZ.INIT=2'h2;
  LUT4 un4_rnd_sat_out_i_3_cZ(.I0(pre_out_i[20:20]),.I1(pre_out_i[21:21]),.I2(pre_out_i[22:22]),.I3(pre_out_i[19:19]),.O(un4_rnd_sat_out_i_3));
defparam un4_rnd_sat_out_i_3_cZ.INIT=16'h8000;
  LUT4 un5_rnd_sat_out_r_3_cZ(.I0(pre_out_r[20:20]),.I1(pre_out_r[21:21]),.I2(pre_out_r[22:22]),.I3(pre_out_r[19:19]),.O(un5_rnd_sat_out_r_3));
defparam un5_rnd_sat_out_r_3_cZ.INIT=16'h8000;
  LUT3 un1_pos_out_r(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.O(un1_pos_out_r_0));
defparam un1_pos_out_r.INIT=8'h04;
  LUT3 un1_pos_out_i(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.O(un1_pos_out_i_0));
defparam un1_pos_out_i.INIT=8'h08;
  LUT6_L desc537(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r_s_12_2),.LO(pos_out_r[11:11]));
defparam desc537.INIT=64'hDBD0DBD00000D0D0;
  LUT6_L desc538(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i_s_12_2),.LO(pos_out_i[11:11]));
defparam desc538.INIT=64'hE7E0E7E00000E0E0;
  LUT6_L desc539(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[10:10]),.LO(pos_out_i_iv_i[10:10]));
defparam desc539.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc540(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[9:9]),.LO(pos_out_i_iv_i[9:9]));
defparam desc540.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc541(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[8:8]),.LO(pos_out_i_iv_i[8:8]));
defparam desc541.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc542(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[7:7]),.LO(pos_out_i_iv_i[7:7]));
defparam desc542.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc543(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[6:6]),.LO(pos_out_i_iv_i[6:6]));
defparam desc543.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc544(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[5:5]),.LO(pos_out_i_iv_i[5:5]));
defparam desc544.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc545(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[4:4]),.LO(pos_out_i_iv_i[4:4]));
defparam desc545.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc546(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[3:3]),.LO(pos_out_i_iv_i[3:3]));
defparam desc546.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc547(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[2:2]),.LO(pos_out_i_iv_i[2:2]));
defparam desc547.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc548(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_1),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[1:1]),.LO(pos_out_i_iv_i[1:1]));
defparam desc548.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc549(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(un1_rnd_out_i[0:0]),.I4(PATTERNDETECT_1),.I5(un4_rnd_sat_out_i_3),.LO(pos_out_i_iv_i[0:0]));
defparam desc549.INIT=64'hFF18FF1F1F181F1F;
  LUT6_L desc550(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[10:10]),.LO(pos_out_r_iv_i[10:10]));
defparam desc550.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc551(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[9:9]),.LO(pos_out_r_iv_i[9:9]));
defparam desc551.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc552(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[8:8]),.LO(pos_out_r_iv_i[8:8]));
defparam desc552.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc553(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[7:7]),.LO(pos_out_r_iv_i[7:7]));
defparam desc553.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc554(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[6:6]),.LO(pos_out_r_iv_i[6:6]));
defparam desc554.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc555(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[5:5]),.LO(pos_out_r_iv_i[5:5]));
defparam desc555.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc556(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[4:4]),.LO(pos_out_r_iv_i[4:4]));
defparam desc556.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc557(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[3:3]),.LO(pos_out_r_iv_i[3:3]));
defparam desc557.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc558(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[2:2]),.LO(pos_out_r_iv_i[2:2]));
defparam desc558.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc559(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_2),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[1:1]),.LO(pos_out_r_iv_i[1:1]));
defparam desc559.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc560(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(un2_rnd_out_r[0:0]),.I4(PATTERNDETECT_2),.I5(un5_rnd_sat_out_r_3),.LO(pos_out_r_iv_i[0:0]));
defparam desc560.INIT=64'hFF24FF2F2F242F2F;
  XORCY un1_rnd_out_i_s_12(.LI(un1_rnd_out_i_axb_12),.CI(un1_rnd_out_i_cry_11),.O(un1_rnd_out_i_s_12_2));
  XORCY un1_rnd_out_i_s_11(.LI(un1_rnd_out_i_axb_11),.CI(un1_rnd_out_i_cry_10),.O(un1_rnd_out_i[10:10]));
  MUXCY_L un1_rnd_out_i_cry_11_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_10),.S(un1_rnd_out_i_axb_11),.LO(un1_rnd_out_i_cry_11));
  XORCY un1_rnd_out_i_s_10(.LI(un1_rnd_out_i_axb_10),.CI(un1_rnd_out_i_cry_9),.O(un1_rnd_out_i[9:9]));
  MUXCY_L un1_rnd_out_i_cry_10_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_9),.S(un1_rnd_out_i_axb_10),.LO(un1_rnd_out_i_cry_10));
  XORCY un1_rnd_out_i_s_9(.LI(un1_rnd_out_i_axb_9),.CI(un1_rnd_out_i_cry_8),.O(un1_rnd_out_i[8:8]));
  MUXCY_L un1_rnd_out_i_cry_9_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_8),.S(un1_rnd_out_i_axb_9),.LO(un1_rnd_out_i_cry_9));
  XORCY un1_rnd_out_i_s_8(.LI(un1_rnd_out_i_axb_8),.CI(un1_rnd_out_i_cry_7),.O(un1_rnd_out_i[7:7]));
  MUXCY_L un1_rnd_out_i_cry_8_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_7),.S(un1_rnd_out_i_axb_8),.LO(un1_rnd_out_i_cry_8));
  XORCY un1_rnd_out_i_s_7(.LI(un1_rnd_out_i_axb_7),.CI(un1_rnd_out_i_cry_6),.O(un1_rnd_out_i[6:6]));
  MUXCY_L un1_rnd_out_i_cry_7_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_6),.S(un1_rnd_out_i_axb_7),.LO(un1_rnd_out_i_cry_7));
  XORCY un1_rnd_out_i_s_6(.LI(un1_rnd_out_i_axb_6),.CI(un1_rnd_out_i_cry_5),.O(un1_rnd_out_i[5:5]));
  MUXCY_L un1_rnd_out_i_cry_6_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_5),.S(un1_rnd_out_i_axb_6),.LO(un1_rnd_out_i_cry_6));
  XORCY un1_rnd_out_i_s_5(.LI(un1_rnd_out_i_axb_5),.CI(un1_rnd_out_i_cry_4),.O(un1_rnd_out_i[4:4]));
  MUXCY_L un1_rnd_out_i_cry_5_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_4),.S(un1_rnd_out_i_axb_5),.LO(un1_rnd_out_i_cry_5));
  XORCY un1_rnd_out_i_s_4(.LI(un1_rnd_out_i_axb_4),.CI(un1_rnd_out_i_cry_3),.O(un1_rnd_out_i[3:3]));
  MUXCY_L un1_rnd_out_i_cry_4_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_3),.S(un1_rnd_out_i_axb_4),.LO(un1_rnd_out_i_cry_4));
  XORCY un1_rnd_out_i_s_3(.LI(un1_rnd_out_i_axb_3),.CI(un1_rnd_out_i_cry_2),.O(un1_rnd_out_i[2:2]));
  MUXCY_L un1_rnd_out_i_cry_3_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_2),.S(un1_rnd_out_i_axb_3),.LO(un1_rnd_out_i_cry_3));
  XORCY un1_rnd_out_i_s_2(.LI(un1_rnd_out_i_axb_2),.CI(un1_rnd_out_i_cry_1),.O(un1_rnd_out_i[1:1]));
  MUXCY_L un1_rnd_out_i_cry_2_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_1),.S(un1_rnd_out_i_axb_2),.LO(un1_rnd_out_i_cry_2));
  XORCY un1_rnd_out_i_s_1(.LI(un1_rnd_out_i_axb_1),.CI(pre_out_i[7:7]),.O(un1_rnd_out_i[0:0]));
  MUXCY_L un1_rnd_out_i_cry_1_cZ(.DI(GND),.CI(pre_out_i[7:7]),.S(un1_rnd_out_i_axb_1),.LO(un1_rnd_out_i_cry_1));
  XORCY un2_rnd_out_r_s_12(.LI(un2_rnd_out_r_axb_12),.CI(un2_rnd_out_r_cry_11),.O(un2_rnd_out_r_s_12_2));
  XORCY un2_rnd_out_r_s_11(.LI(un2_rnd_out_r_axb_11),.CI(un2_rnd_out_r_cry_10),.O(un2_rnd_out_r[10:10]));
  MUXCY_L un2_rnd_out_r_cry_11_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_10),.S(un2_rnd_out_r_axb_11),.LO(un2_rnd_out_r_cry_11));
  XORCY un2_rnd_out_r_s_10(.LI(un2_rnd_out_r_axb_10),.CI(un2_rnd_out_r_cry_9),.O(un2_rnd_out_r[9:9]));
  MUXCY_L un2_rnd_out_r_cry_10_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_9),.S(un2_rnd_out_r_axb_10),.LO(un2_rnd_out_r_cry_10));
  XORCY un2_rnd_out_r_s_9(.LI(un2_rnd_out_r_axb_9),.CI(un2_rnd_out_r_cry_8),.O(un2_rnd_out_r[8:8]));
  MUXCY_L un2_rnd_out_r_cry_9_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_8),.S(un2_rnd_out_r_axb_9),.LO(un2_rnd_out_r_cry_9));
  XORCY un2_rnd_out_r_s_8(.LI(un2_rnd_out_r_axb_8),.CI(un2_rnd_out_r_cry_7),.O(un2_rnd_out_r[7:7]));
  MUXCY_L un2_rnd_out_r_cry_8_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_7),.S(un2_rnd_out_r_axb_8),.LO(un2_rnd_out_r_cry_8));
  XORCY un2_rnd_out_r_s_7(.LI(un2_rnd_out_r_axb_7),.CI(un2_rnd_out_r_cry_6),.O(un2_rnd_out_r[6:6]));
  MUXCY_L un2_rnd_out_r_cry_7_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_6),.S(un2_rnd_out_r_axb_7),.LO(un2_rnd_out_r_cry_7));
  XORCY un2_rnd_out_r_s_6(.LI(un2_rnd_out_r_axb_6),.CI(un2_rnd_out_r_cry_5),.O(un2_rnd_out_r[5:5]));
  MUXCY_L un2_rnd_out_r_cry_6_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_5),.S(un2_rnd_out_r_axb_6),.LO(un2_rnd_out_r_cry_6));
  XORCY un2_rnd_out_r_s_5(.LI(un2_rnd_out_r_axb_5),.CI(un2_rnd_out_r_cry_4),.O(un2_rnd_out_r[4:4]));
  MUXCY_L un2_rnd_out_r_cry_5_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_4),.S(un2_rnd_out_r_axb_5),.LO(un2_rnd_out_r_cry_5));
  XORCY un2_rnd_out_r_s_4(.LI(un2_rnd_out_r_axb_4),.CI(un2_rnd_out_r_cry_3),.O(un2_rnd_out_r[3:3]));
  MUXCY_L un2_rnd_out_r_cry_4_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_3),.S(un2_rnd_out_r_axb_4),.LO(un2_rnd_out_r_cry_4));
  XORCY un2_rnd_out_r_s_3(.LI(un2_rnd_out_r_axb_3),.CI(un2_rnd_out_r_cry_2),.O(un2_rnd_out_r[2:2]));
  MUXCY_L un2_rnd_out_r_cry_3_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_2),.S(un2_rnd_out_r_axb_3),.LO(un2_rnd_out_r_cry_3));
  XORCY un2_rnd_out_r_s_2(.LI(un2_rnd_out_r_axb_2),.CI(un2_rnd_out_r_cry_1),.O(un2_rnd_out_r[1:1]));
  MUXCY_L un2_rnd_out_r_cry_2_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_1),.S(un2_rnd_out_r_axb_2),.LO(un2_rnd_out_r_cry_2));
  XORCY un2_rnd_out_r_s_1(.LI(un2_rnd_out_r_axb_1),.CI(pre_out_r[7:7]),.O(un2_rnd_out_r[0:0]));
  MUXCY_L un2_rnd_out_r_cry_1_cZ(.DI(GND),.CI(pre_out_r[7:7]),.S(un2_rnd_out_r_axb_1),.LO(un2_rnd_out_r_cry_1));
  FDS desc561(.Q(out_i_vec_mult_1[11:11]),.D(pos_out_i[11:11]),.C(clk),.S(un1_pos_out_i_0));
  FDR desc562(.Q(out_i_vec_mult_1[10:10]),.D(pos_out_i_iv_i[10:10]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc563(.Q(out_i_vec_mult_1[9:9]),.D(pos_out_i_iv_i[9:9]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc564(.Q(out_i_vec_mult_1[8:8]),.D(pos_out_i_iv_i[8:8]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc565(.Q(out_i_vec_mult_1[7:7]),.D(pos_out_i_iv_i[7:7]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc566(.Q(out_i_vec_mult_1[6:6]),.D(pos_out_i_iv_i[6:6]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc567(.Q(out_i_vec_mult_1[5:5]),.D(pos_out_i_iv_i[5:5]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc568(.Q(out_i_vec_mult_1[4:4]),.D(pos_out_i_iv_i[4:4]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc569(.Q(out_i_vec_mult_1[3:3]),.D(pos_out_i_iv_i[3:3]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc570(.Q(out_i_vec_mult_1[2:2]),.D(pos_out_i_iv_i[2:2]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc571(.Q(out_i_vec_mult_1[1:1]),.D(pos_out_i_iv_i[1:1]),.C(clk),.R(un1_pos_out_i_0));
  FDR desc572(.Q(out_i_vec_mult_1[0:0]),.D(pos_out_i_iv_i[0:0]),.C(clk),.R(un1_pos_out_i_0));
  FDS desc573(.Q(out_r_vec_mult_1[11:11]),.D(pos_out_r[11:11]),.C(clk),.S(un1_pos_out_r_0));
  FDR desc574(.Q(out_r_vec_mult_1[10:10]),.D(pos_out_r_iv_i[10:10]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc575(.Q(out_r_vec_mult_1[9:9]),.D(pos_out_r_iv_i[9:9]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc576(.Q(out_r_vec_mult_1[8:8]),.D(pos_out_r_iv_i[8:8]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc577(.Q(out_r_vec_mult_1[7:7]),.D(pos_out_r_iv_i[7:7]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc578(.Q(out_r_vec_mult_1[6:6]),.D(pos_out_r_iv_i[6:6]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc579(.Q(out_r_vec_mult_1[5:5]),.D(pos_out_r_iv_i[5:5]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc580(.Q(out_r_vec_mult_1[4:4]),.D(pos_out_r_iv_i[4:4]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc581(.Q(out_r_vec_mult_1[3:3]),.D(pos_out_r_iv_i[3:3]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc582(.Q(out_r_vec_mult_1[2:2]),.D(pos_out_r_iv_i[2:2]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc583(.Q(out_r_vec_mult_1[1:1]),.D(pos_out_r_iv_i[1:1]),.C(clk),.R(un1_pos_out_r_0));
  FDR desc584(.Q(out_r_vec_mult_1[0:0]),.D(pos_out_r_iv_i[0:0]),.C(clk),.R(un1_pos_out_r_0));
  mult_pipe_8_inj mult1(.mult1_out_23(mult1_out[23:23]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_20_0(P_uc_20_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  mult_pipe_9_inj mult2(.mult2_out_23(mult2_out[23:23]),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_10_inj mult3(.mult3_out_23(mult3_out[23:23]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_11_inj mult4(.mult4_out_23(mult4_out[23:23]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_23_0(P_uc_23_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  add_subZ2_2_inj sub(.pre_out_r(pre_out_r[23:7]),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_20_0(P_uc_20_0[47:24]),.PATTERNDETECT_2(PATTERNDETECT_2),.clk(clk));
  add_subZ1_2_inj add(.pre_out_i(pre_out_i[23:7]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_23_0(P_uc_23_0[47:24]),.PATTERNDETECT_1(PATTERNDETECT_1),.clk(clk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module desc591_inj (out_i_vec_mult_0,out_r_vec_mult_0,out_inner_prod_r,vec_out_r_AQ_0,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,vec_out_i_AQ_0,out_inner_prod_i,in_b_i_reg,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output [11:0] out_i_vec_mult_0 ;
output [11:0] out_r_vec_mult_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_0 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input [11:0] vec_out_i_AQ_0 ;
input [11:0] out_inner_prod_i ;
input [11:0] in_b_i_reg ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [23:7] pre_out_r ;
wire [23:7] pre_out_i ;
wire [23:23] mult2_out ;
wire [23:23] mult1_out ;
wire [23:23] mult3_out ;
wire [23:23] mult4_out ;
wire [11:11] pos_out_r ;
wire [11:11] pos_out_i ;
wire [10:0] un1_rnd_out_i ;
wire [10:0] pos_out_i_iv_i ;
wire [10:0] un2_rnd_out_r ;
wire [10:0] pos_out_r_iv_i ;
wire [23:0] mult1_out_0 ;
wire [47:24] P_uc_16_0 ;
wire [23:0] mult4_out_0 ;
wire [47:24] P_uc_19_0 ;
wire un2_rnd_out_r_axb_1 ;
wire un2_rnd_out_r_axb_2 ;
wire un2_rnd_out_r_axb_3 ;
wire un2_rnd_out_r_axb_4 ;
wire un2_rnd_out_r_axb_5 ;
wire un2_rnd_out_r_axb_6 ;
wire un2_rnd_out_r_axb_7 ;
wire un2_rnd_out_r_axb_8 ;
wire un2_rnd_out_r_axb_9 ;
wire un2_rnd_out_r_axb_10 ;
wire un2_rnd_out_r_axb_11 ;
wire un1_rnd_out_i_axb_1 ;
wire un1_rnd_out_i_axb_2 ;
wire un1_rnd_out_i_axb_3 ;
wire un1_rnd_out_i_axb_4 ;
wire un1_rnd_out_i_axb_5 ;
wire un1_rnd_out_i_axb_6 ;
wire un1_rnd_out_i_axb_7 ;
wire un1_rnd_out_i_axb_8 ;
wire un1_rnd_out_i_axb_9 ;
wire un1_rnd_out_i_axb_10 ;
wire un1_rnd_out_i_axb_11 ;
wire un1_rnd_out_i_axb_12 ;
wire un2_rnd_out_r_axb_12 ;
wire un4_rnd_sat_out_i_3 ;
wire un5_rnd_sat_out_r_3 ;
wire un1_pos_out_r_1 ;
wire un1_pos_out_i_1 ;
wire PATTERNDETECT_0 ;
wire un2_rnd_out_r_s_12_0 ;
wire PATTERNDETECT ;
wire un1_rnd_out_i_s_12_0 ;
wire un1_rnd_out_i_cry_11 ;
wire un1_rnd_out_i_cry_10 ;
wire GND ;
wire un1_rnd_out_i_cry_9 ;
wire un1_rnd_out_i_cry_8 ;
wire un1_rnd_out_i_cry_7 ;
wire un1_rnd_out_i_cry_6 ;
wire un1_rnd_out_i_cry_5 ;
wire un1_rnd_out_i_cry_4 ;
wire un1_rnd_out_i_cry_3 ;
wire un1_rnd_out_i_cry_2 ;
wire un1_rnd_out_i_cry_1 ;
wire un2_rnd_out_r_cry_11 ;
wire un2_rnd_out_r_cry_10 ;
wire un2_rnd_out_r_cry_9 ;
wire un2_rnd_out_r_cry_8 ;
wire un2_rnd_out_r_cry_7 ;
wire un2_rnd_out_r_cry_6 ;
wire un2_rnd_out_r_cry_5 ;
wire un2_rnd_out_r_cry_4 ;
wire un2_rnd_out_r_cry_3 ;
wire un2_rnd_out_r_cry_2 ;
wire un2_rnd_out_r_cry_1 ;
wire VCC ;
// instances
  LUT1 un2_rnd_out_r_axb_1_cZ(.I0(pre_out_r[8:8]),.O(un2_rnd_out_r_axb_1));
defparam un2_rnd_out_r_axb_1_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_2_cZ(.I0(pre_out_r[9:9]),.O(un2_rnd_out_r_axb_2));
defparam un2_rnd_out_r_axb_2_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_3_cZ(.I0(pre_out_r[10:10]),.O(un2_rnd_out_r_axb_3));
defparam un2_rnd_out_r_axb_3_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_4_cZ(.I0(pre_out_r[11:11]),.O(un2_rnd_out_r_axb_4));
defparam un2_rnd_out_r_axb_4_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_5_cZ(.I0(pre_out_r[12:12]),.O(un2_rnd_out_r_axb_5));
defparam un2_rnd_out_r_axb_5_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_6_cZ(.I0(pre_out_r[13:13]),.O(un2_rnd_out_r_axb_6));
defparam un2_rnd_out_r_axb_6_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_7_cZ(.I0(pre_out_r[14:14]),.O(un2_rnd_out_r_axb_7));
defparam un2_rnd_out_r_axb_7_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_8_cZ(.I0(pre_out_r[15:15]),.O(un2_rnd_out_r_axb_8));
defparam un2_rnd_out_r_axb_8_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_9_cZ(.I0(pre_out_r[16:16]),.O(un2_rnd_out_r_axb_9));
defparam un2_rnd_out_r_axb_9_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_10_cZ(.I0(pre_out_r[17:17]),.O(un2_rnd_out_r_axb_10));
defparam un2_rnd_out_r_axb_10_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_11_cZ(.I0(pre_out_r[18:18]),.O(un2_rnd_out_r_axb_11));
defparam un2_rnd_out_r_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_1_cZ(.I0(pre_out_i[8:8]),.O(un1_rnd_out_i_axb_1));
defparam un1_rnd_out_i_axb_1_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_2_cZ(.I0(pre_out_i[9:9]),.O(un1_rnd_out_i_axb_2));
defparam un1_rnd_out_i_axb_2_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_3_cZ(.I0(pre_out_i[10:10]),.O(un1_rnd_out_i_axb_3));
defparam un1_rnd_out_i_axb_3_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_4_cZ(.I0(pre_out_i[11:11]),.O(un1_rnd_out_i_axb_4));
defparam un1_rnd_out_i_axb_4_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_5_cZ(.I0(pre_out_i[12:12]),.O(un1_rnd_out_i_axb_5));
defparam un1_rnd_out_i_axb_5_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_6_cZ(.I0(pre_out_i[13:13]),.O(un1_rnd_out_i_axb_6));
defparam un1_rnd_out_i_axb_6_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_7_cZ(.I0(pre_out_i[14:14]),.O(un1_rnd_out_i_axb_7));
defparam un1_rnd_out_i_axb_7_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_8_cZ(.I0(pre_out_i[15:15]),.O(un1_rnd_out_i_axb_8));
defparam un1_rnd_out_i_axb_8_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_9_cZ(.I0(pre_out_i[16:16]),.O(un1_rnd_out_i_axb_9));
defparam un1_rnd_out_i_axb_9_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_10_cZ(.I0(pre_out_i[17:17]),.O(un1_rnd_out_i_axb_10));
defparam un1_rnd_out_i_axb_10_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_11_cZ(.I0(pre_out_i[18:18]),.O(un1_rnd_out_i_axb_11));
defparam un1_rnd_out_i_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_12_cZ(.I0(pre_out_i[19:19]),.O(un1_rnd_out_i_axb_12));
defparam un1_rnd_out_i_axb_12_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_12_cZ(.I0(pre_out_r[19:19]),.O(un2_rnd_out_r_axb_12));
defparam un2_rnd_out_r_axb_12_cZ.INIT=2'h2;
  LUT4 un4_rnd_sat_out_i_3_cZ(.I0(pre_out_i[20:20]),.I1(pre_out_i[21:21]),.I2(pre_out_i[22:22]),.I3(pre_out_i[19:19]),.O(un4_rnd_sat_out_i_3));
defparam un4_rnd_sat_out_i_3_cZ.INIT=16'h8000;
  LUT4 un5_rnd_sat_out_r_3_cZ(.I0(pre_out_r[20:20]),.I1(pre_out_r[21:21]),.I2(pre_out_r[22:22]),.I3(pre_out_r[19:19]),.O(un5_rnd_sat_out_r_3));
defparam un5_rnd_sat_out_r_3_cZ.INIT=16'h8000;
  LUT3 un1_pos_out_r(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.O(un1_pos_out_r_1));
defparam un1_pos_out_r.INIT=8'h04;
  LUT3 un1_pos_out_i(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.O(un1_pos_out_i_1));
defparam un1_pos_out_i.INIT=8'h08;
  LUT6_L desc592(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r_s_12_0),.LO(pos_out_r[11:11]));
defparam desc592.INIT=64'hDBD0DBD00000D0D0;
  LUT6_L desc593(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i_s_12_0),.LO(pos_out_i[11:11]));
defparam desc593.INIT=64'hE7E0E7E00000E0E0;
  LUT6_L desc594(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[10:10]),.LO(pos_out_i_iv_i[10:10]));
defparam desc594.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc595(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[9:9]),.LO(pos_out_i_iv_i[9:9]));
defparam desc595.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc596(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[8:8]),.LO(pos_out_i_iv_i[8:8]));
defparam desc596.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc597(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[7:7]),.LO(pos_out_i_iv_i[7:7]));
defparam desc597.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc598(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[6:6]),.LO(pos_out_i_iv_i[6:6]));
defparam desc598.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc599(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[5:5]),.LO(pos_out_i_iv_i[5:5]));
defparam desc599.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc600(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[4:4]),.LO(pos_out_i_iv_i[4:4]));
defparam desc600.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc601(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[3:3]),.LO(pos_out_i_iv_i[3:3]));
defparam desc601.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc602(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[2:2]),.LO(pos_out_i_iv_i[2:2]));
defparam desc602.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc603(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[1:1]),.LO(pos_out_i_iv_i[1:1]));
defparam desc603.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc604(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(un1_rnd_out_i[0:0]),.I4(PATTERNDETECT),.I5(un4_rnd_sat_out_i_3),.LO(pos_out_i_iv_i[0:0]));
defparam desc604.INIT=64'hFF18FF1F1F181F1F;
  LUT6_L desc605(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[10:10]),.LO(pos_out_r_iv_i[10:10]));
defparam desc605.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc606(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[9:9]),.LO(pos_out_r_iv_i[9:9]));
defparam desc606.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc607(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[8:8]),.LO(pos_out_r_iv_i[8:8]));
defparam desc607.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc608(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[7:7]),.LO(pos_out_r_iv_i[7:7]));
defparam desc608.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc609(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[6:6]),.LO(pos_out_r_iv_i[6:6]));
defparam desc609.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc610(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[5:5]),.LO(pos_out_r_iv_i[5:5]));
defparam desc610.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc611(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[4:4]),.LO(pos_out_r_iv_i[4:4]));
defparam desc611.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc612(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[3:3]),.LO(pos_out_r_iv_i[3:3]));
defparam desc612.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc613(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[2:2]),.LO(pos_out_r_iv_i[2:2]));
defparam desc613.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc614(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_0),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[1:1]),.LO(pos_out_r_iv_i[1:1]));
defparam desc614.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc615(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(un2_rnd_out_r[0:0]),.I4(PATTERNDETECT_0),.I5(un5_rnd_sat_out_r_3),.LO(pos_out_r_iv_i[0:0]));
defparam desc615.INIT=64'hFF24FF2F2F242F2F;
  XORCY un1_rnd_out_i_s_12(.LI(un1_rnd_out_i_axb_12),.CI(un1_rnd_out_i_cry_11),.O(un1_rnd_out_i_s_12_0));
  XORCY un1_rnd_out_i_s_11(.LI(un1_rnd_out_i_axb_11),.CI(un1_rnd_out_i_cry_10),.O(un1_rnd_out_i[10:10]));
  MUXCY_L un1_rnd_out_i_cry_11_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_10),.S(un1_rnd_out_i_axb_11),.LO(un1_rnd_out_i_cry_11));
  XORCY un1_rnd_out_i_s_10(.LI(un1_rnd_out_i_axb_10),.CI(un1_rnd_out_i_cry_9),.O(un1_rnd_out_i[9:9]));
  MUXCY_L un1_rnd_out_i_cry_10_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_9),.S(un1_rnd_out_i_axb_10),.LO(un1_rnd_out_i_cry_10));
  XORCY un1_rnd_out_i_s_9(.LI(un1_rnd_out_i_axb_9),.CI(un1_rnd_out_i_cry_8),.O(un1_rnd_out_i[8:8]));
  MUXCY_L un1_rnd_out_i_cry_9_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_8),.S(un1_rnd_out_i_axb_9),.LO(un1_rnd_out_i_cry_9));
  XORCY un1_rnd_out_i_s_8(.LI(un1_rnd_out_i_axb_8),.CI(un1_rnd_out_i_cry_7),.O(un1_rnd_out_i[7:7]));
  MUXCY_L un1_rnd_out_i_cry_8_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_7),.S(un1_rnd_out_i_axb_8),.LO(un1_rnd_out_i_cry_8));
  XORCY un1_rnd_out_i_s_7(.LI(un1_rnd_out_i_axb_7),.CI(un1_rnd_out_i_cry_6),.O(un1_rnd_out_i[6:6]));
  MUXCY_L un1_rnd_out_i_cry_7_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_6),.S(un1_rnd_out_i_axb_7),.LO(un1_rnd_out_i_cry_7));
  XORCY un1_rnd_out_i_s_6(.LI(un1_rnd_out_i_axb_6),.CI(un1_rnd_out_i_cry_5),.O(un1_rnd_out_i[5:5]));
  MUXCY_L un1_rnd_out_i_cry_6_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_5),.S(un1_rnd_out_i_axb_6),.LO(un1_rnd_out_i_cry_6));
  XORCY un1_rnd_out_i_s_5(.LI(un1_rnd_out_i_axb_5),.CI(un1_rnd_out_i_cry_4),.O(un1_rnd_out_i[4:4]));
  MUXCY_L un1_rnd_out_i_cry_5_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_4),.S(un1_rnd_out_i_axb_5),.LO(un1_rnd_out_i_cry_5));
  XORCY un1_rnd_out_i_s_4(.LI(un1_rnd_out_i_axb_4),.CI(un1_rnd_out_i_cry_3),.O(un1_rnd_out_i[3:3]));
  MUXCY_L un1_rnd_out_i_cry_4_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_3),.S(un1_rnd_out_i_axb_4),.LO(un1_rnd_out_i_cry_4));
  XORCY un1_rnd_out_i_s_3(.LI(un1_rnd_out_i_axb_3),.CI(un1_rnd_out_i_cry_2),.O(un1_rnd_out_i[2:2]));
  MUXCY_L un1_rnd_out_i_cry_3_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_2),.S(un1_rnd_out_i_axb_3),.LO(un1_rnd_out_i_cry_3));
  XORCY un1_rnd_out_i_s_2(.LI(un1_rnd_out_i_axb_2),.CI(un1_rnd_out_i_cry_1),.O(un1_rnd_out_i[1:1]));
  MUXCY_L un1_rnd_out_i_cry_2_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_1),.S(un1_rnd_out_i_axb_2),.LO(un1_rnd_out_i_cry_2));
  XORCY un1_rnd_out_i_s_1(.LI(un1_rnd_out_i_axb_1),.CI(pre_out_i[7:7]),.O(un1_rnd_out_i[0:0]));
  MUXCY_L un1_rnd_out_i_cry_1_cZ(.DI(GND),.CI(pre_out_i[7:7]),.S(un1_rnd_out_i_axb_1),.LO(un1_rnd_out_i_cry_1));
  XORCY un2_rnd_out_r_s_12(.LI(un2_rnd_out_r_axb_12),.CI(un2_rnd_out_r_cry_11),.O(un2_rnd_out_r_s_12_0));
  XORCY un2_rnd_out_r_s_11(.LI(un2_rnd_out_r_axb_11),.CI(un2_rnd_out_r_cry_10),.O(un2_rnd_out_r[10:10]));
  MUXCY_L un2_rnd_out_r_cry_11_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_10),.S(un2_rnd_out_r_axb_11),.LO(un2_rnd_out_r_cry_11));
  XORCY un2_rnd_out_r_s_10(.LI(un2_rnd_out_r_axb_10),.CI(un2_rnd_out_r_cry_9),.O(un2_rnd_out_r[9:9]));
  MUXCY_L un2_rnd_out_r_cry_10_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_9),.S(un2_rnd_out_r_axb_10),.LO(un2_rnd_out_r_cry_10));
  XORCY un2_rnd_out_r_s_9(.LI(un2_rnd_out_r_axb_9),.CI(un2_rnd_out_r_cry_8),.O(un2_rnd_out_r[8:8]));
  MUXCY_L un2_rnd_out_r_cry_9_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_8),.S(un2_rnd_out_r_axb_9),.LO(un2_rnd_out_r_cry_9));
  XORCY un2_rnd_out_r_s_8(.LI(un2_rnd_out_r_axb_8),.CI(un2_rnd_out_r_cry_7),.O(un2_rnd_out_r[7:7]));
  MUXCY_L un2_rnd_out_r_cry_8_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_7),.S(un2_rnd_out_r_axb_8),.LO(un2_rnd_out_r_cry_8));
  XORCY un2_rnd_out_r_s_7(.LI(un2_rnd_out_r_axb_7),.CI(un2_rnd_out_r_cry_6),.O(un2_rnd_out_r[6:6]));
  MUXCY_L un2_rnd_out_r_cry_7_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_6),.S(un2_rnd_out_r_axb_7),.LO(un2_rnd_out_r_cry_7));
  XORCY un2_rnd_out_r_s_6(.LI(un2_rnd_out_r_axb_6),.CI(un2_rnd_out_r_cry_5),.O(un2_rnd_out_r[5:5]));
  MUXCY_L un2_rnd_out_r_cry_6_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_5),.S(un2_rnd_out_r_axb_6),.LO(un2_rnd_out_r_cry_6));
  XORCY un2_rnd_out_r_s_5(.LI(un2_rnd_out_r_axb_5),.CI(un2_rnd_out_r_cry_4),.O(un2_rnd_out_r[4:4]));
  MUXCY_L un2_rnd_out_r_cry_5_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_4),.S(un2_rnd_out_r_axb_5),.LO(un2_rnd_out_r_cry_5));
  XORCY un2_rnd_out_r_s_4(.LI(un2_rnd_out_r_axb_4),.CI(un2_rnd_out_r_cry_3),.O(un2_rnd_out_r[3:3]));
  MUXCY_L un2_rnd_out_r_cry_4_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_3),.S(un2_rnd_out_r_axb_4),.LO(un2_rnd_out_r_cry_4));
  XORCY un2_rnd_out_r_s_3(.LI(un2_rnd_out_r_axb_3),.CI(un2_rnd_out_r_cry_2),.O(un2_rnd_out_r[2:2]));
  MUXCY_L un2_rnd_out_r_cry_3_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_2),.S(un2_rnd_out_r_axb_3),.LO(un2_rnd_out_r_cry_3));
  XORCY un2_rnd_out_r_s_2(.LI(un2_rnd_out_r_axb_2),.CI(un2_rnd_out_r_cry_1),.O(un2_rnd_out_r[1:1]));
  MUXCY_L un2_rnd_out_r_cry_2_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_1),.S(un2_rnd_out_r_axb_2),.LO(un2_rnd_out_r_cry_2));
  XORCY un2_rnd_out_r_s_1(.LI(un2_rnd_out_r_axb_1),.CI(pre_out_r[7:7]),.O(un2_rnd_out_r[0:0]));
  MUXCY_L un2_rnd_out_r_cry_1_cZ(.DI(GND),.CI(pre_out_r[7:7]),.S(un2_rnd_out_r_axb_1),.LO(un2_rnd_out_r_cry_1));
  FDS desc616(.Q(out_i_vec_mult_0[11:11]),.D(pos_out_i[11:11]),.C(clk),.S(un1_pos_out_i_1));
  FDR desc617(.Q(out_i_vec_mult_0[10:10]),.D(pos_out_i_iv_i[10:10]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc618(.Q(out_i_vec_mult_0[9:9]),.D(pos_out_i_iv_i[9:9]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc619(.Q(out_i_vec_mult_0[8:8]),.D(pos_out_i_iv_i[8:8]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc620(.Q(out_i_vec_mult_0[7:7]),.D(pos_out_i_iv_i[7:7]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc621(.Q(out_i_vec_mult_0[6:6]),.D(pos_out_i_iv_i[6:6]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc622(.Q(out_i_vec_mult_0[5:5]),.D(pos_out_i_iv_i[5:5]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc623(.Q(out_i_vec_mult_0[4:4]),.D(pos_out_i_iv_i[4:4]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc624(.Q(out_i_vec_mult_0[3:3]),.D(pos_out_i_iv_i[3:3]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc625(.Q(out_i_vec_mult_0[2:2]),.D(pos_out_i_iv_i[2:2]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc626(.Q(out_i_vec_mult_0[1:1]),.D(pos_out_i_iv_i[1:1]),.C(clk),.R(un1_pos_out_i_1));
  FDR desc627(.Q(out_i_vec_mult_0[0:0]),.D(pos_out_i_iv_i[0:0]),.C(clk),.R(un1_pos_out_i_1));
  FDS desc628(.Q(out_r_vec_mult_0[11:11]),.D(pos_out_r[11:11]),.C(clk),.S(un1_pos_out_r_1));
  FDR desc629(.Q(out_r_vec_mult_0[10:10]),.D(pos_out_r_iv_i[10:10]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc630(.Q(out_r_vec_mult_0[9:9]),.D(pos_out_r_iv_i[9:9]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc631(.Q(out_r_vec_mult_0[8:8]),.D(pos_out_r_iv_i[8:8]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc632(.Q(out_r_vec_mult_0[7:7]),.D(pos_out_r_iv_i[7:7]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc633(.Q(out_r_vec_mult_0[6:6]),.D(pos_out_r_iv_i[6:6]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc634(.Q(out_r_vec_mult_0[5:5]),.D(pos_out_r_iv_i[5:5]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc635(.Q(out_r_vec_mult_0[4:4]),.D(pos_out_r_iv_i[4:4]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc636(.Q(out_r_vec_mult_0[3:3]),.D(pos_out_r_iv_i[3:3]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc637(.Q(out_r_vec_mult_0[2:2]),.D(pos_out_r_iv_i[2:2]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc638(.Q(out_r_vec_mult_0[1:1]),.D(pos_out_r_iv_i[1:1]),.C(clk),.R(un1_pos_out_r_1));
  FDR desc639(.Q(out_r_vec_mult_0[0:0]),.D(pos_out_r_iv_i[0:0]),.C(clk),.R(un1_pos_out_r_1));
  mult_pipe_12_inj mult1(.mult1_out_23(mult1_out[23:23]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_16_0(P_uc_16_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  mult_pipe_13_inj mult2(.mult2_out_23(mult2_out[23:23]),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_14_inj mult3(.mult3_out_23(mult3_out[23:23]),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_15_inj mult4(.mult4_out_23(mult4_out[23:23]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_19_0(P_uc_19_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  add_subZ2_3_inj sub(.pre_out_r(pre_out_r[23:7]),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_16_0(P_uc_16_0[47:24]),.PATTERNDETECT_0(PATTERNDETECT_0),.clk(clk));
  add_subZ1_3_inj add(.pre_out_i(pre_out_i[23:7]),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_19_0(P_uc_19_0[47:24]),.PATTERNDETECT(PATTERNDETECT),.clk(clk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module desc646_inj (out_i_vec_mult_3,out_r_vec_mult_3,out_inner_prod_r,vec_out_r_AQ_3,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,vec_out_i_AQ_3,out_inner_prod_i,in_b_i_reg,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output [11:0] out_i_vec_mult_3 ;
output [11:0] out_r_vec_mult_3 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_3 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input [11:0] vec_out_i_AQ_3 ;
input [11:0] out_inner_prod_i ;
input [11:0] in_b_i_reg ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [23:7] pre_out_r ;
wire [23:7] pre_out_i ;
wire [23:23] mult2_out ;
wire [23:23] mult1_out ;
wire [23:23] mult3_out ;
wire [23:23] mult4_out ;
wire [11:11] pos_out_r ;
wire [11:11] pos_out_i ;
wire [10:0] un1_rnd_out_i ;
wire [10:0] pos_out_i_iv_i ;
wire [10:0] un2_rnd_out_r ;
wire [10:0] pos_out_r_iv_i ;
wire [23:0] mult1_out_0 ;
wire [47:24] P_uc_28_0 ;
wire [23:0] mult4_out_0 ;
wire [47:24] P_uc_31_0 ;
wire un2_rnd_out_r_axb_1 ;
wire un2_rnd_out_r_axb_2 ;
wire un2_rnd_out_r_axb_3 ;
wire un2_rnd_out_r_axb_4 ;
wire un2_rnd_out_r_axb_5 ;
wire un2_rnd_out_r_axb_6 ;
wire un2_rnd_out_r_axb_7 ;
wire un2_rnd_out_r_axb_8 ;
wire un2_rnd_out_r_axb_9 ;
wire un2_rnd_out_r_axb_10 ;
wire un2_rnd_out_r_axb_11 ;
wire un1_rnd_out_i_axb_1 ;
wire un1_rnd_out_i_axb_2 ;
wire un1_rnd_out_i_axb_3 ;
wire un1_rnd_out_i_axb_4 ;
wire un1_rnd_out_i_axb_5 ;
wire un1_rnd_out_i_axb_6 ;
wire un1_rnd_out_i_axb_7 ;
wire un1_rnd_out_i_axb_8 ;
wire un1_rnd_out_i_axb_9 ;
wire un1_rnd_out_i_axb_10 ;
wire un1_rnd_out_i_axb_11 ;
wire un1_rnd_out_i_axb_12 ;
wire un2_rnd_out_r_axb_12 ;
wire un4_rnd_sat_out_i_3 ;
wire un5_rnd_sat_out_r_3 ;
wire un1_pos_out_r_2 ;
wire un1_pos_out_i_2 ;
wire PATTERNDETECT_6 ;
wire un2_rnd_out_r_s_12_1 ;
wire PATTERNDETECT_5 ;
wire un1_rnd_out_i_s_12_1 ;
wire un1_rnd_out_i_cry_11 ;
wire un1_rnd_out_i_cry_10 ;
wire GND ;
wire un1_rnd_out_i_cry_9 ;
wire un1_rnd_out_i_cry_8 ;
wire un1_rnd_out_i_cry_7 ;
wire un1_rnd_out_i_cry_6 ;
wire un1_rnd_out_i_cry_5 ;
wire un1_rnd_out_i_cry_4 ;
wire un1_rnd_out_i_cry_3 ;
wire un1_rnd_out_i_cry_2 ;
wire un1_rnd_out_i_cry_1 ;
wire un2_rnd_out_r_cry_11 ;
wire un2_rnd_out_r_cry_10 ;
wire un2_rnd_out_r_cry_9 ;
wire un2_rnd_out_r_cry_8 ;
wire un2_rnd_out_r_cry_7 ;
wire un2_rnd_out_r_cry_6 ;
wire un2_rnd_out_r_cry_5 ;
wire un2_rnd_out_r_cry_4 ;
wire un2_rnd_out_r_cry_3 ;
wire un2_rnd_out_r_cry_2 ;
wire un2_rnd_out_r_cry_1 ;
wire VCC ;
// instances
  LUT1 un2_rnd_out_r_axb_1_cZ(.I0(pre_out_r[8:8]),.O(un2_rnd_out_r_axb_1));
defparam un2_rnd_out_r_axb_1_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_2_cZ(.I0(pre_out_r[9:9]),.O(un2_rnd_out_r_axb_2));
defparam un2_rnd_out_r_axb_2_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_3_cZ(.I0(pre_out_r[10:10]),.O(un2_rnd_out_r_axb_3));
defparam un2_rnd_out_r_axb_3_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_4_cZ(.I0(pre_out_r[11:11]),.O(un2_rnd_out_r_axb_4));
defparam un2_rnd_out_r_axb_4_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_5_cZ(.I0(pre_out_r[12:12]),.O(un2_rnd_out_r_axb_5));
defparam un2_rnd_out_r_axb_5_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_6_cZ(.I0(pre_out_r[13:13]),.O(un2_rnd_out_r_axb_6));
defparam un2_rnd_out_r_axb_6_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_7_cZ(.I0(pre_out_r[14:14]),.O(un2_rnd_out_r_axb_7));
defparam un2_rnd_out_r_axb_7_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_8_cZ(.I0(pre_out_r[15:15]),.O(un2_rnd_out_r_axb_8));
defparam un2_rnd_out_r_axb_8_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_9_cZ(.I0(pre_out_r[16:16]),.O(un2_rnd_out_r_axb_9));
defparam un2_rnd_out_r_axb_9_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_10_cZ(.I0(pre_out_r[17:17]),.O(un2_rnd_out_r_axb_10));
defparam un2_rnd_out_r_axb_10_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_11_cZ(.I0(pre_out_r[18:18]),.O(un2_rnd_out_r_axb_11));
defparam un2_rnd_out_r_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_1_cZ(.I0(pre_out_i[8:8]),.O(un1_rnd_out_i_axb_1));
defparam un1_rnd_out_i_axb_1_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_2_cZ(.I0(pre_out_i[9:9]),.O(un1_rnd_out_i_axb_2));
defparam un1_rnd_out_i_axb_2_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_3_cZ(.I0(pre_out_i[10:10]),.O(un1_rnd_out_i_axb_3));
defparam un1_rnd_out_i_axb_3_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_4_cZ(.I0(pre_out_i[11:11]),.O(un1_rnd_out_i_axb_4));
defparam un1_rnd_out_i_axb_4_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_5_cZ(.I0(pre_out_i[12:12]),.O(un1_rnd_out_i_axb_5));
defparam un1_rnd_out_i_axb_5_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_6_cZ(.I0(pre_out_i[13:13]),.O(un1_rnd_out_i_axb_6));
defparam un1_rnd_out_i_axb_6_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_7_cZ(.I0(pre_out_i[14:14]),.O(un1_rnd_out_i_axb_7));
defparam un1_rnd_out_i_axb_7_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_8_cZ(.I0(pre_out_i[15:15]),.O(un1_rnd_out_i_axb_8));
defparam un1_rnd_out_i_axb_8_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_9_cZ(.I0(pre_out_i[16:16]),.O(un1_rnd_out_i_axb_9));
defparam un1_rnd_out_i_axb_9_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_10_cZ(.I0(pre_out_i[17:17]),.O(un1_rnd_out_i_axb_10));
defparam un1_rnd_out_i_axb_10_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_11_cZ(.I0(pre_out_i[18:18]),.O(un1_rnd_out_i_axb_11));
defparam un1_rnd_out_i_axb_11_cZ.INIT=2'h2;
  LUT1 un1_rnd_out_i_axb_12_cZ(.I0(pre_out_i[19:19]),.O(un1_rnd_out_i_axb_12));
defparam un1_rnd_out_i_axb_12_cZ.INIT=2'h2;
  LUT1 un2_rnd_out_r_axb_12_cZ(.I0(pre_out_r[19:19]),.O(un2_rnd_out_r_axb_12));
defparam un2_rnd_out_r_axb_12_cZ.INIT=2'h2;
  LUT4 un4_rnd_sat_out_i_3_cZ(.I0(pre_out_i[20:20]),.I1(pre_out_i[21:21]),.I2(pre_out_i[22:22]),.I3(pre_out_i[19:19]),.O(un4_rnd_sat_out_i_3));
defparam un4_rnd_sat_out_i_3_cZ.INIT=16'h8000;
  LUT4 un5_rnd_sat_out_r_3_cZ(.I0(pre_out_r[20:20]),.I1(pre_out_r[21:21]),.I2(pre_out_r[22:22]),.I3(pre_out_r[19:19]),.O(un5_rnd_sat_out_r_3));
defparam un5_rnd_sat_out_r_3_cZ.INIT=16'h8000;
  LUT3 un1_pos_out_r(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.O(un1_pos_out_r_2));
defparam un1_pos_out_r.INIT=8'h04;
  LUT3 un1_pos_out_i(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.O(un1_pos_out_i_2));
defparam un1_pos_out_i.INIT=8'h08;
  LUT6_L desc647(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r_s_12_1),.LO(pos_out_r[11:11]));
defparam desc647.INIT=64'hDBD0DBD00000D0D0;
  LUT6_L desc648(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i_s_12_1),.LO(pos_out_i[11:11]));
defparam desc648.INIT=64'hE7E0E7E00000E0E0;
  LUT6_L desc649(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[10:10]),.LO(pos_out_i_iv_i[10:10]));
defparam desc649.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc650(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[9:9]),.LO(pos_out_i_iv_i[9:9]));
defparam desc650.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc651(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[8:8]),.LO(pos_out_i_iv_i[8:8]));
defparam desc651.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc652(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[7:7]),.LO(pos_out_i_iv_i[7:7]));
defparam desc652.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc653(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[6:6]),.LO(pos_out_i_iv_i[6:6]));
defparam desc653.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc654(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[5:5]),.LO(pos_out_i_iv_i[5:5]));
defparam desc654.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc655(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[4:4]),.LO(pos_out_i_iv_i[4:4]));
defparam desc655.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc656(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[3:3]),.LO(pos_out_i_iv_i[3:3]));
defparam desc656.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc657(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[2:2]),.LO(pos_out_i_iv_i[2:2]));
defparam desc657.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc658(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(PATTERNDETECT_5),.I4(un4_rnd_sat_out_i_3),.I5(un1_rnd_out_i[1:1]),.LO(pos_out_i_iv_i[1:1]));
defparam desc658.INIT=64'hFFFF1F1F181F181F;
  LUT6_L desc659(.I0(mult3_out[23:23]),.I1(mult4_out[23:23]),.I2(pre_out_i[23:23]),.I3(un1_rnd_out_i[0:0]),.I4(PATTERNDETECT_5),.I5(un4_rnd_sat_out_i_3),.LO(pos_out_i_iv_i[0:0]));
defparam desc659.INIT=64'hFF18FF1F1F181F1F;
  LUT6_L desc660(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[10:10]),.LO(pos_out_r_iv_i[10:10]));
defparam desc660.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc661(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[9:9]),.LO(pos_out_r_iv_i[9:9]));
defparam desc661.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc662(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[8:8]),.LO(pos_out_r_iv_i[8:8]));
defparam desc662.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc663(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[7:7]),.LO(pos_out_r_iv_i[7:7]));
defparam desc663.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc664(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[6:6]),.LO(pos_out_r_iv_i[6:6]));
defparam desc664.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc665(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[5:5]),.LO(pos_out_r_iv_i[5:5]));
defparam desc665.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc666(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[4:4]),.LO(pos_out_r_iv_i[4:4]));
defparam desc666.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc667(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[3:3]),.LO(pos_out_r_iv_i[3:3]));
defparam desc667.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc668(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[2:2]),.LO(pos_out_r_iv_i[2:2]));
defparam desc668.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc669(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(PATTERNDETECT_6),.I4(un5_rnd_sat_out_r_3),.I5(un2_rnd_out_r[1:1]),.LO(pos_out_r_iv_i[1:1]));
defparam desc669.INIT=64'hFFFF2F2F242F242F;
  LUT6_L desc670(.I0(mult2_out[23:23]),.I1(mult1_out[23:23]),.I2(pre_out_r[23:23]),.I3(un2_rnd_out_r[0:0]),.I4(PATTERNDETECT_6),.I5(un5_rnd_sat_out_r_3),.LO(pos_out_r_iv_i[0:0]));
defparam desc670.INIT=64'hFF24FF2F2F242F2F;
  XORCY un1_rnd_out_i_s_12(.LI(un1_rnd_out_i_axb_12),.CI(un1_rnd_out_i_cry_11),.O(un1_rnd_out_i_s_12_1));
  XORCY un1_rnd_out_i_s_11(.LI(un1_rnd_out_i_axb_11),.CI(un1_rnd_out_i_cry_10),.O(un1_rnd_out_i[10:10]));
  MUXCY_L un1_rnd_out_i_cry_11_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_10),.S(un1_rnd_out_i_axb_11),.LO(un1_rnd_out_i_cry_11));
  XORCY un1_rnd_out_i_s_10(.LI(un1_rnd_out_i_axb_10),.CI(un1_rnd_out_i_cry_9),.O(un1_rnd_out_i[9:9]));
  MUXCY_L un1_rnd_out_i_cry_10_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_9),.S(un1_rnd_out_i_axb_10),.LO(un1_rnd_out_i_cry_10));
  XORCY un1_rnd_out_i_s_9(.LI(un1_rnd_out_i_axb_9),.CI(un1_rnd_out_i_cry_8),.O(un1_rnd_out_i[8:8]));
  MUXCY_L un1_rnd_out_i_cry_9_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_8),.S(un1_rnd_out_i_axb_9),.LO(un1_rnd_out_i_cry_9));
  XORCY un1_rnd_out_i_s_8(.LI(un1_rnd_out_i_axb_8),.CI(un1_rnd_out_i_cry_7),.O(un1_rnd_out_i[7:7]));
  MUXCY_L un1_rnd_out_i_cry_8_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_7),.S(un1_rnd_out_i_axb_8),.LO(un1_rnd_out_i_cry_8));
  XORCY un1_rnd_out_i_s_7(.LI(un1_rnd_out_i_axb_7),.CI(un1_rnd_out_i_cry_6),.O(un1_rnd_out_i[6:6]));
  MUXCY_L un1_rnd_out_i_cry_7_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_6),.S(un1_rnd_out_i_axb_7),.LO(un1_rnd_out_i_cry_7));
  XORCY un1_rnd_out_i_s_6(.LI(un1_rnd_out_i_axb_6),.CI(un1_rnd_out_i_cry_5),.O(un1_rnd_out_i[5:5]));
  MUXCY_L un1_rnd_out_i_cry_6_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_5),.S(un1_rnd_out_i_axb_6),.LO(un1_rnd_out_i_cry_6));
  XORCY un1_rnd_out_i_s_5(.LI(un1_rnd_out_i_axb_5),.CI(un1_rnd_out_i_cry_4),.O(un1_rnd_out_i[4:4]));
  MUXCY_L un1_rnd_out_i_cry_5_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_4),.S(un1_rnd_out_i_axb_5),.LO(un1_rnd_out_i_cry_5));
  XORCY un1_rnd_out_i_s_4(.LI(un1_rnd_out_i_axb_4),.CI(un1_rnd_out_i_cry_3),.O(un1_rnd_out_i[3:3]));
  MUXCY_L un1_rnd_out_i_cry_4_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_3),.S(un1_rnd_out_i_axb_4),.LO(un1_rnd_out_i_cry_4));
  XORCY un1_rnd_out_i_s_3(.LI(un1_rnd_out_i_axb_3),.CI(un1_rnd_out_i_cry_2),.O(un1_rnd_out_i[2:2]));
  MUXCY_L un1_rnd_out_i_cry_3_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_2),.S(un1_rnd_out_i_axb_3),.LO(un1_rnd_out_i_cry_3));
  XORCY un1_rnd_out_i_s_2(.LI(un1_rnd_out_i_axb_2),.CI(un1_rnd_out_i_cry_1),.O(un1_rnd_out_i[1:1]));
  MUXCY_L un1_rnd_out_i_cry_2_cZ(.DI(GND),.CI(un1_rnd_out_i_cry_1),.S(un1_rnd_out_i_axb_2),.LO(un1_rnd_out_i_cry_2));
  XORCY un1_rnd_out_i_s_1(.LI(un1_rnd_out_i_axb_1),.CI(pre_out_i[7:7]),.O(un1_rnd_out_i[0:0]));
  MUXCY_L un1_rnd_out_i_cry_1_cZ(.DI(GND),.CI(pre_out_i[7:7]),.S(un1_rnd_out_i_axb_1),.LO(un1_rnd_out_i_cry_1));
  XORCY un2_rnd_out_r_s_12(.LI(un2_rnd_out_r_axb_12),.CI(un2_rnd_out_r_cry_11),.O(un2_rnd_out_r_s_12_1));
  XORCY un2_rnd_out_r_s_11(.LI(un2_rnd_out_r_axb_11),.CI(un2_rnd_out_r_cry_10),.O(un2_rnd_out_r[10:10]));
  MUXCY_L un2_rnd_out_r_cry_11_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_10),.S(un2_rnd_out_r_axb_11),.LO(un2_rnd_out_r_cry_11));
  XORCY un2_rnd_out_r_s_10(.LI(un2_rnd_out_r_axb_10),.CI(un2_rnd_out_r_cry_9),.O(un2_rnd_out_r[9:9]));
  MUXCY_L un2_rnd_out_r_cry_10_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_9),.S(un2_rnd_out_r_axb_10),.LO(un2_rnd_out_r_cry_10));
  XORCY un2_rnd_out_r_s_9(.LI(un2_rnd_out_r_axb_9),.CI(un2_rnd_out_r_cry_8),.O(un2_rnd_out_r[8:8]));
  MUXCY_L un2_rnd_out_r_cry_9_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_8),.S(un2_rnd_out_r_axb_9),.LO(un2_rnd_out_r_cry_9));
  XORCY un2_rnd_out_r_s_8(.LI(un2_rnd_out_r_axb_8),.CI(un2_rnd_out_r_cry_7),.O(un2_rnd_out_r[7:7]));
  MUXCY_L un2_rnd_out_r_cry_8_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_7),.S(un2_rnd_out_r_axb_8),.LO(un2_rnd_out_r_cry_8));
  XORCY un2_rnd_out_r_s_7(.LI(un2_rnd_out_r_axb_7),.CI(un2_rnd_out_r_cry_6),.O(un2_rnd_out_r[6:6]));
  MUXCY_L un2_rnd_out_r_cry_7_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_6),.S(un2_rnd_out_r_axb_7),.LO(un2_rnd_out_r_cry_7));
  XORCY un2_rnd_out_r_s_6(.LI(un2_rnd_out_r_axb_6),.CI(un2_rnd_out_r_cry_5),.O(un2_rnd_out_r[5:5]));
  MUXCY_L un2_rnd_out_r_cry_6_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_5),.S(un2_rnd_out_r_axb_6),.LO(un2_rnd_out_r_cry_6));
  XORCY un2_rnd_out_r_s_5(.LI(un2_rnd_out_r_axb_5),.CI(un2_rnd_out_r_cry_4),.O(un2_rnd_out_r[4:4]));
  MUXCY_L un2_rnd_out_r_cry_5_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_4),.S(un2_rnd_out_r_axb_5),.LO(un2_rnd_out_r_cry_5));
  XORCY un2_rnd_out_r_s_4(.LI(un2_rnd_out_r_axb_4),.CI(un2_rnd_out_r_cry_3),.O(un2_rnd_out_r[3:3]));
  MUXCY_L un2_rnd_out_r_cry_4_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_3),.S(un2_rnd_out_r_axb_4),.LO(un2_rnd_out_r_cry_4));
  XORCY un2_rnd_out_r_s_3(.LI(un2_rnd_out_r_axb_3),.CI(un2_rnd_out_r_cry_2),.O(un2_rnd_out_r[2:2]));
  MUXCY_L un2_rnd_out_r_cry_3_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_2),.S(un2_rnd_out_r_axb_3),.LO(un2_rnd_out_r_cry_3));
  XORCY un2_rnd_out_r_s_2(.LI(un2_rnd_out_r_axb_2),.CI(un2_rnd_out_r_cry_1),.O(un2_rnd_out_r[1:1]));
  MUXCY_L un2_rnd_out_r_cry_2_cZ(.DI(GND),.CI(un2_rnd_out_r_cry_1),.S(un2_rnd_out_r_axb_2),.LO(un2_rnd_out_r_cry_2));
  XORCY un2_rnd_out_r_s_1(.LI(un2_rnd_out_r_axb_1),.CI(pre_out_r[7:7]),.O(un2_rnd_out_r[0:0]));
  MUXCY_L un2_rnd_out_r_cry_1_cZ(.DI(GND),.CI(pre_out_r[7:7]),.S(un2_rnd_out_r_axb_1),.LO(un2_rnd_out_r_cry_1));
  FDS desc671(.Q(out_i_vec_mult_3[11:11]),.D(pos_out_i[11:11]),.C(clk),.S(un1_pos_out_i_2));
  FDR desc672(.Q(out_i_vec_mult_3[10:10]),.D(pos_out_i_iv_i[10:10]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc673(.Q(out_i_vec_mult_3[9:9]),.D(pos_out_i_iv_i[9:9]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc674(.Q(out_i_vec_mult_3[8:8]),.D(pos_out_i_iv_i[8:8]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc675(.Q(out_i_vec_mult_3[7:7]),.D(pos_out_i_iv_i[7:7]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc676(.Q(out_i_vec_mult_3[6:6]),.D(pos_out_i_iv_i[6:6]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc677(.Q(out_i_vec_mult_3[5:5]),.D(pos_out_i_iv_i[5:5]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc678(.Q(out_i_vec_mult_3[4:4]),.D(pos_out_i_iv_i[4:4]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc679(.Q(out_i_vec_mult_3[3:3]),.D(pos_out_i_iv_i[3:3]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc680(.Q(out_i_vec_mult_3[2:2]),.D(pos_out_i_iv_i[2:2]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc681(.Q(out_i_vec_mult_3[1:1]),.D(pos_out_i_iv_i[1:1]),.C(clk),.R(un1_pos_out_i_2));
  FDR desc682(.Q(out_i_vec_mult_3[0:0]),.D(pos_out_i_iv_i[0:0]),.C(clk),.R(un1_pos_out_i_2));
  FDS desc683(.Q(out_r_vec_mult_3[11:11]),.D(pos_out_r[11:11]),.C(clk),.S(un1_pos_out_r_2));
  FDR desc684(.Q(out_r_vec_mult_3[10:10]),.D(pos_out_r_iv_i[10:10]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc685(.Q(out_r_vec_mult_3[9:9]),.D(pos_out_r_iv_i[9:9]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc686(.Q(out_r_vec_mult_3[8:8]),.D(pos_out_r_iv_i[8:8]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc687(.Q(out_r_vec_mult_3[7:7]),.D(pos_out_r_iv_i[7:7]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc688(.Q(out_r_vec_mult_3[6:6]),.D(pos_out_r_iv_i[6:6]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc689(.Q(out_r_vec_mult_3[5:5]),.D(pos_out_r_iv_i[5:5]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc690(.Q(out_r_vec_mult_3[4:4]),.D(pos_out_r_iv_i[4:4]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc691(.Q(out_r_vec_mult_3[3:3]),.D(pos_out_r_iv_i[3:3]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc692(.Q(out_r_vec_mult_3[2:2]),.D(pos_out_r_iv_i[2:2]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc693(.Q(out_r_vec_mult_3[1:1]),.D(pos_out_r_iv_i[1:1]),.C(clk),.R(un1_pos_out_r_2));
  FDR desc694(.Q(out_r_vec_mult_3[0:0]),.D(pos_out_r_iv_i[0:0]),.C(clk),.R(un1_pos_out_r_2));
  mult_pipe_16_inj mult1(.mult1_out_23(mult1_out[23:23]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_28_0(P_uc_28_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  mult_pipe_17_inj mult2(.mult2_out_23(mult2_out[23:23]),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_18_inj mult3(.mult3_out_23(mult3_out[23:23]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk));
  mult_pipe_19_inj mult4(.mult4_out_23(mult4_out[23:23]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_31_0(P_uc_31_0[47:24]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  add_subZ2_4_inj sub(.pre_out_r(pre_out_r[23:7]),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult1_out_0(mult1_out_0[23:0]),.P_uc_28_0(P_uc_28_0[47:24]),.PATTERNDETECT_6(PATTERNDETECT_6),.clk(clk));
  add_subZ1_4_inj add(.pre_out_i(pre_out_i[23:7]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.mult4_out_0(mult4_out_0[23:0]),.P_uc_31_0(P_uc_31_0[47:24]),.PATTERNDETECT_5(PATTERNDETECT_5),.clk(clk));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module desc940_inj (un8_rnd_out_un0_P_9,un8_rnd_out_un0_P_10,un8_rnd_out_un0_P_11,un8_rnd_out_un0_P_12,un8_rnd_out_un0_P_13,un8_rnd_out_un0_P_14,un8_rnd_out_un0_P_15,un8_rnd_out_un0_P_16,un8_rnd_out_un0_P_17,un8_rnd_out_un0_P_18,un8_rnd_out_un0_P_19,mult1_out,mult2_out,pre_out_23,un2_output_3,PATTERNDETECT_15);
output un8_rnd_out_un0_P_9 ;
output un8_rnd_out_un0_P_10 ;
output un8_rnd_out_un0_P_11 ;
output un8_rnd_out_un0_P_12 ;
output un8_rnd_out_un0_P_13 ;
output un8_rnd_out_un0_P_14 ;
output un8_rnd_out_un0_P_15 ;
output un8_rnd_out_un0_P_16 ;
output un8_rnd_out_un0_P_17 ;
output un8_rnd_out_un0_P_18 ;
output un8_rnd_out_un0_P_19 ;
input [11:0] mult1_out ;
input [11:0] mult2_out ;
output pre_out_23 ;
output un2_output_3 ;
output PATTERNDETECT_15 ;
wire un8_rnd_out_un0_P_9 ;
wire un8_rnd_out_un0_P_10 ;
wire un8_rnd_out_un0_P_11 ;
wire un8_rnd_out_un0_P_12 ;
wire un8_rnd_out_un0_P_13 ;
wire un8_rnd_out_un0_P_14 ;
wire un8_rnd_out_un0_P_15 ;
wire un8_rnd_out_un0_P_16 ;
wire un8_rnd_out_un0_P_17 ;
wire un8_rnd_out_un0_P_18 ;
wire un8_rnd_out_un0_P_19 ;
wire pre_out_23 ;
wire un2_output_3 ;
wire PATTERNDETECT_15 ;
wire [22:0] pre_out ;
wire [29:0] ACOUT_11 ;
wire [17:0] BCOUT_11 ;
wire [3:0] CARRYOUT_11 ;
wire [8:0] un8_rnd_out_un0_P ;
wire [23:20] P_uc_1 ;
wire [47:24] P_uc_11 ;
wire [47:0] PCOUT_11 ;
wire [29:0] ACOUT_15 ;
wire [17:0] BCOUT_15 ;
wire [3:0] CARRYOUT_15 ;
wire [47:24] P_uc_15 ;
wire [47:0] PCOUT_15 ;
wire CARRYCASCOUT_11 ;
wire MULTSIGNOUT_11 ;
wire OVERFLOW_11 ;
wire PATTERNBDETECT_11 ;
wire PATTERNDETECT_11 ;
wire UNDERFLOW_11 ;
wire VCC ;
wire GND ;
wire CARRYCASCOUT_15 ;
wire MULTSIGNOUT_15 ;
wire OVERFLOW_15 ;
wire PATTERNBDETECT_15 ;
wire UNDERFLOW_15 ;
// instances
  LUT4 desc941(.I0(pre_out[19:19]),.I1(pre_out[20:20]),.I2(pre_out[21:21]),.I3(pre_out[22:22]),.O(un2_output_3));
defparam desc941.INIT=16'h0001;
  DSP48E1 desc942(.ACOUT(ACOUT_11[29:0]),.BCOUT(BCOUT_11[17:0]),.CARRYCASCOUT(CARRYCASCOUT_11),.CARRYOUT(CARRYOUT_11[3:0]),.MULTSIGNOUT(MULTSIGNOUT_11),.OVERFLOW(OVERFLOW_11),.P({P_uc_11[47:24],P_uc_1[23:20],un8_rnd_out_un0_P_19,un8_rnd_out_un0_P_18,un8_rnd_out_un0_P_17,un8_rnd_out_un0_P_16,un8_rnd_out_un0_P_15,un8_rnd_out_un0_P_14,un8_rnd_out_un0_P_13,un8_rnd_out_un0_P_12,un8_rnd_out_un0_P_11,un8_rnd_out_un0_P_10,un8_rnd_out_un0_P_9,un8_rnd_out_un0_P[8:0]}),.PATTERNBDETECT(PATTERNBDETECT_11),.PATTERNDETECT(PATTERNDETECT_11),.PCOUT(PCOUT_11[47:0]),.UNDERFLOW(UNDERFLOW_11),.A({mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,GND,GND,GND,GND,GND,GND,GND}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(GND),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,VCC,VCC,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc942.ACASCREG=0;
defparam desc942.ADREG=0;
defparam desc942.ALUMODEREG=0;
defparam desc942.AREG=0;
defparam desc942.AUTORESET_PATDET="NO_RESET";
defparam desc942.A_INPUT="DIRECT";
defparam desc942.BCASCREG=0;
defparam desc942.BREG=0;
defparam desc942.B_INPUT="DIRECT";
defparam desc942.CARRYINREG=0;
defparam desc942.CARRYINSELREG=0;
defparam desc942.CREG=0;
defparam desc942.DREG=0;
defparam desc942.INMODEREG=0;
defparam desc942.MREG=0;
defparam desc942.OPMODEREG=0;
defparam desc942.PREG=0;
defparam desc942.USE_DPORT="FALSE";
defparam desc942.USE_MULT="MULTIPLY";
defparam desc942.USE_SIMD="ONE48";
  DSP48E1 desc943(.ACOUT(ACOUT_15[29:0]),.BCOUT(BCOUT_15[17:0]),.CARRYCASCOUT(CARRYCASCOUT_15),.CARRYOUT(CARRYOUT_15[3:0]),.MULTSIGNOUT(MULTSIGNOUT_15),.OVERFLOW(OVERFLOW_15),.P({P_uc_15[47:24],pre_out_23,pre_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_15),.PATTERNDETECT(PATTERNDETECT_15),.PCOUT(PCOUT_15[47:0]),.UNDERFLOW(UNDERFLOW_15),.A({mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:11],mult1_out[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:11],mult2_out[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(GND),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc943.ACASCREG=0;
defparam desc943.ADREG=0;
defparam desc943.ALUMODEREG=0;
defparam desc943.AREG=0;
defparam desc943.AUTORESET_PATDET="NO_RESET";
defparam desc943.A_INPUT="DIRECT";
defparam desc943.BCASCREG=0;
defparam desc943.BREG=0;
defparam desc943.B_INPUT="DIRECT";
defparam desc943.CARRYINREG=0;
defparam desc943.CARRYINSELREG=0;
defparam desc943.CREG=1;
defparam desc943.DREG=0;
defparam desc943.INMODEREG=0;
defparam desc943.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc943.MREG=0;
defparam desc943.OPMODEREG=0;
defparam desc943.PATTERN=48'b111111111111111111111111111111111111111111111111;
defparam desc943.PREG=0;
defparam desc943.SEL_MASK="MASK";
defparam desc943.USE_DPORT="FALSE";
defparam desc943.USE_MULT="MULTIPLY";
defparam desc943.USE_PATTERN_DETECT="PATDET";
defparam desc943.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module inner_prod_inj (out_inner_prod_i,out_inner_prod_r,in_a_inner_prod_sel,single_out_r_AQ_7,single_out_r_AQ_0,single_out_r_AQ_1,single_out_r_AQ_4,single_out_r_AQ_2,in_b_inner_prod_sel,vec_in_r_AQ_mux_0_6,vec_in_r_AQ_mux_0_7,vec_in_r_AQ_mux_0_0,vec_in_r_AQ_mux_0_9,vec_in_r_AQ_mux_0_1,vec_in_r_AQ_mux_0_8,vec_in_r_AQ_mux_0_4,vec_in_r_AQ_mux_0_3,vec_in_r_AQ_mux_0_2,vec_in_r_AQ_mux_0_10,vec_in_i_AQ_mux_0_7,vec_in_i_AQ_mux_0_1,vec_in_i_AQ_mux_0_0,vec_in_i_AQ_mux_0_6,vec_in_i_AQ_mux_0_8,vec_in_i_AQ_mux_0_10,vec_in_i_AQ_mux_0_5,vec_in_i_AQ_mux_0_9,vec_in_i_AQ_mux_0_4,vec_in_i_AQ_mux_0_11,single_out_i_AQ_1,single_out_i_AQ_0,single_out_i_AQ_8,single_out_i_AQ_10,single_out_i_AQ_9,single_out_i_AQ_4,single_out_i_AQ_11,output_iv,single_out_r_AQ2_4,single_out_r_AQ2_0,single_out_r_AQ2_1,single_out_r_AQ2_6,output_iv_0_4,output_iv_0_7,output_iv_0_0,output_iv_0_9,output_iv_0_1,output_iv_0_6,output_iv_0_3,output_iv_0_2,output_iv_0_8,out_r_vec_sub_0,out_i_vec_sub_0,single_out_i_AQ2_0,single_out_i_AQ2_5,single_out_i_AQ2_4,single_out_i_AQ2_1,single_out_i_AQ2_11,start_inner_prod,red_mat_reg,clk,rst,done_inner_prod,N_623,N_568,N_622,N_507,N_549,N_505,N_597,N_567,N_596,N_628,N_637,N_566,N_506,N_585,N_584,N_612,N_583,N_595,N_508,N_501,N_605,N_624,N_607,N_552,N_555,N_586,N_645,N_641,N_582,N_606,N_632,N_500,N_571,p_desc318_p_O_FDC,p_desc319_p_O_FDC,p_desc320_p_O_FDC,p_desc321_p_O_FDC,p_desc322_p_O_FDC,p_in_reg_enable_fsm_Z_p_O_FDC,p_done_Z_p_O_FDC,p_acc_enable_Z_p_O_FDC,p_desc325_p_O_FDC,p_desc326_p_O_FDC,p_desc327_p_O_FDC,p_desc328_p_O_FDC,p_desc329_p_O_FDC,p_desc330_p_O_FDC,p_desc331_p_O_FDC,p_desc332_p_O_FDC,p_desc333_p_O_FDC,p_desc334_p_O_FDC,p_desc335_p_O_FDC,p_desc336_p_O_FDC,p_desc337_p_O_FDC,p_desc338_p_O_FDC,p_desc339_p_O_FDC,p_desc340_p_O_FDC,p_desc341_p_O_FDC,p_desc342_p_O_FDC,p_desc343_p_O_FDC,p_desc344_p_O_FDC,p_desc345_p_O_FDC,p_desc346_p_O_FDC,p_desc347_p_O_FDC,p_desc348_p_O_FDC,p_desc349_p_O_FDC,p_desc350_p_O_FDC,p_desc375_p_O_FDC,p_desc376_p_O_FDC,p_desc377_p_O_FDC,p_desc378_p_O_FDC,p_desc379_p_O_FDC,p_desc380_p_O_FDC,p_desc381_p_O_FDC,p_desc382_p_O_FDC,p_desc383_p_O_FDC,p_desc384_p_O_FDC,p_desc385_p_O_FDC,p_desc386_p_O_FDC,p_desc387_p_O_FDC,p_desc388_p_O_FDC,p_desc389_p_O_FDC,p_desc390_p_O_FDC,p_desc391_p_O_FDC,p_desc392_p_O_FDC,p_desc393_p_O_FDC,p_desc394_p_O_FDC,p_desc395_p_O_FDC,p_desc396_p_O_FDC,p_desc397_p_O_FDC,p_desc398_p_O_FDC,p_acc_clear_Z_p_O_FDP,p_desc324_p_O_FDCE,p_desc351_p_O_FDCE,p_desc352_p_O_FDCE,p_desc353_p_O_FDCE,p_desc354_p_O_FDCE,p_desc355_p_O_FDCE,p_desc356_p_O_FDCE,p_desc357_p_O_FDCE,p_desc358_p_O_FDCE,p_desc359_p_O_FDCE,p_desc360_p_O_FDCE,p_desc361_p_O_FDCE,p_desc362_p_O_FDCE,p_desc363_p_O_FDCE,p_desc364_p_O_FDCE,p_desc365_p_O_FDCE,p_desc366_p_O_FDCE,p_desc367_p_O_FDCE,p_desc368_p_O_FDCE,p_desc369_p_O_FDCE,p_desc370_p_O_FDCE,p_desc371_p_O_FDCE,p_desc372_p_O_FDCE,p_desc373_p_O_FDCE,p_desc374_p_O_FDCE);
output [11:0] out_inner_prod_i ;
output [11:0] out_inner_prod_r ;
input in_a_inner_prod_sel ;
input single_out_r_AQ_7 ;
input single_out_r_AQ_0 ;
input single_out_r_AQ_1 ;
input single_out_r_AQ_4 ;
input single_out_r_AQ_2 ;
input in_b_inner_prod_sel ;
input vec_in_r_AQ_mux_0_6 ;
input vec_in_r_AQ_mux_0_7 ;
input vec_in_r_AQ_mux_0_0 ;
input vec_in_r_AQ_mux_0_9 ;
input vec_in_r_AQ_mux_0_1 ;
input vec_in_r_AQ_mux_0_8 ;
input vec_in_r_AQ_mux_0_4 ;
input vec_in_r_AQ_mux_0_3 ;
input vec_in_r_AQ_mux_0_2 ;
input vec_in_r_AQ_mux_0_10 ;
input vec_in_i_AQ_mux_0_7 ;
input vec_in_i_AQ_mux_0_1 ;
input vec_in_i_AQ_mux_0_0 ;
input vec_in_i_AQ_mux_0_6 ;
input vec_in_i_AQ_mux_0_8 ;
input vec_in_i_AQ_mux_0_10 ;
input vec_in_i_AQ_mux_0_5 ;
input vec_in_i_AQ_mux_0_9 ;
input vec_in_i_AQ_mux_0_4 ;
input vec_in_i_AQ_mux_0_11 ;
input single_out_i_AQ_1 ;
input single_out_i_AQ_0 ;
input single_out_i_AQ_8 ;
input single_out_i_AQ_10 ;
input single_out_i_AQ_9 ;
input single_out_i_AQ_4 ;
input single_out_i_AQ_11 ;
input [10:0] output_iv ;
input single_out_r_AQ2_4 ;
input single_out_r_AQ2_0 ;
input single_out_r_AQ2_1 ;
input single_out_r_AQ2_6 ;
input output_iv_0_4 ;
input output_iv_0_7 ;
input output_iv_0_0 ;
input output_iv_0_9 ;
input output_iv_0_1 ;
input output_iv_0_6 ;
input output_iv_0_3 ;
input output_iv_0_2 ;
input output_iv_0_8 ;
input [11:11] out_r_vec_sub_0 ;
input [11:11] out_i_vec_sub_0 ;
input single_out_i_AQ2_0 ;
input single_out_i_AQ2_5 ;
input single_out_i_AQ2_4 ;
input single_out_i_AQ2_1 ;
input single_out_i_AQ2_11 ;
input start_inner_prod ;
input red_mat_reg ;
input clk ;
input rst ;
output done_inner_prod ;
input N_623 ;
input N_568 ;
input N_622 ;
input N_507 ;
input N_549 ;
input N_505 ;
input N_597 ;
input N_567 ;
input N_596 ;
input N_628 ;
input N_637 ;
input N_566 ;
input N_506 ;
input N_585 ;
input N_584 ;
input N_612 ;
input N_583 ;
input N_595 ;
input N_508 ;
input N_501 ;
input N_605 ;
input N_624 ;
input N_607 ;
input N_552 ;
input N_555 ;
input N_586 ;
input N_645 ;
input N_641 ;
input N_582 ;
input N_606 ;
input N_632 ;
input N_500 ;
input N_571 ;
wire single_out_r_AQ_7 ;
wire single_out_r_AQ_0 ;
wire single_out_r_AQ_1 ;
wire single_out_r_AQ_4 ;
wire single_out_r_AQ_2 ;
wire vec_in_r_AQ_mux_0_6 ;
wire vec_in_r_AQ_mux_0_7 ;
wire vec_in_r_AQ_mux_0_0 ;
wire vec_in_r_AQ_mux_0_9 ;
wire vec_in_r_AQ_mux_0_1 ;
wire vec_in_r_AQ_mux_0_8 ;
wire vec_in_r_AQ_mux_0_4 ;
wire vec_in_r_AQ_mux_0_3 ;
wire vec_in_r_AQ_mux_0_2 ;
wire vec_in_r_AQ_mux_0_10 ;
wire vec_in_i_AQ_mux_0_7 ;
wire vec_in_i_AQ_mux_0_1 ;
wire vec_in_i_AQ_mux_0_0 ;
wire vec_in_i_AQ_mux_0_6 ;
wire vec_in_i_AQ_mux_0_8 ;
wire vec_in_i_AQ_mux_0_10 ;
wire vec_in_i_AQ_mux_0_5 ;
wire vec_in_i_AQ_mux_0_9 ;
wire vec_in_i_AQ_mux_0_4 ;
wire vec_in_i_AQ_mux_0_11 ;
wire single_out_i_AQ_1 ;
wire single_out_i_AQ_0 ;
wire single_out_i_AQ_8 ;
wire single_out_i_AQ_10 ;
wire single_out_i_AQ_9 ;
wire single_out_i_AQ_4 ;
wire single_out_i_AQ_11 ;
wire single_out_r_AQ2_4 ;
wire single_out_r_AQ2_0 ;
wire single_out_r_AQ2_1 ;
wire single_out_r_AQ2_6 ;
wire output_iv_0_4 ;
wire output_iv_0_7 ;
wire output_iv_0_0 ;
wire output_iv_0_9 ;
wire output_iv_0_1 ;
wire output_iv_0_6 ;
wire output_iv_0_3 ;
wire output_iv_0_2 ;
wire output_iv_0_8 ;
wire single_out_i_AQ2_0 ;
wire single_out_i_AQ2_5 ;
wire single_out_i_AQ2_4 ;
wire single_out_i_AQ2_1 ;
wire single_out_i_AQ2_11 ;
wire start_inner_prod ;
wire red_mat_reg ;
wire clk ;
wire rst ;
wire done_inner_prod ;
wire N_623 ;
wire N_568 ;
wire N_622 ;
wire N_507 ;
wire N_549 ;
wire N_505 ;
wire N_597 ;
wire N_567 ;
wire N_596 ;
wire N_628 ;
wire N_637 ;
wire N_566 ;
wire N_506 ;
wire N_585 ;
wire N_584 ;
wire N_612 ;
wire N_583 ;
wire N_595 ;
wire N_508 ;
wire N_501 ;
wire N_605 ;
wire N_624 ;
wire N_607 ;
wire N_552 ;
wire N_555 ;
wire N_586 ;
wire N_645 ;
wire N_641 ;
wire N_582 ;
wire N_606 ;
wire N_632 ;
wire N_500 ;
wire N_571 ;
wire [11:0] mult_out_i ;
wire [10:1] un2_pre_out ;
wire [11:0] acc_i_2 ;
wire [2:0] pipe_counter ;
wire [1:0] state ;
wire [2:0] in_counter ;
wire [2:1] pipe_counter_4_0_a2 ;
wire state_i_0 ;
wire [11:0] in_a_i_reg ;
wire [11:0] in_a_i_reg_2 ;
wire [11:0] in_a_r_reg ;
wire [8:1] in_a_r_reg_3 ;
wire [1:0] state_ns ;
wire [11:0] in_b_i_reg ;
wire [11:0] in_b_i_reg_2 ;
wire [11:0] in_b_r_reg ;
wire [11:1] in_b_r_reg_2 ;
wire [11:0] mult_out_r ;
wire [10:1] un2_pre_out_0 ;
wire acc_clear ;
wire un2_pre_out_s_11_0 ;
wire VCC ;
wire acc_enable ;
wire un1_state_4_0_0_lut6_2_O6 ;
wire acc_enable_0 ;
wire in_reg_enable_fsm_0_sqmuxa ;
wire un1_state_8_0_0_a2_lut6_2_O5 ;
wire un7_acc_enable_lut6_2_O6 ;
wire acc_clear_0 ;
wire in_counter_5_43_i_i_a2 ;
wire N_113_i_0 ;
wire in_reg_enable_fsm ;
wire in_reg_enable_fsm_0 ;
wire done ;
wire N_516_i_0 ;
wire N_518_i ;
wire N_519_i_0 ;
wire N_520_i ;
wire N_523_i ;
wire N_193_i ;
wire N_524_i ;
wire N_183_i ;
wire N_195_i ;
wire N_191_i ;
wire N_26_i ;
wire N_24_i ;
wire N_22_i ;
wire N_20_i ;
wire N_18_i ;
wire N_16_i ;
wire N_14_i ;
wire N_12_i ;
wire N_10_i ;
wire N_8_i ;
wire N_6_i ;
wire N_4_i ;
wire N_521_i ;
wire N_517_i_0 ;
wire N_522_i ;
wire N_185_i ;
wire un2_pre_out_s_11 ;
wire N_27 ;
wire N_26 ;
wire N_25 ;
wire GND ;
input p_desc318_p_O_FDC ;
input p_desc319_p_O_FDC ;
input p_desc320_p_O_FDC ;
input p_desc321_p_O_FDC ;
input p_desc322_p_O_FDC ;
input p_in_reg_enable_fsm_Z_p_O_FDC ;
input p_done_Z_p_O_FDC ;
input p_acc_enable_Z_p_O_FDC ;
input p_desc325_p_O_FDC ;
input p_desc326_p_O_FDC ;
input p_desc327_p_O_FDC ;
input p_desc328_p_O_FDC ;
input p_desc329_p_O_FDC ;
input p_desc330_p_O_FDC ;
input p_desc331_p_O_FDC ;
input p_desc332_p_O_FDC ;
input p_desc333_p_O_FDC ;
input p_desc334_p_O_FDC ;
input p_desc335_p_O_FDC ;
input p_desc336_p_O_FDC ;
input p_desc337_p_O_FDC ;
input p_desc338_p_O_FDC ;
input p_desc339_p_O_FDC ;
input p_desc340_p_O_FDC ;
input p_desc341_p_O_FDC ;
input p_desc342_p_O_FDC ;
input p_desc343_p_O_FDC ;
input p_desc344_p_O_FDC ;
input p_desc345_p_O_FDC ;
input p_desc346_p_O_FDC ;
input p_desc347_p_O_FDC ;
input p_desc348_p_O_FDC ;
input p_desc349_p_O_FDC ;
input p_desc350_p_O_FDC ;
input p_desc375_p_O_FDC ;
input p_desc376_p_O_FDC ;
input p_desc377_p_O_FDC ;
input p_desc378_p_O_FDC ;
input p_desc379_p_O_FDC ;
input p_desc380_p_O_FDC ;
input p_desc381_p_O_FDC ;
input p_desc382_p_O_FDC ;
input p_desc383_p_O_FDC ;
input p_desc384_p_O_FDC ;
input p_desc385_p_O_FDC ;
input p_desc386_p_O_FDC ;
input p_desc387_p_O_FDC ;
input p_desc388_p_O_FDC ;
input p_desc389_p_O_FDC ;
input p_desc390_p_O_FDC ;
input p_desc391_p_O_FDC ;
input p_desc392_p_O_FDC ;
input p_desc393_p_O_FDC ;
input p_desc394_p_O_FDC ;
input p_desc395_p_O_FDC ;
input p_desc396_p_O_FDC ;
input p_desc397_p_O_FDC ;
input p_desc398_p_O_FDC ;
input p_acc_clear_Z_p_O_FDP ;
input p_desc324_p_O_FDCE ;
input p_desc351_p_O_FDCE ;
input p_desc352_p_O_FDCE ;
input p_desc353_p_O_FDCE ;
input p_desc354_p_O_FDCE ;
input p_desc355_p_O_FDCE ;
input p_desc356_p_O_FDCE ;
input p_desc357_p_O_FDCE ;
input p_desc358_p_O_FDCE ;
input p_desc359_p_O_FDCE ;
input p_desc360_p_O_FDCE ;
input p_desc361_p_O_FDCE ;
input p_desc362_p_O_FDCE ;
input p_desc363_p_O_FDCE ;
input p_desc364_p_O_FDCE ;
input p_desc365_p_O_FDCE ;
input p_desc366_p_O_FDCE ;
input p_desc367_p_O_FDCE ;
input p_desc368_p_O_FDCE ;
input p_desc369_p_O_FDCE ;
input p_desc370_p_O_FDCE ;
input p_desc371_p_O_FDCE ;
input p_desc372_p_O_FDCE ;
input p_desc373_p_O_FDCE ;
input p_desc374_p_O_FDCE ;
// instances
  p_O_FDC desc318(.Q(in_counter[2:2]),.D(in_counter_5_43_i_i_a2),.C(clk),.CLR(rst),.E(p_desc318_p_O_FDC));
  p_O_FDC desc319(.Q(in_counter[1:1]),.D(N_113_i_0),.C(clk),.CLR(rst),.E(p_desc319_p_O_FDC));
  p_O_FDC desc320(.Q(in_counter[0:0]),.D(state_i_0),.C(clk),.CLR(rst),.E(p_desc320_p_O_FDC));
  p_O_FDC desc321(.Q(pipe_counter[2:2]),.D(pipe_counter_4_0_a2[2:2]),.C(clk),.CLR(rst),.E(p_desc321_p_O_FDC));
  p_O_FDC desc322(.Q(pipe_counter[1:1]),.D(pipe_counter_4_0_a2[1:1]),.C(clk),.CLR(rst),.E(p_desc322_p_O_FDC));
  LUT4 desc323(.I0(in_counter[0:0]),.I1(state[0:0]),.I2(in_counter[1:1]),.I3(un1_state_4_0_0_lut6_2_O6),.O(N_113_i_0));
defparam desc323.INIT=16'h88F0;
  p_O_FDCE desc324(.Q(pipe_counter[0:0]),.D(in_reg_enable_fsm_0_sqmuxa),.C(clk),.CLR(rst),.CE(un1_state_8_0_0_a2_lut6_2_O5),.E(p_desc324_p_O_FDCE));
  p_O_FDC in_reg_enable_fsm_Z(.Q(in_reg_enable_fsm),.D(in_reg_enable_fsm_0),.C(clk),.CLR(rst),.E(p_in_reg_enable_fsm_Z_p_O_FDC));
  p_O_FDC done_Z(.Q(done_inner_prod),.D(done),.C(clk),.CLR(rst),.E(p_done_Z_p_O_FDC));
  p_O_FDC acc_enable_Z(.Q(acc_enable),.D(acc_enable_0),.C(clk),.CLR(rst),.E(p_acc_enable_Z_p_O_FDC));
  p_O_FDP acc_clear_Z(.Q(acc_clear),.D(acc_clear_0),.C(clk),.PRE(rst),.E(p_acc_clear_Z_p_O_FDP));
  p_O_FDC desc325(.Q(in_a_i_reg[0:0]),.D(in_a_i_reg_2[0:0]),.C(clk),.CLR(rst),.E(p_desc325_p_O_FDC));
  p_O_FDC desc326(.Q(in_a_i_reg[1:1]),.D(in_a_i_reg_2[1:1]),.C(clk),.CLR(rst),.E(p_desc326_p_O_FDC));
  p_O_FDC desc327(.Q(in_a_i_reg[2:2]),.D(N_516_i_0),.C(clk),.CLR(rst),.E(p_desc327_p_O_FDC));
  p_O_FDC desc328(.Q(in_a_i_reg[3:3]),.D(N_518_i),.C(clk),.CLR(rst),.E(p_desc328_p_O_FDC));
  p_O_FDC desc329(.Q(in_a_i_reg[4:4]),.D(in_a_i_reg_2[4:4]),.C(clk),.CLR(rst),.E(p_desc329_p_O_FDC));
  p_O_FDC desc330(.Q(in_a_i_reg[5:5]),.D(in_a_i_reg_2[5:5]),.C(clk),.CLR(rst),.E(p_desc330_p_O_FDC));
  p_O_FDC desc331(.Q(in_a_i_reg[6:6]),.D(N_519_i_0),.C(clk),.CLR(rst),.E(p_desc331_p_O_FDC));
  p_O_FDC desc332(.Q(in_a_i_reg[7:7]),.D(N_520_i),.C(clk),.CLR(rst),.E(p_desc332_p_O_FDC));
  p_O_FDC desc333(.Q(in_a_i_reg[8:8]),.D(in_a_i_reg_2[8:8]),.C(clk),.CLR(rst),.E(p_desc333_p_O_FDC));
  p_O_FDC desc334(.Q(in_a_i_reg[9:9]),.D(in_a_i_reg_2[9:9]),.C(clk),.CLR(rst),.E(p_desc334_p_O_FDC));
  p_O_FDC desc335(.Q(in_a_i_reg[10:10]),.D(in_a_i_reg_2[10:10]),.C(clk),.CLR(rst),.E(p_desc335_p_O_FDC));
  p_O_FDC desc336(.Q(in_a_i_reg[11:11]),.D(in_a_i_reg_2[11:11]),.C(clk),.CLR(rst),.E(p_desc336_p_O_FDC));
  p_O_FDC desc337(.Q(in_a_r_reg[3:3]),.D(in_a_r_reg_3[3:3]),.C(clk),.CLR(rst),.E(p_desc337_p_O_FDC));
  p_O_FDC desc338(.Q(in_a_r_reg[4:4]),.D(in_a_r_reg_3[4:4]),.C(clk),.CLR(rst),.E(p_desc338_p_O_FDC));
  p_O_FDC desc339(.Q(in_a_r_reg[5:5]),.D(in_a_r_reg_3[5:5]),.C(clk),.CLR(rst),.E(p_desc339_p_O_FDC));
  p_O_FDC desc340(.Q(in_a_r_reg[6:6]),.D(N_523_i),.C(clk),.CLR(rst),.E(p_desc340_p_O_FDC));
  p_O_FDC desc341(.Q(in_a_r_reg[7:7]),.D(N_193_i),.C(clk),.CLR(rst),.E(p_desc341_p_O_FDC));
  p_O_FDC desc342(.Q(in_a_r_reg[8:8]),.D(in_a_r_reg_3[8:8]),.C(clk),.CLR(rst),.E(p_desc342_p_O_FDC));
  p_O_FDC desc343(.Q(in_a_r_reg[9:9]),.D(N_524_i),.C(clk),.CLR(rst),.E(p_desc343_p_O_FDC));
  p_O_FDC desc344(.Q(in_a_r_reg[10:10]),.D(N_183_i),.C(clk),.CLR(rst),.E(p_desc344_p_O_FDC));
  p_O_FDC desc345(.Q(in_a_r_reg[11:11]),.D(N_195_i),.C(clk),.CLR(rst),.E(p_desc345_p_O_FDC));
  p_O_FDC desc346(.Q(in_a_r_reg[0:0]),.D(N_191_i),.C(clk),.CLR(rst),.E(p_desc346_p_O_FDC));
  p_O_FDC desc347(.Q(in_a_r_reg[1:1]),.D(in_a_r_reg_3[1:1]),.C(clk),.CLR(rst),.E(p_desc347_p_O_FDC));
  p_O_FDC desc348(.Q(in_a_r_reg[2:2]),.D(in_a_r_reg_3[2:2]),.C(clk),.CLR(rst),.E(p_desc348_p_O_FDC));
  p_O_FDC desc349(.Q(state[0:0]),.D(state_ns[0:0]),.C(clk),.CLR(rst),.E(p_desc349_p_O_FDC));
  p_O_FDC desc350(.Q(state[1:1]),.D(state_ns[1:1]),.C(clk),.CLR(rst),.E(p_desc350_p_O_FDC));
  p_O_FDCE desc351(.Q(out_inner_prod_i[11:11]),.D(acc_i_2[11:11]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc351_p_O_FDCE));
  p_O_FDCE desc352(.Q(out_inner_prod_i[10:10]),.D(acc_i_2[10:10]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc352_p_O_FDCE));
  p_O_FDCE desc353(.Q(out_inner_prod_i[9:9]),.D(acc_i_2[9:9]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc353_p_O_FDCE));
  p_O_FDCE desc354(.Q(out_inner_prod_i[8:8]),.D(acc_i_2[8:8]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc354_p_O_FDCE));
  p_O_FDCE desc355(.Q(out_inner_prod_i[7:7]),.D(acc_i_2[7:7]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc355_p_O_FDCE));
  p_O_FDCE desc356(.Q(out_inner_prod_i[6:6]),.D(acc_i_2[6:6]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc356_p_O_FDCE));
  p_O_FDCE desc357(.Q(out_inner_prod_i[5:5]),.D(acc_i_2[5:5]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc357_p_O_FDCE));
  p_O_FDCE desc358(.Q(out_inner_prod_i[4:4]),.D(acc_i_2[4:4]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc358_p_O_FDCE));
  p_O_FDCE desc359(.Q(out_inner_prod_i[3:3]),.D(acc_i_2[3:3]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc359_p_O_FDCE));
  p_O_FDCE desc360(.Q(out_inner_prod_i[2:2]),.D(acc_i_2[2:2]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc360_p_O_FDCE));
  p_O_FDCE desc361(.Q(out_inner_prod_i[1:1]),.D(acc_i_2[1:1]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc361_p_O_FDCE));
  p_O_FDCE desc362(.Q(out_inner_prod_i[0:0]),.D(acc_i_2[0:0]),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc362_p_O_FDCE));
  p_O_FDCE desc363(.Q(out_inner_prod_r[11:11]),.D(N_26_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc363_p_O_FDCE));
  p_O_FDCE desc364(.Q(out_inner_prod_r[10:10]),.D(N_24_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc364_p_O_FDCE));
  p_O_FDCE desc365(.Q(out_inner_prod_r[9:9]),.D(N_22_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc365_p_O_FDCE));
  p_O_FDCE desc366(.Q(out_inner_prod_r[8:8]),.D(N_20_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc366_p_O_FDCE));
  p_O_FDCE desc367(.Q(out_inner_prod_r[7:7]),.D(N_18_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc367_p_O_FDCE));
  p_O_FDCE desc368(.Q(out_inner_prod_r[6:6]),.D(N_16_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc368_p_O_FDCE));
  p_O_FDCE desc369(.Q(out_inner_prod_r[5:5]),.D(N_14_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc369_p_O_FDCE));
  p_O_FDCE desc370(.Q(out_inner_prod_r[4:4]),.D(N_12_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc370_p_O_FDCE));
  p_O_FDCE desc371(.Q(out_inner_prod_r[3:3]),.D(N_10_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc371_p_O_FDCE));
  p_O_FDCE desc372(.Q(out_inner_prod_r[2:2]),.D(N_8_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc372_p_O_FDCE));
  p_O_FDCE desc373(.Q(out_inner_prod_r[1:1]),.D(N_6_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc373_p_O_FDCE));
  p_O_FDCE desc374(.Q(out_inner_prod_r[0:0]),.D(N_4_i),.C(clk),.CLR(rst),.CE(un7_acc_enable_lut6_2_O6),.E(p_desc374_p_O_FDCE));
  p_O_FDC desc375(.Q(in_b_i_reg[11:11]),.D(in_b_i_reg_2[11:11]),.C(clk),.CLR(rst),.E(p_desc375_p_O_FDC));
  p_O_FDC desc376(.Q(in_b_i_reg[10:10]),.D(in_b_i_reg_2[10:10]),.C(clk),.CLR(rst),.E(p_desc376_p_O_FDC));
  p_O_FDC desc377(.Q(in_b_i_reg[9:9]),.D(in_b_i_reg_2[9:9]),.C(clk),.CLR(rst),.E(p_desc377_p_O_FDC));
  p_O_FDC desc378(.Q(in_b_i_reg[8:8]),.D(in_b_i_reg_2[8:8]),.C(clk),.CLR(rst),.E(p_desc378_p_O_FDC));
  p_O_FDC desc379(.Q(in_b_i_reg[7:7]),.D(in_b_i_reg_2[7:7]),.C(clk),.CLR(rst),.E(p_desc379_p_O_FDC));
  p_O_FDC desc380(.Q(in_b_i_reg[6:6]),.D(in_b_i_reg_2[6:6]),.C(clk),.CLR(rst),.E(p_desc380_p_O_FDC));
  p_O_FDC desc381(.Q(in_b_i_reg[5:5]),.D(in_b_i_reg_2[5:5]),.C(clk),.CLR(rst),.E(p_desc381_p_O_FDC));
  p_O_FDC desc382(.Q(in_b_i_reg[4:4]),.D(in_b_i_reg_2[4:4]),.C(clk),.CLR(rst),.E(p_desc382_p_O_FDC));
  p_O_FDC desc383(.Q(in_b_i_reg[3:3]),.D(N_521_i),.C(clk),.CLR(rst),.E(p_desc383_p_O_FDC));
  p_O_FDC desc384(.Q(in_b_i_reg[2:2]),.D(N_517_i_0),.C(clk),.CLR(rst),.E(p_desc384_p_O_FDC));
  p_O_FDC desc385(.Q(in_b_i_reg[1:1]),.D(in_b_i_reg_2[1:1]),.C(clk),.CLR(rst),.E(p_desc385_p_O_FDC));
  p_O_FDC desc386(.Q(in_b_i_reg[0:0]),.D(in_b_i_reg_2[0:0]),.C(clk),.CLR(rst),.E(p_desc386_p_O_FDC));
  p_O_FDC desc387(.Q(in_b_r_reg[11:11]),.D(in_b_r_reg_2[11:11]),.C(clk),.CLR(rst),.E(p_desc387_p_O_FDC));
  p_O_FDC desc388(.Q(in_b_r_reg[10:10]),.D(in_b_r_reg_2[10:10]),.C(clk),.CLR(rst),.E(p_desc388_p_O_FDC));
  p_O_FDC desc389(.Q(in_b_r_reg[9:9]),.D(in_b_r_reg_2[9:9]),.C(clk),.CLR(rst),.E(p_desc389_p_O_FDC));
  p_O_FDC desc390(.Q(in_b_r_reg[8:8]),.D(in_b_r_reg_2[8:8]),.C(clk),.CLR(rst),.E(p_desc390_p_O_FDC));
  p_O_FDC desc391(.Q(in_b_r_reg[7:7]),.D(in_b_r_reg_2[7:7]),.C(clk),.CLR(rst),.E(p_desc391_p_O_FDC));
  p_O_FDC desc392(.Q(in_b_r_reg[6:6]),.D(N_522_i),.C(clk),.CLR(rst),.E(p_desc392_p_O_FDC));
  p_O_FDC desc393(.Q(in_b_r_reg[5:5]),.D(in_b_r_reg_2[5:5]),.C(clk),.CLR(rst),.E(p_desc393_p_O_FDC));
  p_O_FDC desc394(.Q(in_b_r_reg[4:4]),.D(in_b_r_reg_2[4:4]),.C(clk),.CLR(rst),.E(p_desc394_p_O_FDC));
  p_O_FDC desc395(.Q(in_b_r_reg[3:3]),.D(in_b_r_reg_2[3:3]),.C(clk),.CLR(rst),.E(p_desc395_p_O_FDC));
  p_O_FDC desc396(.Q(in_b_r_reg[2:2]),.D(in_b_r_reg_2[2:2]),.C(clk),.CLR(rst),.E(p_desc396_p_O_FDC));
  p_O_FDC desc397(.Q(in_b_r_reg[1:1]),.D(in_b_r_reg_2[1:1]),.C(clk),.CLR(rst),.E(p_desc397_p_O_FDC));
  p_O_FDC desc398(.Q(in_b_r_reg[0:0]),.D(N_185_i),.C(clk),.CLR(rst),.E(p_desc398_p_O_FDC));
  LUT5_L desc399(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_623),.I4(vec_in_r_AQ_mux_0_6),.LO(N_193_i));
defparam desc399.INIT=32'hFC54A800;
  LUT5_L desc400(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_r_AQ_7),.I4(vec_in_r_AQ_mux_0_7),.LO(in_a_r_reg_3[8:8]));
defparam desc400.INIT=32'hFC54A800;
  LUT5_L desc401(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_r_AQ_0),.I4(vec_in_r_AQ_mux_0_0),.LO(in_a_r_reg_3[1:1]));
defparam desc401.INIT=32'hFC54A800;
  LUT5_L desc402(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_568),.I4(vec_in_i_AQ_mux_0_7),.LO(N_520_i));
defparam desc402.INIT=32'hFC54A800;
  LUT5_L desc403(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_622),.I4(N_507),.LO(N_191_i));
defparam desc403.INIT=32'hFC54A800;
  LUT5_L desc404(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_1),.I4(vec_in_i_AQ_mux_0_1),.LO(in_a_i_reg_2[1:1]));
defparam desc404.INIT=32'hFC54A800;
  LUT5_L desc405(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_0),.I4(vec_in_i_AQ_mux_0_0),.LO(in_a_i_reg_2[0:0]));
defparam desc405.INIT=32'hFC54A800;
  LUT5_L desc406(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_549),.I4(N_505),.LO(N_516_i_0));
defparam desc406.INIT=32'hFC54A800;
  LUT5_L desc407(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_597),.I4(vec_in_r_AQ_mux_0_9),.LO(N_183_i));
defparam desc407.INIT=32'hFC54A800;
  LUT5_L desc408(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_567),.I4(vec_in_i_AQ_mux_0_6),.LO(N_519_i_0));
defparam desc408.INIT=32'hFC54A800;
  LUT5_L desc409(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_r_AQ_1),.I4(vec_in_r_AQ_mux_0_1),.LO(in_a_r_reg_3[2:2]));
defparam desc409.INIT=32'hFC54A800;
  LUT5_L desc410(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_596),.I4(vec_in_r_AQ_mux_0_8),.LO(N_524_i));
defparam desc410.INIT=32'hFC54A800;
  LUT5_L desc411(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_8),.I4(vec_in_i_AQ_mux_0_8),.LO(in_a_i_reg_2[8:8]));
defparam desc411.INIT=32'hFC54A800;
  LUT5_L desc412(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_10),.I4(vec_in_i_AQ_mux_0_10),.LO(in_a_i_reg_2[10:10]));
defparam desc412.INIT=32'hFC54A800;
  LUT5_L desc413(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_628),.I4(vec_in_i_AQ_mux_0_5),.LO(in_a_i_reg_2[5:5]));
defparam desc413.INIT=32'hFC54A800;
  LUT5_L desc414(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_r_AQ_4),.I4(vec_in_r_AQ_mux_0_4),.LO(in_a_r_reg_3[5:5]));
defparam desc414.INIT=32'hFC54A800;
  LUT5_L desc415(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_637),.I4(vec_in_r_AQ_mux_0_3),.LO(in_a_r_reg_3[4:4]));
defparam desc415.INIT=32'hFC54A800;
  LUT5_L desc416(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_9),.I4(vec_in_i_AQ_mux_0_9),.LO(in_a_i_reg_2[9:9]));
defparam desc416.INIT=32'hFC54A800;
  LUT5_L desc417(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_i_AQ_4),.I4(vec_in_i_AQ_mux_0_4),.LO(in_a_i_reg_2[4:4]));
defparam desc417.INIT=32'hFC54A800;
  LUT5_L desc418(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(single_out_r_AQ_2),.I4(vec_in_r_AQ_mux_0_2),.LO(in_a_r_reg_3[3:3]));
defparam desc418.INIT=32'hFC54A800;
  LUT5_L desc419(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_566),.I4(N_506),.LO(N_518_i));
defparam desc419.INIT=32'hFC54A800;
  LUT5_L desc420(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[9:9]),.I4(N_585),.LO(in_b_i_reg_2[9:9]));
defparam desc420.INIT=32'hA8FC0054;
  LUT5_L desc421(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[5:5]),.I4(single_out_r_AQ2_4),.LO(in_b_r_reg_2[5:5]));
defparam desc421.INIT=32'hA8FC0054;
  LUT5_L desc422(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[7:7]),.I4(N_584),.LO(in_b_i_reg_2[7:7]));
defparam desc422.INIT=32'hA8FC0054;
  LUT5_L desc423(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[8:8]),.I4(N_612),.LO(in_b_i_reg_2[8:8]));
defparam desc423.INIT=32'hA8FC0054;
  LUT5_L desc424(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[6:6]),.I4(N_583),.LO(in_b_i_reg_2[6:6]));
defparam desc424.INIT=32'hA8FC0054;
  LUT5_L desc425(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_595),.I4(N_508),.LO(N_523_i));
defparam desc425.INIT=32'hFC54A800;
  LUT5_L desc426(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[1:1]),.I4(single_out_r_AQ2_0),.LO(in_b_r_reg_2[1:1]));
defparam desc426.INIT=32'hA8FC0054;
  LUT5_L desc427(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[0:0]),.I4(single_out_i_AQ2_0),.LO(in_b_i_reg_2[0:0]));
defparam desc427.INIT=32'hA8FC0054;
  LUT5_L desc428(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_4),.I4(single_out_i_AQ2_5),.LO(in_b_i_reg_2[5:5]));
defparam desc428.INIT=32'hA8FC0054;
  LUT5_L desc429(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_501),.I4(N_605),.LO(N_185_i));
defparam desc429.INIT=32'hA8FC0054;
  LUT5_L desc430(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(vec_in_r_AQ_mux_0_10),.I4(N_624),.LO(N_195_i));
defparam desc430.INIT=32'hFCA85400;
  LUT5_L desc431(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[4:4]),.I4(single_out_i_AQ2_4),.LO(in_b_i_reg_2[4:4]));
defparam desc431.INIT=32'hA8FC0054;
  LUT5_L desc432(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[10:10]),.I4(N_607),.LO(in_b_r_reg_2[10:10]));
defparam desc432.INIT=32'hA8FC0054;
  LUT5_L desc433(.I0(in_a_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(vec_in_i_AQ_mux_0_11),.I4(single_out_i_AQ_11),.LO(in_a_i_reg_2[11:11]));
defparam desc433.INIT=32'hFCA85400;
  LUT5_L desc434(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_7),.I4(N_552),.LO(in_b_r_reg_2[8:8]));
defparam desc434.INIT=32'hA8FC0054;
  LUT5_L desc435(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[2:2]),.I4(N_555),.LO(N_517_i_0));
defparam desc435.INIT=32'hA8FC0054;
  LUT5_L desc436(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_0),.I4(single_out_i_AQ2_1),.LO(in_b_i_reg_2[1:1]));
defparam desc436.INIT=32'hA8FC0054;
  LUT5_L desc437(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_9),.I4(N_586),.LO(in_b_i_reg_2[10:10]));
defparam desc437.INIT=32'hA8FC0054;
  LUT5_L desc438(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv[3:3]),.I4(N_645),.LO(in_b_r_reg_2[3:3]));
defparam desc438.INIT=32'hA8FC0054;
  LUT5_L desc439(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_1),.I4(single_out_r_AQ2_1),.LO(in_b_r_reg_2[2:2]));
defparam desc439.INIT=32'hA8FC0054;
  LUT5_L desc440(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_6),.I4(single_out_r_AQ2_6),.LO(in_b_r_reg_2[7:7]));
defparam desc440.INIT=32'hA8FC0054;
  LUT5_L desc441(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_3),.I4(N_641),.LO(in_b_r_reg_2[4:4]));
defparam desc441.INIT=32'hA8FC0054;
  LUT5_L desc442(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_2),.I4(N_582),.LO(N_521_i));
defparam desc442.INIT=32'hA8FC0054;
  LUT5_L desc443(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(output_iv_0_8),.I4(N_606),.LO(in_b_r_reg_2[9:9]));
defparam desc443.INIT=32'hA8FC0054;
  LUT5_L desc444(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(out_r_vec_sub_0[11:11]),.I4(N_632),.LO(in_b_r_reg_2[11:11]));
defparam desc444.INIT=32'hFCA85400;
  LUT5_L desc445(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(out_i_vec_sub_0[11:11]),.I4(single_out_i_AQ2_11),.LO(in_b_i_reg_2[11:11]));
defparam desc445.INIT=32'hFCA85400;
  LUT5_L desc446(.I0(in_b_inner_prod_sel),.I1(in_reg_enable_fsm),.I2(start_inner_prod),.I3(N_500),.I4(N_571),.LO(N_522_i));
defparam desc446.INIT=32'hA8FC0054;
  LUT5_L desc447(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[7:7]),.I4(un2_pre_out_s_11),.LO(N_18_i));
defparam desc447.INIT=32'h33011300;
  LUT5_L desc448(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[6:6]),.I4(un2_pre_out_s_11),.LO(N_16_i));
defparam desc448.INIT=32'h33011300;
  LUT5_L desc449(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[5:5]),.I4(un2_pre_out_s_11),.LO(N_14_i));
defparam desc449.INIT=32'h33011300;
  LUT5_L desc450(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[4:4]),.I4(un2_pre_out_s_11),.LO(N_12_i));
defparam desc450.INIT=32'h33011300;
  LUT6_L desc451(.I0(mult_out_r[0:0]),.I1(mult_out_r[11:11]),.I2(out_inner_prod_r[0:0]),.I3(acc_clear),.I4(out_inner_prod_r[11:11]),.I5(un2_pre_out_s_11),.LO(N_4_i));
defparam desc451.INIT=64'h005A007B0012005A;
  LUT5_L desc452(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[9:9]),.I4(un2_pre_out_s_11),.LO(N_22_i));
defparam desc452.INIT=32'h33011300;
  LUT5_L desc453(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[3:3]),.I4(un2_pre_out_s_11),.LO(N_10_i));
defparam desc453.INIT=32'h33011300;
  LUT5_L desc454(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[2:2]),.I4(un2_pre_out_s_11),.LO(N_8_i));
defparam desc454.INIT=32'h33011300;
  LUT5_L desc455(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out[1:1]),.I4(un2_pre_out_s_11),.LO(N_6_i));
defparam desc455.INIT=32'h33011300;
  LUT5_L desc456(.I0(mult_out_r[11:11]),.I1(acc_clear),.I2(out_inner_prod_r[11:11]),.I3(un2_pre_out_0[10:10]),.I4(un2_pre_out_s_11),.LO(N_24_i));
defparam desc456.INIT=32'h33011300;
  LUT6_L desc457(.I0(mult_out_i[0:0]),.I1(out_inner_prod_i[0:0]),.I2(mult_out_i[11:11]),.I3(acc_clear),.I4(out_inner_prod_i[11:11]),.I5(un2_pre_out_s_11_0),.LO(acc_i_2[0:0]));
defparam desc457.INIT=64'h0066006F00060066;
  LUT6_L desc458(.I0(pipe_counter[2:2]),.I1(in_counter[2:2]),.I2(in_counter[0:0]),.I3(state[1:1]),.I4(state[0:0]),.I5(red_mat_reg),.LO(state_ns[1:1]));
defparam desc458.INIT=64'hF0F05500CCCC5500;
  LUT4_L done_e(.I0(pipe_counter[2:2]),.I1(state[1:1]),.I2(done_inner_prod),.I3(state[0:0]),.LO(done));
defparam done_e.INIT=16'hF0C8;
  LUT6_L desc459(.I0(in_counter[2:2]),.I1(in_counter[0:0]),.I2(state[1:1]),.I3(state[0:0]),.I4(red_mat_reg),.I5(start_inner_prod),.LO(state_ns[0:0]));
defparam desc459.INIT=64'h330F550F33005500;
  LUT5_L in_reg_enable_fsm_e(.I0(state[1:1]),.I1(state[0:0]),.I2(in_reg_enable_fsm),.I3(start_inner_prod),.I4(in_reg_enable_fsm_0_sqmuxa),.LO(in_reg_enable_fsm_0));
defparam in_reg_enable_fsm_e.INIT=32'h3333F1F0;
  LUT5_L desc460(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out[8:8]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[8:8]));
defparam desc460.INIT=32'h33011300;
  LUT5_L desc461(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[4:4]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[4:4]));
defparam desc461.INIT=32'h33011300;
  LUT5_L desc462(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[7:7]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[7:7]));
defparam desc462.INIT=32'h33011300;
  LUT5_L desc463(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[3:3]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[3:3]));
defparam desc463.INIT=32'h33011300;
  LUT5_L desc464(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[5:5]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[5:5]));
defparam desc464.INIT=32'h33011300;
  LUT5_L desc465(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[1:1]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[1:1]));
defparam desc465.INIT=32'h33011300;
  LUT5_L desc466(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[2:2]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[2:2]));
defparam desc466.INIT=32'h33011300;
  LUT5_L desc467(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[9:9]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[9:9]));
defparam desc467.INIT=32'h33011300;
  LUT5_L desc468(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_0[6:6]),.I4(un2_pre_out_s_11_0),.LO(acc_i_2[6:6]));
defparam desc468.INIT=32'h33011300;
  complex_mult_pipe_prod_inj cp_mult(.mult_out_r(mult_out_r[11:0]),.mult_out_i(mult_out_i[11:0]),.in_a_r_reg(in_a_r_reg[11:0]),.in_b_r_reg(in_b_r_reg[11:0]),.in_a_i_reg(in_a_i_reg[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk));
  add_subZ0_add_r_inj add_r(.mult_out_r(mult_out_r[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.un2_pre_out_10(un2_pre_out_0[10:10]),.un2_pre_out_9(un2_pre_out[9:9]),.un2_pre_out_7(un2_pre_out[7:7]),.un2_pre_out_6(un2_pre_out[6:6]),.un2_pre_out_5(un2_pre_out[5:5]),.un2_pre_out_4(un2_pre_out[4:4]),.un2_pre_out_3(un2_pre_out[3:3]),.un2_pre_out_2(un2_pre_out[2:2]),.un2_pre_out_1(un2_pre_out[1:1]),.acc_clear(acc_clear),.un2_pre_out_s_11(un2_pre_out_s_11),.N_26_i(N_26_i),.N_20_i(N_20_i));
  add_subZ0_add_r_1_inj add_i(.mult_out_i(mult_out_i[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.un2_pre_out_10(un2_pre_out[10:10]),.un2_pre_out_9(un2_pre_out_0[9:9]),.un2_pre_out_8(un2_pre_out[8:8]),.un2_pre_out_7(un2_pre_out_0[7:7]),.un2_pre_out_6(un2_pre_out_0[6:6]),.un2_pre_out_5(un2_pre_out_0[5:5]),.un2_pre_out_4(un2_pre_out_0[4:4]),.un2_pre_out_3(un2_pre_out_0[3:3]),.un2_pre_out_2(un2_pre_out_0[2:2]),.un2_pre_out_1(un2_pre_out_0[1:1]),.un2_pre_out_s_11_0(un2_pre_out_s_11_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc469(.I0(in_counter[1:1]),.I1(in_counter[2:2]),.I2(state[0:0]),.I3(un1_state_4_0_0_lut6_2_O6),.O(in_counter_5_43_i_i_a2));
defparam desc469.INIT=16'hA0CC;
  LUT3 desc470(.I0(in_counter[0:0]),.I1(state[0:0]),.I2(un1_state_4_0_0_lut6_2_O6),.O(state_i_0));
defparam desc470.INIT=8'h3A;
  LUT4 desc471(.I0(pipe_counter[1:1]),.I1(pipe_counter[2:2]),.I2(state[0:0]),.I3(un1_state_8_0_0_a2_lut6_2_O5),.O(pipe_counter_4_0_a2[2:2]));
defparam desc471.INIT=16'h0ACC;
  LUT4 desc472(.I0(pipe_counter[0:0]),.I1(pipe_counter[1:1]),.I2(state[0:0]),.I3(un1_state_8_0_0_a2_lut6_2_O5),.O(pipe_counter_4_0_a2[1:1]));
defparam desc472.INIT=16'h0ACC;
  LUT2 un7_acc_enable_lut6_2_o6(.I0(acc_enable),.I1(acc_clear),.O(un7_acc_enable_lut6_2_O6));
defparam un7_acc_enable_lut6_2_o6.INIT=4'hE;
  LUT4 un7_acc_enable_lut6_2_o5(.I0(state[1:1]),.I1(state[0:0]),.I2(acc_clear),.I3(start_inner_prod),.O(acc_clear_0));
defparam un7_acc_enable_lut6_2_o5.INIT=16'hB1A0;
  LUT4 un1_state_8_0_0_a2_lut6_2_o6(.I0(in_counter[2:2]),.I1(in_counter[0:0]),.I2(state[0:0]),.I3(red_mat_reg),.O(in_reg_enable_fsm_0_sqmuxa));
defparam un1_state_8_0_0_a2_lut6_2_o6.INIT=16'hC0A0;
  LUT5 un1_state_8_0_0_a2_lut6_2_o5(.I0(in_counter[2:2]),.I1(in_counter[0:0]),.I2(state[1:1]),.I3(state[0:0]),.I4(red_mat_reg),.O(un1_state_8_0_0_a2_lut6_2_O5));
defparam un1_state_8_0_0_a2_lut6_2_o5.INIT=32'hFCF0FAF0;
  LUT3 un1_state_4_0_0_lut6_2_o6(.I0(state[1:1]),.I1(state[0:0]),.I2(start_inner_prod),.O(un1_state_4_0_0_lut6_2_O6));
defparam un1_state_4_0_0_lut6_2_o6.INIT=8'hDC;
  LUT4 un1_state_4_0_0_lut6_2_o5(.I0(acc_enable),.I1(pipe_counter[2:2]),.I2(state[1:1]),.I3(state[0:0]),.O(acc_enable_0));
defparam un1_state_4_0_0_lut6_2_o5.INIT=16'hFF2A;
  LUT4 desc473(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out_s_11_0),.O(acc_i_2[11:11]));
defparam desc473.INIT=16'h3220;
  LUT5 desc474(.I0(mult_out_i[11:11]),.I1(acc_clear),.I2(out_inner_prod_i[11:11]),.I3(un2_pre_out[10:10]),.I4(un2_pre_out_s_11_0),.O(acc_i_2[10:10]));
defparam desc474.INIT=32'h33011300;
endmodule
module inv_sqrt_inj (out_inner_prod_r,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_8,out_inv_sqrt_7,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_11,out_inv_sqrt_0,done_inv_sqrt,clk,rst,start_inv_sqrt,N_434_i,N_431_i,N_428_i,N_425_i,p_output_reg_pipe_13_Z_p_O_FDshifterZ0_,p_output_reg_pipe_12_Z_p_O_FDshifterZ0_,p_output_reg_pipe_Z_p_O_FDshifterZ0_,p_desc951_p_O_FDE,p_desc952_p_O_FDE,p_desc953_p_O_FDE,p_desc954_p_O_FDE,p_desc955_p_O_FDE,p_desc956_p_O_FDE,p_desc957_p_O_FDE,p_desc958_p_O_FDE,p_desc959_p_O_FDE,p_desc960_p_O_FDE,p_desc961_p_O_FDE,p_desc962_p_O_FDE,p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_,p_output_reg_pipe_Z_p_O_FDRE,p_output_reg_pipe_3_Z_p_O_FDRE,p_output_reg_pipe_6_Z_p_O_FDRE,p_output_reg_pipe_9_Z_p_O_FDRE,p_output_reg_pipe_12_Z_p_O_FDRE,p_output_reg_pipe_15_Z_p_O_FDRE,p_output_reg_pipe_16_Z_p_O_FDRE,p_output_reg_pipe_17_Z_p_O_FDRE,p_output_reg_pipe_18_Z_p_O_FDRE,p_output_reg_pipe_21_Z_p_O_FDRE,p_done_Z_p_O_FDC,p_desc946_p_O_FDC,p_desc947_p_O_FDC,p_desc948_p_O_FDC,p_desc949_p_O_FDC,p_desc950_p_O_FDC);
input [11:0] out_inner_prod_r ;
output out_inv_sqrt_9 ;
output out_inv_sqrt_10 ;
output out_inv_sqrt_8 ;
output out_inv_sqrt_7 ;
output out_inv_sqrt_2 ;
output out_inv_sqrt_1 ;
output out_inv_sqrt_11 ;
output out_inv_sqrt_0 ;
output done_inv_sqrt ;
input clk ;
input rst ;
input start_inv_sqrt ;
output N_434_i ;
output N_431_i ;
output N_428_i ;
output N_425_i ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_11 ;
wire out_inv_sqrt_0 ;
wire done_inv_sqrt ;
wire clk ;
wire rst ;
wire start_inv_sqrt ;
wire N_434_i ;
wire N_431_i ;
wire N_428_i ;
wire N_425_i ;
wire [2:2] ret_val_m10 ;
wire [3:1] ret_val ;
wire [11:11] un1_poly_odd_s_lut6_2_O6 ;
wire [11:0] input_reg ;
wire [3:0] counter ;
wire state ;
wire [3:1] counter_4 ;
wire [11:0] un14_pos_outputf ;
wire [11:0] pre_outputf ;
wire [1:1] out_shift_amount ;
wire [6:5] un7_output_2_1 ;
wire [6:5] un11_output ;
wire [11:0] pre_output ;
wire [7:1] un26_output ;
wire [7:4] un1_input_shifted ;
wire state_i ;
wire [11:1] un14_pos_output ;
wire [9:9] un11_output_6_d_0 ;
wire [11:0] z_5 ;
wire [3:3] ret_val_m2 ;
wire [1:1] ret_val_d_a1 ;
wire [1:1] ret_val_d_a0 ;
wire [10:7] un1_poly_odd ;
wire [10:9] un7 ;
wire [6:2] input_shifted ;
wire ret_val_d_0 ;
wire [1:1] shift_amount_1 ;
wire [2:2] shift_amount_1_i ;
wire [11:11] z_5_i ;
wire [19:9] un8_rnd_out_un0_P ;
wire [23:23] pre_out ;
wire [14:14] un20_output_2 ;
wire [11:11] un1_poly_odd_d ;
wire [6:6] un26_output_0_iv_3 ;
wire [6:6] un26_output_0_iv_2_0 ;
wire [4:4] output_d ;
wire [6:6] un7_output_2_0_0 ;
wire [6:6] un1_poly_odd_i ;
wire [11:0] mult1_out ;
wire [11:0] mult2_out ;
wire N_454 ;
wire un3_shift_right_c2_0_0_a0_1 ;
wire un9_0_axb_8 ;
wire VCC ;
wire m9_a1_1 ;
wire GND ;
wire N_439 ;
wire done ;
wire output_reg_pipe_11 ;
wire N_419 ;
wire un3_shift_right ;
wire z_5_axb_5 ;
wire N_71 ;
wire N_50_i ;
wire output_reg_pipe_12_RNIPJ901_O6 ;
wire N_420 ;
wire output_reg_pipe_17 ;
wire z_axb_0_i ;
wire un9_0_s_2 ;
wire m9_0_0 ;
wire CO1 ;
wire N_62 ;
wire z_5_8_d ;
wire N_414 ;
wire N_417 ;
wire N_33 ;
wire N_31 ;
wire z_5_axb_10 ;
wire un1_apply_nrlt8_1 ;
wire SUM1_0_i_a2_a0_1 ;
wire SUM1_0_i_1_1 ;
wire ret_val_ss0 ;
wire N_458 ;
wire N_378 ;
wire N_13_0 ;
wire N_410 ;
wire N_413 ;
wire N_18_0 ;
wire z_5_axb_7 ;
wire N_80 ;
wire N_51 ;
wire z_5_axb_3 ;
wire N_65 ;
wire un9_0_o5_2 ;
wire N_72 ;
wire un9_0_axb_1 ;
wire un9_0_o5_1 ;
wire un9_0_cry_0_RNO ;
wire N_100_i ;
wire N_79 ;
wire N_50 ;
wire z_5_axb_2 ;
wire un9_0_axb_3 ;
wire un9_0_axb_2 ;
wire ret_val_sm0 ;
wire un4_overflow_2 ;
wire get_m8_0_o4_2 ;
wire N_441 ;
wire un3_shift_right_axb0_i ;
wire un9_0_cry_0_cy ;
wire ret_val_ss3 ;
wire un4_overflow_0 ;
wire PATTERNDETECT_15 ;
wire un2_output_3 ;
wire z_axb_10 ;
wire un1_apply_nrlt7 ;
wire z_axb_9 ;
wire z_axb_8 ;
wire z_axb_7 ;
wire z_axb_6 ;
wire z_axb_5 ;
wire z_axb_4 ;
wire z_axb_3 ;
wire z_axb_2 ;
wire z_axb_1 ;
wire z_axb_0 ;
wire N_45 ;
wire N_70 ;
wire N_73 ;
wire un20_output_0_0_a2_0_0_lut6_2_O5 ;
wire z_5_axb_8 ;
wire un9_0_axb_0 ;
wire N_56 ;
wire N_49 ;
wire z_5_axb_1 ;
wire N_33_0 ;
wire z_5_axb_4 ;
wire z_5_axb_6 ;
wire z_5_axb_9 ;
wire z_5_cry_10 ;
wire z_5_cry_9 ;
wire z_5_cry_8 ;
wire z_5_cry_7 ;
wire z_5_cry_6 ;
wire z_5_cry_5 ;
wire z_5_cry_4 ;
wire z_5_cry_3 ;
wire z_5_cry_2 ;
wire z_5_cry_1 ;
wire z_5_cry_0 ;
wire z_cry_10 ;
wire z_cry_9 ;
wire z_cry_8 ;
wire z_cry_7 ;
wire z_cry_6 ;
wire z_cry_5 ;
wire z_cry_4 ;
wire z_cry_3 ;
wire z_cry_2 ;
wire z_cry_1 ;
wire z_cry_0 ;
wire un9_0_cry_7 ;
wire un9_0_s_8 ;
wire un9_0_cry_6 ;
wire un9_0_s_7 ;
wire N_2502_i ;
wire un9_0_cry_5 ;
wire un9_0_s_6 ;
wire un9_0_cry_4 ;
wire un9_0_s_5 ;
wire un9_0_axb_4 ;
wire un9_0_cry_3 ;
wire un9_0_s_4 ;
wire un9_0_cry_2 ;
wire un9_0_s_3 ;
wire un9_0_cry_1 ;
wire un9_0_cry_0 ;
wire un9_0_s_1 ;
wire un9_0_s_0 ;
input p_output_reg_pipe_13_Z_p_O_FDshifterZ0_ ;
input p_output_reg_pipe_12_Z_p_O_FDshifterZ0_ ;
input p_output_reg_pipe_Z_p_O_FDshifterZ0_ ;
input p_desc951_p_O_FDE ;
input p_desc952_p_O_FDE ;
input p_desc953_p_O_FDE ;
input p_desc954_p_O_FDE ;
input p_desc955_p_O_FDE ;
input p_desc956_p_O_FDE ;
input p_desc957_p_O_FDE ;
input p_desc958_p_O_FDE ;
input p_desc959_p_O_FDE ;
input p_desc960_p_O_FDE ;
input p_desc961_p_O_FDE ;
input p_desc962_p_O_FDE ;
input p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_ ;
input p_output_reg_pipe_Z_p_O_FDRE ;
input p_output_reg_pipe_3_Z_p_O_FDRE ;
input p_output_reg_pipe_6_Z_p_O_FDRE ;
input p_output_reg_pipe_9_Z_p_O_FDRE ;
input p_output_reg_pipe_12_Z_p_O_FDRE ;
input p_output_reg_pipe_15_Z_p_O_FDRE ;
input p_output_reg_pipe_16_Z_p_O_FDRE ;
input p_output_reg_pipe_17_Z_p_O_FDRE ;
input p_output_reg_pipe_18_Z_p_O_FDRE ;
input p_output_reg_pipe_21_Z_p_O_FDRE ;
input p_done_Z_p_O_FDC ;
input p_desc946_p_O_FDC ;
input p_desc947_p_O_FDC ;
input p_desc948_p_O_FDC ;
input p_desc949_p_O_FDC ;
input p_desc950_p_O_FDC ;
// instances
  LUT4 desc944(.I0(un3_shift_right),.I1(un7_output_2_1[5:5]),.I2(un11_output[5:5]),.I3(pre_output[6:6]),.O(z_5_axb_5));
defparam desc944.INIT=16'h27D8;
  LUT4 desc945(.I0(N_71),.I1(un26_output[4:4]),.I2(un3_shift_right),.I3(un9_0_axb_8),.O(un1_input_shifted[7:7]));
defparam desc945.INIT=16'hFFAC;
  p_O_FDC done_Z(.Q(done_inv_sqrt),.D(done),.C(clk),.CLR(rst),.E(p_done_Z_p_O_FDC));
  p_O_FDC desc946(.Q(counter[0:0]),.D(state_i),.C(clk),.CLR(rst),.E(p_desc946_p_O_FDC));
  p_O_FDC desc947(.Q(counter[1:1]),.D(counter_4[1:1]),.C(clk),.CLR(rst),.E(p_desc947_p_O_FDC));
  p_O_FDC desc948(.Q(counter[2:2]),.D(counter_4[2:2]),.C(clk),.CLR(rst),.E(p_desc948_p_O_FDC));
  p_O_FDC desc949(.Q(counter[3:3]),.D(counter_4[3:3]),.C(clk),.CLR(rst),.E(p_desc949_p_O_FDC));
  p_O_FDC desc950(.Q(state),.D(N_50_i),.C(clk),.CLR(rst),.E(p_desc950_p_O_FDC));
  p_O_FDE desc951(.Q(input_reg[11:11]),.D(out_inner_prod_r[11:11]),.C(clk),.CE(start_inv_sqrt),.E(p_desc951_p_O_FDE));
  p_O_FDE desc952(.Q(input_reg[10:10]),.D(out_inner_prod_r[10:10]),.C(clk),.CE(start_inv_sqrt),.E(p_desc952_p_O_FDE));
  p_O_FDE desc953(.Q(input_reg[9:9]),.D(out_inner_prod_r[9:9]),.C(clk),.CE(start_inv_sqrt),.E(p_desc953_p_O_FDE));
  p_O_FDE desc954(.Q(input_reg[8:8]),.D(out_inner_prod_r[8:8]),.C(clk),.CE(start_inv_sqrt),.E(p_desc954_p_O_FDE));
  p_O_FDE desc955(.Q(input_reg[7:7]),.D(out_inner_prod_r[7:7]),.C(clk),.CE(start_inv_sqrt),.E(p_desc955_p_O_FDE));
  p_O_FDE desc956(.Q(input_reg[6:6]),.D(out_inner_prod_r[6:6]),.C(clk),.CE(start_inv_sqrt),.E(p_desc956_p_O_FDE));
  p_O_FDE desc957(.Q(input_reg[5:5]),.D(out_inner_prod_r[5:5]),.C(clk),.CE(start_inv_sqrt),.E(p_desc957_p_O_FDE));
  p_O_FDE desc958(.Q(input_reg[4:4]),.D(out_inner_prod_r[4:4]),.C(clk),.CE(start_inv_sqrt),.E(p_desc958_p_O_FDE));
  p_O_FDE desc959(.Q(input_reg[3:3]),.D(out_inner_prod_r[3:3]),.C(clk),.CE(start_inv_sqrt),.E(p_desc959_p_O_FDE));
  p_O_FDE desc960(.Q(input_reg[2:2]),.D(out_inner_prod_r[2:2]),.C(clk),.CE(start_inv_sqrt),.E(p_desc960_p_O_FDE));
  p_O_FDE desc961(.Q(input_reg[1:1]),.D(out_inner_prod_r[1:1]),.C(clk),.CE(start_inv_sqrt),.E(p_desc961_p_O_FDE));
  p_O_FDE desc962(.Q(input_reg[0:0]),.D(out_inner_prod_r[0:0]),.C(clk),.CE(start_inv_sqrt),.E(p_desc962_p_O_FDE));
  p_O_FDRE output_reg_pipe_Z(.Q(pre_outputf[1:1]),.D(pre_output[1:1]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_Z_p_O_FDRE));
  FDSE output_reg_pipe_1_Z(.Q(un14_pos_outputf[1:1]),.D(un14_pos_output[1:1]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_3_Z(.Q(pre_outputf[2:2]),.D(pre_output[2:2]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_3_Z_p_O_FDRE));
  FDSE output_reg_pipe_4_Z(.Q(un14_pos_outputf[2:2]),.D(un14_pos_output[2:2]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_6_Z(.Q(pre_outputf[7:7]),.D(pre_output[7:7]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_6_Z_p_O_FDRE));
  FDSE output_reg_pipe_7_Z(.Q(un14_pos_outputf[7:7]),.D(un14_pos_output[7:7]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_9_Z(.Q(pre_outputf[8:8]),.D(pre_output[8:8]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_9_Z_p_O_FDRE));
  FDSE output_reg_pipe_10_Z(.Q(un14_pos_outputf[8:8]),.D(un14_pos_output[8:8]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  FDSE output_reg_pipe_11_Z(.Q(output_reg_pipe_11),.D(N_420),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_12_Z(.Q(pre_outputf[10:10]),.D(pre_output[10:10]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_12_Z_p_O_FDRE));
  FDSE output_reg_pipe_13_Z(.Q(un14_pos_outputf[10:10]),.D(un14_pos_output[10:10]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_15_Z(.Q(pre_outputf[11:11]),.D(pre_output[11:11]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_15_Z_p_O_FDRE));
  p_O_FDRE output_reg_pipe_16_Z(.Q(un14_pos_outputf[11:11]),.D(un14_pos_output[11:11]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_16_Z_p_O_FDRE));
  p_O_FDRE output_reg_pipe_17_Z(.Q(output_reg_pipe_17),.D(N_420),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_17_Z_p_O_FDRE));
  p_O_FDRE output_reg_pipe_18_Z(.Q(pre_outputf[0:0]),.D(pre_output[0:0]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_18_Z_p_O_FDRE));
  FDSE output_reg_pipe_19_Z(.Q(un14_pos_outputf[0:0]),.D(z_axb_0_i),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  p_O_FDRE output_reg_pipe_21_Z(.Q(pre_outputf[9:9]),.D(pre_output[9:9]),.C(clk),.R(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt),.E(p_output_reg_pipe_21_Z_p_O_FDRE));
  FDSE output_reg_pipe_22_Z(.Q(un14_pos_outputf[9:9]),.D(un14_pos_output[9:9]),.C(clk),.S(output_reg_pipe_12_RNIPJ901_O6),.CE(done_inv_sqrt));
  LUT4 desc963(.I0(ret_val[3:3]),.I1(m9_a1_1),.I2(un9_0_s_2),.I3(m9_0_0),.O(pre_output[0:0]));
defparam desc963.INIT=16'h5540;
  LUT5 desc964(.I0(ret_val[2:2]),.I1(ret_val[3:3]),.I2(CO1),.I3(un11_output_6_d_0[9:9]),.I4(N_62),.O(z_5_8_d));
defparam desc964.INIT=32'hFE24DA00;
  LUT5 desc965(.I0(ret_val[3:3]),.I1(N_414),.I2(N_417),.I3(N_33),.I4(N_31),.O(z_5_axb_10));
defparam desc965.INIT=32'h0F0FF2F8;
  LUT5 desc966(.I0(ret_val[3:3]),.I1(m9_a1_1),.I2(un9_0_s_2),.I3(m9_0_0),.I4(pre_output[1:1]),.O(z_5[0:0]));
defparam desc966.INIT=32'hAABF5540;
  LUT4 desc967(.I0(un3_shift_right),.I1(un7_output_2_1[6:6]),.I2(un11_output[6:6]),.I3(pre_output[7:7]),.O(un1_apply_nrlt8_1));
defparam desc967.INIT=16'hD800;
  LUT6 desc968(.I0(input_reg[3:3]),.I1(input_reg[4:4]),.I2(input_reg[5:5]),.I3(input_reg[6:6]),.I4(ret_val_m2[3:3]),.I5(N_454),.O(ret_val[3:3]));
defparam desc968.INIT=64'h0003000200000000;
  LUT6 desc969(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(input_reg[10:10]),.I3(input_reg[11:11]),.I4(ret_val_m2[3:3]),.I5(SUM1_0_i_a2_a0_1),.O(SUM1_0_i_1_1));
defparam desc969.INIT=64'hFFF0FFF1FFF0FFF0;
  LUT6 desc970(.I0(ret_val_ss0),.I1(ret_val_d_a1[1:1]),.I2(N_458),.I3(ret_val_d_a0[1:1]),.I4(N_454),.I5(un9_0_axb_8),.O(N_378));
defparam desc970.INIT=64'h5F5CFFCCA0A30033;
  LUT6 desc971(.I0(ret_val_ss0),.I1(ret_val_d_a1[1:1]),.I2(N_458),.I3(ret_val_d_a0[1:1]),.I4(N_454),.I5(un9_0_axb_8),.O(CO1));
defparam desc971.INIT=64'h5F5CFFCC00000000;
  LUT6 desc972(.I0(ret_val[3:3]),.I1(CO1),.I2(N_13_0),.I3(N_410),.I4(N_413),.I5(N_18_0),.O(z_5_axb_7));
defparam desc972.INIT=64'h08807FF77FF70880;
  LUT6 desc973(.I0(ret_val[3:3]),.I1(CO1),.I2(un3_shift_right),.I3(N_80),.I4(N_51),.I5(pre_output[4:4]),.O(z_5_axb_3));
defparam desc973.INIT=64'h080FF8FFF7F00700;
  LUT6 un9_0_o5_2_cZ(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_65),.I3(un26_output[7:7]),.I4(un1_input_shifted[5:5]),.I5(un1_poly_odd[9:9]),.O(un9_0_o5_2));
defparam un9_0_o5_2_cZ.INIT=64'hFFFF5D7F5D7F0000;
  LUT6 un9_0_axb_1_cZ(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_72),.I3(un26_output[5:5]),.I4(un7[10:10]),.I5(un1_poly_odd[10:10]),.O(un9_0_axb_1));
defparam un9_0_axb_1_cZ.INIT=64'h5140AEBFAEBF5140;
  LUT6 un9_0_o5_1_cZ(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_72),.I3(un26_output[5:5]),.I4(un7[10:10]),.I5(un1_poly_odd[10:10]),.O(un9_0_o5_1));
defparam un9_0_o5_1_cZ.INIT=64'hFFFF514051400000;
  LUT4 un9_0_cry_0_RNO_cZ(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_72),.I3(un26_output[5:5]),.O(un9_0_cry_0_RNO));
defparam un9_0_cry_0_RNO_cZ.INIT=16'h082A;
  LUT5 un9_0_cry_4_RNO(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_72),.I3(un26_output[5:5]),.I4(input_shifted[6:6]),.O(un1_poly_odd[7:7]));
defparam un9_0_cry_4_RNO.INIT=32'h0415AEBF;
  LUT6 desc974(.I0(N_100_i),.I1(un3_shift_right),.I2(N_79),.I3(N_50),.I4(N_80),.I5(N_51),.O(z_5_axb_2));
defparam desc974.INIT=64'h02CE20ECCE02EC20;
  LUT6 un9_0_axb_3_cZ(.I0(un9_0_axb_8),.I1(un1_input_shifted[4:4]),.I2(un7[9:9]),.I3(un1_poly_odd[8:8]),.I4(un1_input_shifted[5:5]),.I5(un1_poly_odd[9:9]),.O(un9_0_axb_3));
defparam un9_0_axb_3_cZ.INIT=64'h6699699669969966;
  LUT6 un9_0_axb_2_cZ(.I0(un1_input_shifted[6:6]),.I1(un7[9:9]),.I2(un1_input_shifted[5:5]),.I3(un7[10:10]),.I4(un1_poly_odd[10:10]),.I5(un1_poly_odd[9:9]),.O(un9_0_axb_2));
defparam un9_0_axb_2_cZ.INIT=64'h3C6969C3C396963C;
  LUT6 desc975(.I0(ret_val_sm0),.I1(un4_overflow_2),.I2(get_m8_0_o4_2),.I3(ret_val_ss0),.I4(N_441),.I5(ret_val_d_0),.O(un3_shift_right_axb0_i));
defparam desc975.INIT=64'h00000408FFFFF7FB;
  MUXCY_L un9_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_input_shifted[7:7]),.LO(un9_0_cry_0_cy));
  LUT5 desc976(.I0(ret_val_ss0),.I1(ret_val_d_a1[1:1]),.I2(N_458),.I3(ret_val_d_a0[1:1]),.I4(N_454),.O(ret_val[1:1]));
defparam desc976.INIT=32'h5F5CFFCC;
  LUT4 desc977(.I0(N_454),.I1(SUM1_0_i_1_1),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(shift_amount_1[1:1]));
defparam desc977.INIT=16'hCFEC;
  LUT5 desc978(.I0(N_454),.I1(un3_shift_right_c2_0_0_a0_1),.I2(ret_val[2:2]),.I3(ret_val[1:1]),.I4(un9_0_axb_8),.O(shift_amount_1_i[2:2]));
defparam desc978.INIT=32'h0F7D7D7D;
  LUT4 desc979(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_65),.I3(un26_output[7:7]),.O(un1_input_shifted[4:4]));
defparam desc979.INIT=16'hFBEA;
  LUT4 desc980(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_65),.I3(un26_output[7:7]),.O(un7[9:9]));
defparam desc980.INIT=16'h5D7F;
  LUT1_L desc981(.I0(z_5[11:11]),.LO(z_5_i[11:11]));
defparam desc981.INIT=2'h1;
  LUT2 desc982(.I0(input_reg[1:1]),.I1(input_reg[2:2]),.O(ret_val_sm0));
defparam desc982.INIT=4'hE;
  LUT2 desc983(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.O(un4_overflow_2));
defparam desc983.INIT=4'h1;
  LUT1_L desc984(.I0(state),.LO(state_i));
defparam desc984.INIT=2'h1;
  LUT3 desc985(.I0(un14_pos_outputf[11:11]),.I1(output_reg_pipe_17),.I2(pre_outputf[11:11]),.O(out_inv_sqrt_11));
defparam desc985.INIT=8'hB8;
  LUT3 desc986(.I0(un14_pos_outputf[0:0]),.I1(pre_outputf[0:0]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_0));
defparam desc986.INIT=8'hAC;
  LUT4 desc987(.I0(input_reg[3:3]),.I1(input_reg[7:7]),.I2(input_reg[11:11]),.I3(input_reg[6:6]),.O(get_m8_0_o4_2));
defparam desc987.INIT=16'hFFFE;
  LUT4 desc988(.I0(input_reg[3:3]),.I1(input_reg[4:4]),.I2(input_reg[5:5]),.I3(input_reg[6:6]),.O(N_458));
defparam desc988.INIT=16'h0001;
  LUT3 desc989(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(input_reg[2:2]),.O(ret_val_m2[3:3]));
defparam desc989.INIT=8'hFE;
  LUT4 desc990(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[10:10]),.I3(input_reg[11:11]),.O(ret_val_d_a1[1:1]));
defparam desc990.INIT=16'h000E;
  LUT3 desc991(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[10:10]),.O(N_441));
defparam desc991.INIT=8'hFE;
  LUT3_L desc992(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(input_reg[6:6]),.LO(ret_val_ss3));
defparam desc992.INIT=8'hF2;
  LUT3 desc993(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(input_reg[2:2]),.O(ret_val_ss0));
defparam desc993.INIT=8'hF1;
  LUT3_L desc994(.I0(counter[3:3]),.I1(state),.I2(start_inv_sqrt),.LO(N_50_i));
defparam desc994.INIT=8'h74;
  LUT5_L desc995(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[3:3]),.I3(input_reg[7:7]),.I4(input_reg[6:6]),.LO(SUM1_0_i_a2_a0_1));
defparam desc995.INIT=32'h00000001;
  LUT5 desc996(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[7:7]),.I3(input_reg[10:10]),.I4(input_reg[11:11]),.O(N_454));
defparam desc996.INIT=32'h00000001;
  LUT6 desc997(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(input_reg[7:7]),.I3(input_reg[10:10]),.I4(input_reg[11:11]),.I5(input_reg[6:6]),.O(ret_val_d_a0[1:1]));
defparam desc997.INIT=64'h000000000000000E;
  LUT6 desc998(.I0(input_reg[2:2]),.I1(input_reg[3:3]),.I2(input_reg[7:7]),.I3(input_reg[6:6]),.I4(N_439),.I5(un4_overflow_2),.O(un4_overflow_0));
defparam desc998.INIT=64'h0000000100000000;
  LUT6 desc999(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[7:7]),.I3(input_reg[10:10]),.I4(input_reg[11:11]),.I5(ret_val_ss3),.O(ret_val_d_0));
defparam desc999.INIT=64'h0000FF450000FF44;
  LUT6 desc1000(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(input_reg[7:7]),.I3(input_reg[11:11]),.I4(input_reg[6:6]),.I5(N_441),.O(ret_val[2:2]));
defparam desc1000.INIT=64'h0000000000FF00FE;
  LUT6 desc1001(.I0(input_reg[3:3]),.I1(input_reg[7:7]),.I2(input_reg[6:6]),.I3(un4_overflow_2),.I4(ret_val_m2[3:3]),.I5(N_441),.O(un3_shift_right_c2_0_0_a0_1));
defparam desc1001.INIT=64'h00000F0000000D00;
  LUT5_L desc1002(.I0(z_5[10:10]),.I1(un8_rnd_out_un0_P[19:19]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_10));
defparam desc1002.INIT=32'h99A995A5;
  LUT6 desc1003(.I0(pre_output[0:0]),.I1(pre_output[1:1]),.I2(pre_output[2:2]),.I3(pre_output[4:4]),.I4(pre_output[3:3]),.I5(pre_output[5:5]),.O(un1_apply_nrlt7));
defparam desc1003.INIT=64'hFFFFFFFFFF00E000;
  LUT6 desc1004(.I0(ret_val_sm0),.I1(un4_overflow_2),.I2(get_m8_0_o4_2),.I3(ret_val_ss0),.I4(N_441),.I5(ret_val_d_0),.O(un9_0_axb_8));
defparam desc1004.INIT=64'hFFFFFBF700000804;
  LUT5_L desc1005(.I0(z_5[9:9]),.I1(un8_rnd_out_un0_P[18:18]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_9));
defparam desc1005.INIT=32'h99599A5A;
  LUT5_L desc1006(.I0(z_5[8:8]),.I1(un8_rnd_out_un0_P[17:17]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_8));
defparam desc1006.INIT=32'h99599A5A;
  LUT5_L desc1007(.I0(z_5[7:7]),.I1(un8_rnd_out_un0_P[16:16]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_7));
defparam desc1007.INIT=32'h99599A5A;
  LUT5_L desc1008(.I0(z_5[6:6]),.I1(un8_rnd_out_un0_P[15:15]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_6));
defparam desc1008.INIT=32'h99599A5A;
  LUT5_L desc1009(.I0(z_5[5:5]),.I1(un8_rnd_out_un0_P[14:14]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_5));
defparam desc1009.INIT=32'h99599A5A;
  LUT5_L desc1010(.I0(z_5[4:4]),.I1(un8_rnd_out_un0_P[13:13]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_4));
defparam desc1010.INIT=32'h99599A5A;
  LUT5_L desc1011(.I0(z_5[3:3]),.I1(un8_rnd_out_un0_P[12:12]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_3));
defparam desc1011.INIT=32'h99599A5A;
  LUT5_L desc1012(.I0(z_5[2:2]),.I1(un8_rnd_out_un0_P[11:11]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_2));
defparam desc1012.INIT=32'h99599A5A;
  LUT5_L desc1013(.I0(z_5[1:1]),.I1(un8_rnd_out_un0_P[10:10]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_1));
defparam desc1013.INIT=32'h99599A5A;
  LUT5 desc1014(.I0(z_5[0:0]),.I1(un8_rnd_out_un0_P[9:9]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.O(z_axb_0));
defparam desc1014.INIT=32'h99599A5A;
  LUT5_L desc1015(.I0(z_5[0:0]),.I1(un8_rnd_out_un0_P[9:9]),.I2(pre_out[23:23]),.I3(PATTERNDETECT_15),.I4(un2_output_3),.LO(z_axb_0_i));
defparam desc1015.INIT=32'h66A665A5;
  LUT5 desc1016(.I0(ret_val_m10[2:2]),.I1(N_454),.I2(un3_shift_right_c2_0_0_a0_1),.I3(ret_val[1:1]),.I4(un9_0_axb_8),.O(un3_shift_right));
defparam desc1016.INIT=32'h00D1D1D1;
  LUT6 desc1017(.I0(input_reg[2:2]),.I1(un9_0_axb_8),.I2(un20_output_2[14:14]),.I3(N_45),.I4(shift_amount_1[1:1]),.I5(input_shifted[2:2]),.O(un1_poly_odd_d[11:11]));
defparam desc1017.INIT=64'h03331313CFFFDFDF;
  LUT5 desc1018(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(input_shifted[2:2]),.I3(N_70),.I4(un26_output[3:3]),.O(un1_poly_odd[10:10]));
defparam desc1018.INIT=32'h058D27AF;
  LUT4 desc1019(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_72),.I3(un26_output[5:5]),.O(un1_input_shifted[6:6]));
defparam desc1019.INIT=16'h5140;
  LUT6 desc1020(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_70),.I3(N_71),.I4(un26_output[4:4]),.I5(un26_output[3:3]),.O(un1_poly_odd[9:9]));
defparam desc1020.INIT=64'h048C26AE159D37BF;
  LUT6 desc1021(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_71),.I3(un26_output[4:4]),.I4(N_72),.I5(un26_output[5:5]),.O(un1_poly_odd[8:8]));
defparam desc1021.INIT=64'h04158C9D2637AEBF;
  LUT5 desc1022(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_73),.I3(un26_output_0_iv_3[6:6]),.I4(un26_output_0_iv_2_0[6:6]),.O(un1_input_shifted[5:5]));
defparam desc1022.INIT=32'h51515140;
  LUT5 desc1023(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_73),.I3(un26_output_0_iv_3[6:6]),.I4(un26_output_0_iv_2_0[6:6]),.O(un7[10:10]));
defparam desc1023.INIT=32'h0808082A;
  LUT5 desc1024(.I0(un20_output_0_0_a2_0_0_lut6_2_O5),.I1(un3_shift_right),.I2(un11_output_6_d_0[9:9]),.I3(N_62),.I4(pre_output[8:8]),.O(z_5_axb_8));
defparam desc1024.INIT=32'hCDEF3210;
  LUT5 desc1025(.I0(un9_0_axb_8),.I1(un1_poly_odd_s_lut6_2_O6[11:11]),.I2(un26_output[1:1]),.I3(un1_poly_odd_d[11:11]),.I4(input_shifted[5:5]),.O(un9_0_axb_0));
defparam desc1025.INIT=32'h3F0C95A6;
  LUT5 desc1026(.I0(un20_output_2[14:14]),.I1(un3_shift_right),.I2(N_56),.I3(N_49),.I4(pre_output[2:2]),.O(z_5_axb_1));
defparam desc1026.INIT=32'h13DFEC20;
  LUT5 desc1027(.I0(N_419),.I1(un3_shift_right),.I2(N_33_0),.I3(output_d[4:4]),.I4(pre_output[5:5]),.O(z_5_axb_4));
defparam desc1027.INIT=32'h087FF780;
  LUT5 desc1028(.I0(un3_shift_right),.I1(un7_output_2_0_0[6:6]),.I2(un7_output_2_1[6:6]),.I3(un11_output[6:6]),.I4(pre_output[7:7]),.O(z_5_axb_6));
defparam desc1028.INIT=32'h2A7FD580;
  LUT5 desc1029(.I0(un20_output_0_0_a2_0_0_lut6_2_O5),.I1(un3_shift_right),.I2(un11_output_6_d_0[9:9]),.I3(N_62),.I4(pre_output[10:10]),.O(z_5_axb_9));
defparam desc1029.INIT=32'hCDEF3210;
  XORCY desc1030(.LI(pre_output[11:11]),.CI(z_5_cry_10),.O(z_5[11:11]));
  XORCY desc1031(.LI(z_5_axb_10),.CI(z_5_cry_9),.O(z_5[10:10]));
  MUXCY_L desc1032(.DI(pre_output[10:10]),.CI(z_5_cry_9),.S(z_5_axb_10),.LO(z_5_cry_10));
  XORCY desc1033(.LI(z_5_axb_9),.CI(z_5_cry_8),.O(z_5[9:9]));
  MUXCY_L desc1034(.DI(z_5_8_d),.CI(z_5_cry_8),.S(z_5_axb_9),.LO(z_5_cry_9));
  XORCY desc1035(.LI(z_5_axb_8),.CI(z_5_cry_7),.O(z_5[8:8]));
  MUXCY_L desc1036(.DI(z_5_8_d),.CI(z_5_cry_7),.S(z_5_axb_8),.LO(z_5_cry_8));
  XORCY desc1037(.LI(z_5_axb_7),.CI(z_5_cry_6),.O(z_5[7:7]));
  MUXCY_L desc1038(.DI(pre_output[7:7]),.CI(z_5_cry_6),.S(z_5_axb_7),.LO(z_5_cry_7));
  XORCY desc1039(.LI(z_5_axb_6),.CI(z_5_cry_5),.O(z_5[6:6]));
  MUXCY_L desc1040(.DI(pre_output[6:6]),.CI(z_5_cry_5),.S(z_5_axb_6),.LO(z_5_cry_6));
  XORCY desc1041(.LI(z_5_axb_5),.CI(z_5_cry_4),.O(z_5[5:5]));
  MUXCY_L desc1042(.DI(pre_output[5:5]),.CI(z_5_cry_4),.S(z_5_axb_5),.LO(z_5_cry_5));
  XORCY desc1043(.LI(z_5_axb_4),.CI(z_5_cry_3),.O(z_5[4:4]));
  MUXCY_L desc1044(.DI(pre_output[4:4]),.CI(z_5_cry_3),.S(z_5_axb_4),.LO(z_5_cry_4));
  XORCY desc1045(.LI(z_5_axb_3),.CI(z_5_cry_2),.O(z_5[3:3]));
  MUXCY_L desc1046(.DI(pre_output[3:3]),.CI(z_5_cry_2),.S(z_5_axb_3),.LO(z_5_cry_3));
  XORCY desc1047(.LI(z_5_axb_2),.CI(z_5_cry_1),.O(z_5[2:2]));
  MUXCY_L desc1048(.DI(pre_output[2:2]),.CI(z_5_cry_1),.S(z_5_axb_2),.LO(z_5_cry_2));
  XORCY desc1049(.LI(z_5_axb_1),.CI(z_5_cry_0),.O(z_5[1:1]));
  MUXCY_L desc1050(.DI(pre_output[1:1]),.CI(z_5_cry_0),.S(z_5_axb_1),.LO(z_5_cry_1));
  MUXCY_L desc1051(.DI(pre_output[0:0]),.CI(GND),.S(z_5[0:0]),.LO(z_5_cry_0));
  XORCY desc1052(.LI(z_5_i[11:11]),.CI(z_cry_10),.O(un14_pos_output[11:11]));
  XORCY desc1053(.LI(z_axb_10),.CI(z_cry_9),.O(un14_pos_output[10:10]));
  MUXCY_L desc1054(.DI(z_5[10:10]),.CI(z_cry_9),.S(z_axb_10),.LO(z_cry_10));
  XORCY desc1055(.LI(z_axb_9),.CI(z_cry_8),.O(un14_pos_output[9:9]));
  MUXCY_L desc1056(.DI(z_5[9:9]),.CI(z_cry_8),.S(z_axb_9),.LO(z_cry_9));
  XORCY desc1057(.LI(z_axb_8),.CI(z_cry_7),.O(un14_pos_output[8:8]));
  MUXCY_L desc1058(.DI(z_5[8:8]),.CI(z_cry_7),.S(z_axb_8),.LO(z_cry_8));
  XORCY desc1059(.LI(z_axb_7),.CI(z_cry_6),.O(un14_pos_output[7:7]));
  MUXCY_L desc1060(.DI(z_5[7:7]),.CI(z_cry_6),.S(z_axb_7),.LO(z_cry_7));
  XORCY desc1061(.LI(z_axb_6),.CI(z_cry_5),.O(un14_pos_output[6:6]));
  MUXCY_L desc1062(.DI(z_5[6:6]),.CI(z_cry_5),.S(z_axb_6),.LO(z_cry_6));
  XORCY desc1063(.LI(z_axb_5),.CI(z_cry_4),.O(un14_pos_output[5:5]));
  MUXCY_L desc1064(.DI(z_5[5:5]),.CI(z_cry_4),.S(z_axb_5),.LO(z_cry_5));
  XORCY desc1065(.LI(z_axb_4),.CI(z_cry_3),.O(un14_pos_output[4:4]));
  MUXCY_L desc1066(.DI(z_5[4:4]),.CI(z_cry_3),.S(z_axb_4),.LO(z_cry_4));
  XORCY desc1067(.LI(z_axb_3),.CI(z_cry_2),.O(un14_pos_output[3:3]));
  MUXCY_L desc1068(.DI(z_5[3:3]),.CI(z_cry_2),.S(z_axb_3),.LO(z_cry_3));
  XORCY desc1069(.LI(z_axb_2),.CI(z_cry_1),.O(un14_pos_output[2:2]));
  MUXCY_L desc1070(.DI(z_5[2:2]),.CI(z_cry_1),.S(z_axb_2),.LO(z_cry_2));
  XORCY desc1071(.LI(z_axb_1),.CI(z_cry_0),.O(un14_pos_output[1:1]));
  MUXCY_L desc1072(.DI(z_5[1:1]),.CI(z_cry_0),.S(z_axb_1),.LO(z_cry_1));
  MUXCY_L desc1073(.DI(z_5[0:0]),.CI(VCC),.S(z_axb_0),.LO(z_cry_0));
  XORCY un9_0_s_8_cZ(.LI(un9_0_axb_8),.CI(un9_0_cry_7),.O(un9_0_s_8));
  XORCY un9_0_s_7_cZ(.LI(un3_shift_right_axb0_i),.CI(un9_0_cry_6),.O(un9_0_s_7));
  MUXCY_L un9_0_cry_7_cZ(.DI(VCC),.CI(un9_0_cry_6),.S(un3_shift_right_axb0_i),.LO(un9_0_cry_7));
  XORCY un9_0_s_6_cZ(.LI(N_2502_i),.CI(un9_0_cry_5),.O(un9_0_s_6));
  MUXCY_L un9_0_cry_6_cZ(.DI(VCC),.CI(un9_0_cry_5),.S(N_2502_i),.LO(un9_0_cry_6));
  XORCY un9_0_s_5_cZ(.LI(un1_poly_odd_i[6:6]),.CI(un9_0_cry_4),.O(un9_0_s_5));
  MUXCY_L un9_0_cry_5_cZ(.DI(VCC),.CI(un9_0_cry_4),.S(un1_poly_odd_i[6:6]),.LO(un9_0_cry_5));
  XORCY un9_0_s_4_cZ(.LI(un9_0_axb_4),.CI(un9_0_cry_3),.O(un9_0_s_4));
  MUXCY_L un9_0_cry_4_cZ(.DI(un1_poly_odd[7:7]),.CI(un9_0_cry_3),.S(un9_0_axb_4),.LO(un9_0_cry_4));
  XORCY un9_0_s_3_cZ(.LI(un9_0_axb_3),.CI(un9_0_cry_2),.O(un9_0_s_3));
  MUXCY_L un9_0_cry_3_cZ(.DI(un9_0_o5_2),.CI(un9_0_cry_2),.S(un9_0_axb_3),.LO(un9_0_cry_3));
  XORCY un9_0_s_2_cZ(.LI(un9_0_axb_2),.CI(un9_0_cry_1),.O(un9_0_s_2));
  MUXCY_L un9_0_cry_2_cZ(.DI(un9_0_o5_1),.CI(un9_0_cry_1),.S(un9_0_axb_2),.LO(un9_0_cry_2));
  XORCY un9_0_s_1_cZ(.LI(un9_0_axb_1),.CI(un9_0_cry_0),.O(un9_0_s_1));
  MUXCY_L un9_0_cry_1_cZ(.DI(GND),.CI(un9_0_cry_0),.S(un9_0_axb_1),.LO(un9_0_cry_1));
  XORCY un9_0_s_0_cZ(.LI(un9_0_axb_0),.CI(un9_0_cry_0_cy),.O(un9_0_s_0));
  MUXCY_L un9_0_cry_0_cZ(.DI(un9_0_cry_0_RNO),.CI(un9_0_cry_0_cy),.S(un9_0_axb_0),.LO(un9_0_cry_0));
  shifterZ1_inj in_shift(.ret_val(ret_val[3:1]),.un20_output_2(un20_output_2[14:14]),.ret_val_m2(ret_val_m2[3:3]),.shift_amount_1(shift_amount_1[1:1]),.un26_output_0_iv_3(un26_output_0_iv_3[6:6]),.ret_val_d_a1(ret_val_d_a1[1:1]),.ret_val_d_a0(ret_val_d_a0[1:1]),.un26_output_6(un26_output[7:7]),.un26_output_2(un26_output[3:3]),.un26_output_4(un26_output[5:5]),.un26_output_3(un26_output[4:4]),.un26_output_0(un26_output[1:1]),.un1_poly_odd_i(un1_poly_odd_i[6:6]),.input_reg(input_reg[11:0]),.un26_output_0_iv_2_0_1(un26_output_0_iv_2_0[6:6]),.input_shifted_4(input_shifted[6:6]),.input_shifted_0(input_shifted[2:2]),.input_shifted_3(input_shifted[5:5]),.un1_input_shifted(un1_input_shifted[4:4]),.un1_poly_odd(un1_poly_odd[8:8]),.un9_0_axb_8(un9_0_axb_8),.un20_output_0_0_a2_0_0_lut6_2_O5(un20_output_0_0_a2_0_0_lut6_2_O5),.N_100_i(N_100_i),.N_65(N_65),.un3_shift_right(un3_shift_right),.N_2502_i(N_2502_i),.un4_overflow_2(un4_overflow_2),.N_454(N_454),.N_72(N_72),.ret_val_ss0(ret_val_ss0),.N_458(N_458),.N_45(N_45),.N_70(N_70),.N_73(N_73),.N_71(N_71),.N_441(N_441),.un9_0_axb_4(un9_0_axb_4));
  shifterZ0_inj out_shift(.input_reg(input_reg[11:10]),.shift_amount_1(shift_amount_1[1:1]),.un14_pos_output(un14_pos_output[6:3]),.ret_val(ret_val[3:1]),.un11_output_6_d_0(un11_output_6_d_0[9:9]),.out_shift_amount(out_shift_amount[1:1]),.un7_output_2_0_0(un7_output_2_0_0[6:6]),.un7_output_2_1(un7_output_2_1[6:5]),.output_d(output_d[4:4]),.shift_amount_1_i(shift_amount_1_i[2:2]),.un11_output_1(un11_output[5:5]),.un11_output_2(un11_output[6:6]),.un20_output_2(un20_output_2[14:14]),.pre_output(pre_output[11:1]),.done_inv_sqrt(done_inv_sqrt),.un4_overflow_0(un4_overflow_0),.output_reg_pipe_12_RNIPJ901_O6(output_reg_pipe_12_RNIPJ901_O6),.un9_0_axb_8(un9_0_axb_8),.un9_0_s_6(un9_0_s_6),.un9_0_s_7(un9_0_s_7),.N_414(N_414),.N_33(N_33),.clk(clk),.N_420(N_420),.un3_shift_right(un3_shift_right),.N_410(N_410),.un9_0_s_5(un9_0_s_5),.un9_0_s_8(un9_0_s_8),.N_79(N_79),.N_50(N_50),.un9_0_s_4(un9_0_s_4),.un9_0_s_3(un9_0_s_3),.N_13_0(N_13_0),.N_100_i(N_100_i),.N_31(N_31),.N_18_0(N_18_0),.N_378(N_378),.N_33_0(N_33_0),.N_80(N_80),.N_51(N_51),.un9_0_s_0(un9_0_s_0),.un9_0_s_1(un9_0_s_1),.m9_0_0(m9_0_0),.N_417(N_417),.N_62(N_62),.N_454(N_454),.SUM1_0_i_1_1(SUM1_0_i_1_1),.N_56(N_56),.N_434_i(N_434_i),.N_431_i(N_431_i),.N_428_i(N_428_i),.N_425_i(N_425_i),.un9_0_s_2(un9_0_s_2),.N_419(N_419),.N_49(N_49),.N_413(N_413),.un20_output_0_0_a2_0_0_lut6_2_O5(un20_output_0_0_a2_0_0_lut6_2_O5),.un1_apply_nrlt8_1(un1_apply_nrlt8_1),.un1_apply_nrlt7(un1_apply_nrlt7),.p_output_reg_pipe_13_Z_p_O_FD(p_output_reg_pipe_13_Z_p_O_FDshifterZ0_),.p_output_reg_pipe_12_Z_p_O_FD(p_output_reg_pipe_12_Z_p_O_FDshifterZ0_),.p_output_reg_pipe_Z_p_O_FD(p_output_reg_pipe_Z_p_O_FDshifterZ0_),.p_output_reg_pipe_1_Z_p_O_FDE(p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_4_Z_p_O_FDE(p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_5_Z_p_O_FDE(p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_6_Z_p_O_FDE(p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_9_Z_p_O_FDE(p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_10_Z_p_O_FDE(p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_11_Z_p_O_FDE(p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_14_Z_p_O_FDE(p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_15_Z_p_O_FDE(p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_16_Z_p_O_FDE(p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_),.p_output_reg_pipe_19_Z_p_O_FDE(p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_));
  multiplier_inj desc1074(.mult1_out(mult1_out[11:0]),.pre_output(pre_output[11:0]));
  multiplier_1_inj desc1075(.mult2_out(mult2_out[11:0]),.pre_output(pre_output[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.start_inv_sqrt(start_inv_sqrt),.clk(clk));
  desc940_inj desc1076(.un8_rnd_out_un0_P_9(un8_rnd_out_un0_P[9:9]),.un8_rnd_out_un0_P_10(un8_rnd_out_un0_P[10:10]),.un8_rnd_out_un0_P_11(un8_rnd_out_un0_P[11:11]),.un8_rnd_out_un0_P_12(un8_rnd_out_un0_P[12:12]),.un8_rnd_out_un0_P_13(un8_rnd_out_un0_P[13:13]),.un8_rnd_out_un0_P_14(un8_rnd_out_un0_P[14:14]),.un8_rnd_out_un0_P_15(un8_rnd_out_un0_P[15:15]),.un8_rnd_out_un0_P_16(un8_rnd_out_un0_P[16:16]),.un8_rnd_out_un0_P_17(un8_rnd_out_un0_P[17:17]),.un8_rnd_out_un0_P_18(un8_rnd_out_un0_P[18:18]),.un8_rnd_out_un0_P_19(un8_rnd_out_un0_P[19:19]),.mult1_out(mult1_out[11:0]),.mult2_out(mult2_out[11:0]),.pre_out_23(pre_out[23:23]),.un2_output_3(un2_output_3),.PATTERNDETECT_15(PATTERNDETECT_15));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 desc1077(.I0(N_454),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(out_shift_amount[1:1]));
defparam desc1077.INIT=16'hC623;
  LUT4 desc1078(.I0(N_454),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(N_419));
defparam desc1078.INIT=16'h1DDC;
  LUT2 desc1079(.I0(counter[1:1]),.I1(state),.O(counter_4[2:2]));
defparam desc1079.INIT=4'h8;
  LUT2 desc1080(.I0(counter[2:2]),.I1(state),.O(counter_4[3:3]));
defparam desc1080.INIT=4'h8;
  LUT3 desc1081(.I0(un14_pos_outputf[2:2]),.I1(pre_outputf[2:2]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_2));
defparam desc1081.INIT=8'hAC;
  LUT3 desc1082(.I0(un14_pos_outputf[1:1]),.I1(pre_outputf[1:1]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_1));
defparam desc1082.INIT=8'hAC;
  LUT3 desc1083(.I0(un14_pos_outputf[8:8]),.I1(pre_outputf[8:8]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_8));
defparam desc1083.INIT=8'hAC;
  LUT3 desc1084(.I0(un14_pos_outputf[7:7]),.I1(pre_outputf[7:7]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_7));
defparam desc1084.INIT=8'hAC;
  LUT3 desc1085(.I0(un14_pos_outputf[9:9]),.I1(pre_outputf[9:9]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_9));
defparam desc1085.INIT=8'hAC;
  LUT3 desc1086(.I0(un14_pos_outputf[10:10]),.I1(pre_outputf[10:10]),.I2(output_reg_pipe_11),.O(out_inv_sqrt_10));
defparam desc1086.INIT=8'hAC;
  LUT3 done_e_lut6_2_o6(.I0(counter[3:3]),.I1(state),.I2(done_inv_sqrt),.O(done));
defparam done_e_lut6_2_o6.INIT=8'hC8;
  LUT2 done_e_lut6_2_o5(.I0(counter[0:0]),.I1(state),.O(counter_4[1:1]));
defparam done_e_lut6_2_o5.INIT=4'h8;
  LUT4 desc1087(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[10:10]),.I3(input_reg[11:11]),.O(ret_val_m10[2:2]));
defparam desc1087.INIT=16'h0001;
  LUT2 desc1088(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.O(N_439));
defparam desc1088.INIT=4'hE;
  LUT4 desc1089(.I0(ret_val_m10[2:2]),.I1(N_454),.I2(un3_shift_right_c2_0_0_a0_1),.I3(un9_0_axb_8),.O(un1_poly_odd_s_lut6_2_O6[11:11]));
defparam desc1089.INIT=16'h002E;
  LUT5 desc1090(.I0(ret_val_m10[2:2]),.I1(N_454),.I2(un3_shift_right_c2_0_0_a0_1),.I3(ret_val[1:1]),.I4(un9_0_axb_8),.O(m9_a1_1));
defparam desc1090.INIT=32'h000000D1;
endmodule
module mat_regs_inj (col_sel_AQ2_mux_i_m3_lut6_2_O6,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ_int,w_col_sel_AQ_mux_i_m3_lut6_2_O6,w_col_sel_AQ_mux_i_m3_lut6_2_O5,vec_out_r_AQ_0,vec_in_r_AQ_mux_0_4,vec_in_r_AQ_mux_0_9,vec_in_r_AQ_mux_0_6,vec_in_r_AQ_mux_0_0,vec_in_r_AQ_mux_0_1,vec_in_r_AQ_mux_0_2,vec_in_r_AQ_mux_0_3,vec_in_r_AQ_mux_0_10,vec_in_r_AQ_mux_0_7,vec_in_r_AQ_mux_0_8,vec_out_r_AQ_3,vec_in_r_AQ_mux_3,out_Q_r,vec_out_r_AQ_2,vec_out_r_AQ_1,vec_in_r_AQ_mux_2,vec_in_r_AQ_mux_1,vec_out_i_AQ_0,vec_in_i_AQ_mux_0_5,vec_in_i_AQ_mux_0_10,vec_in_i_AQ_mux_0_7,vec_in_i_AQ_mux_0_0,vec_in_i_AQ_mux_0_1,vec_in_i_AQ_mux_0_4,vec_in_i_AQ_mux_0_6,vec_in_i_AQ_mux_0_11,vec_in_i_AQ_mux_0_8,vec_in_i_AQ_mux_0_9,vec_out_i_AQ_3,vec_in_i_AQ_mux_3,out_Q_i,vec_out_i_AQ_2,vec_out_i_AQ_1,vec_in_i_AQ_mux_2,vec_in_i_AQ_mux_1,row_sel_AQ,single_out_r_AQ2_1,single_out_r_AQ2_6,single_out_r_AQ2_4,single_out_r_AQ2_0,single_out_i_AQ2_1,single_out_i_AQ2_5,single_out_i_AQ2_4,single_out_i_AQ2_0,single_out_i_AQ2_11,single_out_i_AQ_1,single_out_i_AQ_0,single_out_i_AQ_8,single_out_i_AQ_10,single_out_i_AQ_11,single_out_i_AQ_9,single_out_i_AQ_4,single_out_r_AQ_4,single_out_r_AQ_2,single_out_r_AQ_7,single_out_r_AQ_1,single_out_r_AQ_0,clk,wr_en_AQ_mux_i_m3_lut6_2_O6,N_507,N_508,N_505,N_506,N_645,N_641,N_637,N_632,N_628,N_624,N_623,N_622,N_612,N_607,N_606,N_605,N_597,N_596,N_595,N_586,N_585,N_584,N_583,N_582,N_571,N_568,N_567,N_566,N_555,N_552,N_549);
input col_sel_AQ2_mux_i_m3_lut6_2_O6 ;
input col_sel_AQ2_mux_i_m3_lut6_2_O5 ;
input [1:0] col_sel_AQ_int ;
input w_col_sel_AQ_mux_i_m3_lut6_2_O6 ;
input w_col_sel_AQ_mux_i_m3_lut6_2_O5 ;
output [11:0] vec_out_r_AQ_0 ;
input vec_in_r_AQ_mux_0_4 ;
input vec_in_r_AQ_mux_0_9 ;
input vec_in_r_AQ_mux_0_6 ;
input vec_in_r_AQ_mux_0_0 ;
input vec_in_r_AQ_mux_0_1 ;
input vec_in_r_AQ_mux_0_2 ;
input vec_in_r_AQ_mux_0_3 ;
input vec_in_r_AQ_mux_0_10 ;
input vec_in_r_AQ_mux_0_7 ;
input vec_in_r_AQ_mux_0_8 ;
output [11:0] vec_out_r_AQ_3 ;
input [11:0] vec_in_r_AQ_mux_3 ;
output [47:0] out_Q_r ;
output [11:0] vec_out_r_AQ_2 ;
output [11:0] vec_out_r_AQ_1 ;
input [11:0] vec_in_r_AQ_mux_2 ;
input [11:0] vec_in_r_AQ_mux_1 ;
output [11:0] vec_out_i_AQ_0 ;
input vec_in_i_AQ_mux_0_5 ;
input vec_in_i_AQ_mux_0_10 ;
input vec_in_i_AQ_mux_0_7 ;
input vec_in_i_AQ_mux_0_0 ;
input vec_in_i_AQ_mux_0_1 ;
input vec_in_i_AQ_mux_0_4 ;
input vec_in_i_AQ_mux_0_6 ;
input vec_in_i_AQ_mux_0_11 ;
input vec_in_i_AQ_mux_0_8 ;
input vec_in_i_AQ_mux_0_9 ;
output [11:0] vec_out_i_AQ_3 ;
input [11:0] vec_in_i_AQ_mux_3 ;
output [47:0] out_Q_i ;
output [11:0] vec_out_i_AQ_2 ;
output [11:0] vec_out_i_AQ_1 ;
input [11:0] vec_in_i_AQ_mux_2 ;
input [11:0] vec_in_i_AQ_mux_1 ;
input [1:0] row_sel_AQ ;
output single_out_r_AQ2_1 ;
output single_out_r_AQ2_6 ;
output single_out_r_AQ2_4 ;
output single_out_r_AQ2_0 ;
output single_out_i_AQ2_1 ;
output single_out_i_AQ2_5 ;
output single_out_i_AQ2_4 ;
output single_out_i_AQ2_0 ;
output single_out_i_AQ2_11 ;
output single_out_i_AQ_1 ;
output single_out_i_AQ_0 ;
output single_out_i_AQ_8 ;
output single_out_i_AQ_10 ;
output single_out_i_AQ_11 ;
output single_out_i_AQ_9 ;
output single_out_i_AQ_4 ;
output single_out_r_AQ_4 ;
output single_out_r_AQ_2 ;
output single_out_r_AQ_7 ;
output single_out_r_AQ_1 ;
output single_out_r_AQ_0 ;
input clk ;
input wr_en_AQ_mux_i_m3_lut6_2_O6 ;
input N_507 ;
input N_508 ;
input N_505 ;
input N_506 ;
output N_645 ;
output N_641 ;
output N_637 ;
output N_632 ;
output N_628 ;
output N_624 ;
output N_623 ;
output N_622 ;
output N_612 ;
output N_607 ;
output N_606 ;
output N_605 ;
output N_597 ;
output N_596 ;
output N_595 ;
output N_586 ;
output N_585 ;
output N_584 ;
output N_583 ;
output N_582 ;
output N_571 ;
output N_568 ;
output N_567 ;
output N_566 ;
output N_555 ;
output N_552 ;
output N_549 ;
wire vec_in_r_AQ_mux_0_4 ;
wire vec_in_r_AQ_mux_0_9 ;
wire vec_in_r_AQ_mux_0_6 ;
wire vec_in_r_AQ_mux_0_0 ;
wire vec_in_r_AQ_mux_0_1 ;
wire vec_in_r_AQ_mux_0_2 ;
wire vec_in_r_AQ_mux_0_3 ;
wire vec_in_r_AQ_mux_0_10 ;
wire vec_in_r_AQ_mux_0_7 ;
wire vec_in_r_AQ_mux_0_8 ;
wire vec_in_i_AQ_mux_0_5 ;
wire vec_in_i_AQ_mux_0_10 ;
wire vec_in_i_AQ_mux_0_7 ;
wire vec_in_i_AQ_mux_0_0 ;
wire vec_in_i_AQ_mux_0_1 ;
wire vec_in_i_AQ_mux_0_4 ;
wire vec_in_i_AQ_mux_0_6 ;
wire vec_in_i_AQ_mux_0_11 ;
wire vec_in_i_AQ_mux_0_8 ;
wire vec_in_i_AQ_mux_0_9 ;
wire single_out_r_AQ2_1 ;
wire single_out_r_AQ2_6 ;
wire single_out_r_AQ2_4 ;
wire single_out_r_AQ2_0 ;
wire single_out_i_AQ2_1 ;
wire single_out_i_AQ2_5 ;
wire single_out_i_AQ2_4 ;
wire single_out_i_AQ2_0 ;
wire single_out_i_AQ2_11 ;
wire single_out_i_AQ_1 ;
wire single_out_i_AQ_0 ;
wire single_out_i_AQ_8 ;
wire single_out_i_AQ_10 ;
wire single_out_i_AQ_11 ;
wire single_out_i_AQ_9 ;
wire single_out_i_AQ_4 ;
wire single_out_r_AQ_4 ;
wire single_out_r_AQ_2 ;
wire single_out_r_AQ_7 ;
wire single_out_r_AQ_1 ;
wire single_out_r_AQ_0 ;
wire clk ;
wire wr_en_AQ_mux_i_m3_lut6_2_O6 ;
wire N_507 ;
wire N_508 ;
wire N_505 ;
wire N_506 ;
wire N_645 ;
wire N_641 ;
wire N_637 ;
wire N_632 ;
wire N_628 ;
wire N_624 ;
wire N_623 ;
wire N_622 ;
wire N_612 ;
wire N_607 ;
wire N_606 ;
wire N_605 ;
wire N_597 ;
wire N_596 ;
wire N_595 ;
wire N_586 ;
wire N_585 ;
wire N_584 ;
wire N_583 ;
wire N_582 ;
wire N_571 ;
wire N_568 ;
wire N_567 ;
wire N_566 ;
wire N_555 ;
wire N_552 ;
wire N_549 ;
wire [1:0] mat_r_1_I_47_DOC ;
wire [1:0] mat_r_1_I_47_DOD ;
wire [1:0] mat_r_1_I_45_DOC ;
wire [1:0] mat_r_1_I_45_DOD ;
wire [1:0] mat_r_1_I_43_DOC ;
wire [1:0] mat_r_1_I_43_DOD ;
wire [1:0] mat_r_1_I_41_DOC ;
wire [1:0] mat_r_1_I_41_DOD ;
wire [1:0] mat_r_1_I_39_DOC ;
wire [1:0] mat_r_1_I_39_DOD ;
wire [1:0] mat_r_1_I_37_DOC ;
wire [1:0] mat_r_1_I_37_DOD ;
wire [1:0] mat_r_1_I_35_DOC ;
wire [1:0] mat_r_1_I_35_DOD ;
wire [1:0] mat_r_1_I_33_DOC ;
wire [1:0] mat_r_1_I_33_DOD ;
wire [1:0] mat_r_1_I_31_DOC ;
wire [1:0] mat_r_1_I_31_DOD ;
wire [1:0] mat_r_1_I_29_DOC ;
wire [1:0] mat_r_1_I_29_DOD ;
wire [1:0] mat_r_1_I_27_DOC ;
wire [1:0] mat_r_1_I_27_DOD ;
wire [1:0] mat_r_1_I_25_DOC ;
wire [1:0] mat_r_1_I_25_DOD ;
wire [1:0] mat_r_1_I_23_DOC ;
wire [1:0] mat_r_1_I_23_DOD ;
wire [1:0] mat_r_1_I_21_DOC ;
wire [1:0] mat_r_1_I_21_DOD ;
wire [1:0] mat_r_1_I_19_DOC ;
wire [1:0] mat_r_1_I_19_DOD ;
wire [1:0] mat_r_1_I_17_DOC ;
wire [1:0] mat_r_1_I_17_DOD ;
wire [1:0] mat_r_1_I_15_DOC ;
wire [1:0] mat_r_1_I_15_DOD ;
wire [1:0] mat_r_1_I_13_DOC ;
wire [1:0] mat_r_1_I_13_DOD ;
wire [1:0] mat_r_1_I_11_DOC ;
wire [1:0] mat_r_1_I_11_DOD ;
wire [1:0] mat_r_1_I_9_DOC ;
wire [1:0] mat_r_1_I_9_DOD ;
wire [1:0] mat_r_1_I_7_DOC ;
wire [1:0] mat_r_1_I_7_DOD ;
wire [1:0] mat_r_1_I_5_DOC ;
wire [1:0] mat_r_1_I_5_DOD ;
wire [1:0] mat_r_1_I_3_DOC ;
wire [1:0] mat_r_1_I_3_DOD ;
wire [1:0] mat_r_1_I_1_DOC ;
wire [1:0] mat_r_1_I_1_DOD ;
wire [1:0] mat_i_1_I_47_DOC ;
wire [1:0] mat_i_1_I_47_DOD ;
wire [1:0] mat_i_1_I_45_DOC ;
wire [1:0] mat_i_1_I_45_DOD ;
wire [1:0] mat_i_1_I_43_DOC ;
wire [1:0] mat_i_1_I_43_DOD ;
wire [1:0] mat_i_1_I_41_DOC ;
wire [1:0] mat_i_1_I_41_DOD ;
wire [1:0] mat_i_1_I_39_DOC ;
wire [1:0] mat_i_1_I_39_DOD ;
wire [1:0] mat_i_1_I_37_DOC ;
wire [1:0] mat_i_1_I_37_DOD ;
wire [1:0] mat_i_1_I_35_DOC ;
wire [1:0] mat_i_1_I_35_DOD ;
wire [1:0] mat_i_1_I_33_DOC ;
wire [1:0] mat_i_1_I_33_DOD ;
wire [1:0] mat_i_1_I_31_DOC ;
wire [1:0] mat_i_1_I_31_DOD ;
wire [1:0] mat_i_1_I_29_DOC ;
wire [1:0] mat_i_1_I_29_DOD ;
wire [1:0] mat_i_1_I_27_DOC ;
wire [1:0] mat_i_1_I_27_DOD ;
wire [1:0] mat_i_1_I_25_DOC ;
wire [1:0] mat_i_1_I_25_DOD ;
wire [1:0] mat_i_1_I_23_DOC ;
wire [1:0] mat_i_1_I_23_DOD ;
wire [1:0] mat_i_1_I_21_DOC ;
wire [1:0] mat_i_1_I_21_DOD ;
wire [1:0] mat_i_1_I_19_DOC ;
wire [1:0] mat_i_1_I_19_DOD ;
wire [1:0] mat_i_1_I_17_DOC ;
wire [1:0] mat_i_1_I_17_DOD ;
wire [1:0] mat_i_1_I_15_DOC ;
wire [1:0] mat_i_1_I_15_DOD ;
wire [1:0] mat_i_1_I_13_DOC ;
wire [1:0] mat_i_1_I_13_DOD ;
wire [1:0] mat_i_1_I_11_DOC ;
wire [1:0] mat_i_1_I_11_DOD ;
wire [1:0] mat_i_1_I_9_DOC ;
wire [1:0] mat_i_1_I_9_DOD ;
wire [1:0] mat_i_1_I_7_DOC ;
wire [1:0] mat_i_1_I_7_DOD ;
wire [1:0] mat_i_1_I_5_DOC ;
wire [1:0] mat_i_1_I_5_DOD ;
wire [1:0] mat_i_1_I_3_DOC ;
wire [1:0] mat_i_1_I_3_DOD ;
wire [1:0] mat_i_1_I_1_DOC ;
wire [1:0] mat_i_1_I_1_DOD ;
wire GND ;
wire VCC ;
// instances
  RAM32M mat_r_1_I_47(.DOA({out_Q_r[8:8],out_Q_r[5:5]}),.DOB({vec_out_r_AQ_3[8:8],vec_out_r_AQ_3[5:5]}),.DOC(mat_r_1_I_47_DOC[1:0]),.DOD(mat_r_1_I_47_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[8:8],vec_in_r_AQ_mux_3[5:5]}),.DIB({vec_in_r_AQ_mux_3[8:8],vec_in_r_AQ_mux_3[5:5]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_47.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_47.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_47.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_47.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_45(.DOA({out_Q_r[41:41],out_Q_r[19:19]}),.DOB({vec_out_r_AQ_0[5:5],vec_out_r_AQ_2[7:7]}),.DOC(mat_r_1_I_45_DOC[1:0]),.DOD(mat_r_1_I_45_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_4,vec_in_r_AQ_mux_2[7:7]}),.DIB({vec_in_r_AQ_mux_0_4,vec_in_r_AQ_mux_2[7:7]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_45.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_45.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_45.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_45.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_43(.DOA({out_Q_r[46:46],out_Q_r[2:2]}),.DOB({vec_out_r_AQ_0[10:10],vec_out_r_AQ_3[2:2]}),.DOC(mat_r_1_I_43_DOC[1:0]),.DOD(mat_r_1_I_43_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_9,vec_in_r_AQ_mux_3[2:2]}),.DIB({vec_in_r_AQ_mux_0_9,vec_in_r_AQ_mux_3[2:2]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_43.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_43.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_43.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_43.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_41(.DOA({out_Q_r[32:32],out_Q_r[20:20]}),.DOB({vec_out_r_AQ_1[8:8],vec_out_r_AQ_2[8:8]}),.DOC(mat_r_1_I_41_DOC[1:0]),.DOD(mat_r_1_I_41_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_1[8:8],vec_in_r_AQ_mux_2[8:8]}),.DIB({vec_in_r_AQ_mux_1[8:8],vec_in_r_AQ_mux_2[8:8]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_41.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_41.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_41.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_41.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_39(.DOA({out_Q_r[43:43],out_Q_r[21:21]}),.DOB({vec_out_r_AQ_0[7:7],vec_out_r_AQ_2[9:9]}),.DOC(mat_r_1_I_39_DOC[1:0]),.DOD(mat_r_1_I_39_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_6,vec_in_r_AQ_mux_2[9:9]}),.DIB({vec_in_r_AQ_mux_0_6,vec_in_r_AQ_mux_2[9:9]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_39.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_39.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_39.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_39.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_37(.DOA({out_Q_r[26:26],out_Q_r[35:35]}),.DOB({vec_out_r_AQ_1[2:2],vec_out_r_AQ_1[11:11]}),.DOC(mat_r_1_I_37_DOC[1:0]),.DOD(mat_r_1_I_37_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_1[2:2],vec_in_r_AQ_mux_1[11:11]}),.DIB({vec_in_r_AQ_mux_1[2:2],vec_in_r_AQ_mux_1[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_37.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_37.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_37.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_37.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_35(.DOA({out_Q_r[22:22],out_Q_r[18:18]}),.DOB({vec_out_r_AQ_2[10:10],vec_out_r_AQ_2[6:6]}),.DOC(mat_r_1_I_35_DOC[1:0]),.DOD(mat_r_1_I_35_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_2[10:10],vec_in_r_AQ_mux_2[6:6]}),.DIB({vec_in_r_AQ_mux_2[10:10],vec_in_r_AQ_mux_2[6:6]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_35.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_35.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_35.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_35.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_33(.DOA({out_Q_r[36:36],out_Q_r[23:23]}),.DOB({vec_out_r_AQ_0[0:0],vec_out_r_AQ_2[11:11]}),.DOC(mat_r_1_I_33_DOC[1:0]),.DOD(mat_r_1_I_33_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({N_507,vec_in_r_AQ_mux_2[11:11]}),.DIB({N_507,vec_in_r_AQ_mux_2[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_33.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_33.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_33.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_33.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_31(.DOA({out_Q_r[10:10],out_Q_r[37:37]}),.DOB({vec_out_r_AQ_3[10:10],vec_out_r_AQ_0[1:1]}),.DOC(mat_r_1_I_31_DOC[1:0]),.DOD(mat_r_1_I_31_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[10:10],vec_in_r_AQ_mux_0_0}),.DIB({vec_in_r_AQ_mux_3[10:10],vec_in_r_AQ_mux_0_0}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_31.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_31.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_31.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_31.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_29(.DOA({out_Q_r[24:24],out_Q_r[11:11]}),.DOB({vec_out_r_AQ_1[0:0],vec_out_r_AQ_3[11:11]}),.DOC(mat_r_1_I_29_DOC[1:0]),.DOD(mat_r_1_I_29_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_1[0:0],vec_in_r_AQ_mux_3[11:11]}),.DIB({vec_in_r_AQ_mux_1[0:0],vec_in_r_AQ_mux_3[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_29.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_29.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_29.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_29.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_27(.DOA({out_Q_r[38:38],out_Q_r[25:25]}),.DOB({vec_out_r_AQ_0[2:2],vec_out_r_AQ_1[1:1]}),.DOC(mat_r_1_I_27_DOC[1:0]),.DOD(mat_r_1_I_27_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_1,vec_in_r_AQ_mux_1[1:1]}),.DIB({vec_in_r_AQ_mux_0_1,vec_in_r_AQ_mux_1[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_27.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_27.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_27.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_27.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_25(.DOA({out_Q_r[12:12],out_Q_r[39:39]}),.DOB({vec_out_r_AQ_2[0:0],vec_out_r_AQ_0[3:3]}),.DOC(mat_r_1_I_25_DOC[1:0]),.DOD(mat_r_1_I_25_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_2[0:0],vec_in_r_AQ_mux_0_2}),.DIB({vec_in_r_AQ_mux_2[0:0],vec_in_r_AQ_mux_0_2}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_25.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_25.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_25.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_25.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_23(.DOA({out_Q_r[9:9],out_Q_r[13:13]}),.DOB({vec_out_r_AQ_3[9:9],vec_out_r_AQ_2[1:1]}),.DOC(mat_r_1_I_23_DOC[1:0]),.DOD(mat_r_1_I_23_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[9:9],vec_in_r_AQ_mux_2[1:1]}),.DIB({vec_in_r_AQ_mux_3[9:9],vec_in_r_AQ_mux_2[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_23.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_23.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_23.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_23.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_21(.DOA({out_Q_r[40:40],out_Q_r[27:27]}),.DOB({vec_out_r_AQ_0[4:4],vec_out_r_AQ_1[3:3]}),.DOC(mat_r_1_I_21_DOC[1:0]),.DOD(mat_r_1_I_21_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_3,vec_in_r_AQ_mux_1[3:3]}),.DIB({vec_in_r_AQ_mux_0_3,vec_in_r_AQ_mux_1[3:3]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_21.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_21.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_21.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_21.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_19(.DOA({out_Q_r[14:14],out_Q_r[0:0]}),.DOB({vec_out_r_AQ_2[2:2],vec_out_r_AQ_3[0:0]}),.DOC(mat_r_1_I_19_DOC[1:0]),.DOD(mat_r_1_I_19_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_2[2:2],vec_in_r_AQ_mux_3[0:0]}),.DIB({vec_in_r_AQ_mux_2[2:2],vec_in_r_AQ_mux_3[0:0]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_19.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_19.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_19.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_19.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_17(.DOA({out_Q_r[6:6],out_Q_r[34:34]}),.DOB({vec_out_r_AQ_3[6:6],vec_out_r_AQ_1[10:10]}),.DOC(mat_r_1_I_17_DOC[1:0]),.DOD(mat_r_1_I_17_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[6:6],vec_in_r_AQ_mux_1[10:10]}),.DIB({vec_in_r_AQ_mux_3[6:6],vec_in_r_AQ_mux_1[10:10]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_17.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_17.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_17.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_17.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_15(.DOA({out_Q_r[42:42],out_Q_r[1:1]}),.DOB({vec_out_r_AQ_0[6:6],vec_out_r_AQ_3[1:1]}),.DOC(mat_r_1_I_15_DOC[1:0]),.DOD(mat_r_1_I_15_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({N_508,vec_in_r_AQ_mux_3[1:1]}),.DIB({N_508,vec_in_r_AQ_mux_3[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_15.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_15.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_15.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_15.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_13(.DOA({out_Q_r[7:7],out_Q_r[47:47]}),.DOB({vec_out_r_AQ_3[7:7],vec_out_r_AQ_0[11:11]}),.DOC(mat_r_1_I_13_DOC[1:0]),.DOD(mat_r_1_I_13_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[7:7],vec_in_r_AQ_mux_0_10}),.DIB({vec_in_r_AQ_mux_3[7:7],vec_in_r_AQ_mux_0_10}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_13.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_13.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_13.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_13.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_11(.DOA({out_Q_r[30:30],out_Q_r[17:17]}),.DOB({vec_out_r_AQ_1[6:6],vec_out_r_AQ_2[5:5]}),.DOC(mat_r_1_I_11_DOC[1:0]),.DOD(mat_r_1_I_11_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_1[6:6],vec_in_r_AQ_mux_2[5:5]}),.DIB({vec_in_r_AQ_mux_1[6:6],vec_in_r_AQ_mux_2[5:5]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_11.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_11.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_11.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_11.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_9(.DOA({out_Q_r[44:44],out_Q_r[31:31]}),.DOB({vec_out_r_AQ_0[8:8],vec_out_r_AQ_1[7:7]}),.DOC(mat_r_1_I_9_DOC[1:0]),.DOD(mat_r_1_I_9_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_0_7,vec_in_r_AQ_mux_1[7:7]}),.DIB({vec_in_r_AQ_mux_0_7,vec_in_r_AQ_mux_1[7:7]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_9.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_9.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_9.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_9.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_7(.DOA({out_Q_r[3:3],out_Q_r[45:45]}),.DOB({vec_out_r_AQ_3[3:3],vec_out_r_AQ_0[9:9]}),.DOC(mat_r_1_I_7_DOC[1:0]),.DOD(mat_r_1_I_7_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[3:3],vec_in_r_AQ_mux_0_8}),.DIB({vec_in_r_AQ_mux_3[3:3],vec_in_r_AQ_mux_0_8}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_7.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_7.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_7.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_7.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_5(.DOA({out_Q_r[4:4],out_Q_r[28:28]}),.DOB({vec_out_r_AQ_3[4:4],vec_out_r_AQ_1[4:4]}),.DOC(mat_r_1_I_5_DOC[1:0]),.DOD(mat_r_1_I_5_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_3[4:4],vec_in_r_AQ_mux_1[4:4]}),.DIB({vec_in_r_AQ_mux_3[4:4],vec_in_r_AQ_mux_1[4:4]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_5.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_5.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_5.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_5.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_3(.DOA({out_Q_r[15:15],out_Q_r[33:33]}),.DOB({vec_out_r_AQ_2[3:3],vec_out_r_AQ_1[9:9]}),.DOC(mat_r_1_I_3_DOC[1:0]),.DOD(mat_r_1_I_3_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_2[3:3],vec_in_r_AQ_mux_1[9:9]}),.DIB({vec_in_r_AQ_mux_2[3:3],vec_in_r_AQ_mux_1[9:9]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_3.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_3.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_3.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_3.INIT_D=64'h0000000000000000;
  RAM32M mat_r_1_I_1(.DOA({out_Q_r[29:29],out_Q_r[16:16]}),.DOB({vec_out_r_AQ_1[5:5],vec_out_r_AQ_2[4:4]}),.DOC(mat_r_1_I_1_DOC[1:0]),.DOD(mat_r_1_I_1_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_r_AQ_mux_1[5:5],vec_in_r_AQ_mux_2[4:4]}),.DIB({vec_in_r_AQ_mux_1[5:5],vec_in_r_AQ_mux_2[4:4]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_r_1_I_1.INIT_A=64'h0000000000000000;
defparam mat_r_1_I_1.INIT_B=64'h0000000000000000;
defparam mat_r_1_I_1.INIT_C=64'h0000000000000000;
defparam mat_r_1_I_1.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_47(.DOA({out_Q_i[8:8],out_Q_i[5:5]}),.DOB({vec_out_i_AQ_3[8:8],vec_out_i_AQ_3[5:5]}),.DOC(mat_i_1_I_47_DOC[1:0]),.DOD(mat_i_1_I_47_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[8:8],vec_in_i_AQ_mux_3[5:5]}),.DIB({vec_in_i_AQ_mux_3[8:8],vec_in_i_AQ_mux_3[5:5]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_47.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_47.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_47.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_47.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_45(.DOA({out_Q_i[41:41],out_Q_i[19:19]}),.DOB({vec_out_i_AQ_0[5:5],vec_out_i_AQ_2[7:7]}),.DOC(mat_i_1_I_45_DOC[1:0]),.DOD(mat_i_1_I_45_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_5,vec_in_i_AQ_mux_2[7:7]}),.DIB({vec_in_i_AQ_mux_0_5,vec_in_i_AQ_mux_2[7:7]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_45.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_45.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_45.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_45.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_43(.DOA({out_Q_i[46:46],out_Q_i[2:2]}),.DOB({vec_out_i_AQ_0[10:10],vec_out_i_AQ_3[2:2]}),.DOC(mat_i_1_I_43_DOC[1:0]),.DOD(mat_i_1_I_43_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_10,vec_in_i_AQ_mux_3[2:2]}),.DIB({vec_in_i_AQ_mux_0_10,vec_in_i_AQ_mux_3[2:2]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_43.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_43.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_43.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_43.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_41(.DOA({out_Q_i[32:32],out_Q_i[20:20]}),.DOB({vec_out_i_AQ_1[8:8],vec_out_i_AQ_2[8:8]}),.DOC(mat_i_1_I_41_DOC[1:0]),.DOD(mat_i_1_I_41_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_1[8:8],vec_in_i_AQ_mux_2[8:8]}),.DIB({vec_in_i_AQ_mux_1[8:8],vec_in_i_AQ_mux_2[8:8]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_41.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_41.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_41.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_41.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_39(.DOA({out_Q_i[43:43],out_Q_i[21:21]}),.DOB({vec_out_i_AQ_0[7:7],vec_out_i_AQ_2[9:9]}),.DOC(mat_i_1_I_39_DOC[1:0]),.DOD(mat_i_1_I_39_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_7,vec_in_i_AQ_mux_2[9:9]}),.DIB({vec_in_i_AQ_mux_0_7,vec_in_i_AQ_mux_2[9:9]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_39.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_39.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_39.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_39.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_37(.DOA({out_Q_i[26:26],out_Q_i[35:35]}),.DOB({vec_out_i_AQ_1[2:2],vec_out_i_AQ_1[11:11]}),.DOC(mat_i_1_I_37_DOC[1:0]),.DOD(mat_i_1_I_37_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_1[2:2],vec_in_i_AQ_mux_1[11:11]}),.DIB({vec_in_i_AQ_mux_1[2:2],vec_in_i_AQ_mux_1[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_37.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_37.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_37.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_37.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_35(.DOA({out_Q_i[22:22],out_Q_i[18:18]}),.DOB({vec_out_i_AQ_2[10:10],vec_out_i_AQ_2[6:6]}),.DOC(mat_i_1_I_35_DOC[1:0]),.DOD(mat_i_1_I_35_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_2[10:10],vec_in_i_AQ_mux_2[6:6]}),.DIB({vec_in_i_AQ_mux_2[10:10],vec_in_i_AQ_mux_2[6:6]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_35.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_35.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_35.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_35.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_33(.DOA({out_Q_i[36:36],out_Q_i[23:23]}),.DOB({vec_out_i_AQ_0[0:0],vec_out_i_AQ_2[11:11]}),.DOC(mat_i_1_I_33_DOC[1:0]),.DOD(mat_i_1_I_33_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_0,vec_in_i_AQ_mux_2[11:11]}),.DIB({vec_in_i_AQ_mux_0_0,vec_in_i_AQ_mux_2[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_33.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_33.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_33.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_33.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_31(.DOA({out_Q_i[10:10],out_Q_i[37:37]}),.DOB({vec_out_i_AQ_3[10:10],vec_out_i_AQ_0[1:1]}),.DOC(mat_i_1_I_31_DOC[1:0]),.DOD(mat_i_1_I_31_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[10:10],vec_in_i_AQ_mux_0_1}),.DIB({vec_in_i_AQ_mux_3[10:10],vec_in_i_AQ_mux_0_1}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_31.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_31.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_31.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_31.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_29(.DOA({out_Q_i[24:24],out_Q_i[11:11]}),.DOB({vec_out_i_AQ_1[0:0],vec_out_i_AQ_3[11:11]}),.DOC(mat_i_1_I_29_DOC[1:0]),.DOD(mat_i_1_I_29_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_1[0:0],vec_in_i_AQ_mux_3[11:11]}),.DIB({vec_in_i_AQ_mux_1[0:0],vec_in_i_AQ_mux_3[11:11]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_29.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_29.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_29.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_29.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_27(.DOA({out_Q_i[38:38],out_Q_i[25:25]}),.DOB({vec_out_i_AQ_0[2:2],vec_out_i_AQ_1[1:1]}),.DOC(mat_i_1_I_27_DOC[1:0]),.DOD(mat_i_1_I_27_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({N_505,vec_in_i_AQ_mux_1[1:1]}),.DIB({N_505,vec_in_i_AQ_mux_1[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_27.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_27.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_27.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_27.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_25(.DOA({out_Q_i[12:12],out_Q_i[39:39]}),.DOB({vec_out_i_AQ_2[0:0],vec_out_i_AQ_0[3:3]}),.DOC(mat_i_1_I_25_DOC[1:0]),.DOD(mat_i_1_I_25_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_2[0:0],N_506}),.DIB({vec_in_i_AQ_mux_2[0:0],N_506}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_25.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_25.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_25.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_25.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_23(.DOA({out_Q_i[9:9],out_Q_i[13:13]}),.DOB({vec_out_i_AQ_3[9:9],vec_out_i_AQ_2[1:1]}),.DOC(mat_i_1_I_23_DOC[1:0]),.DOD(mat_i_1_I_23_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[9:9],vec_in_i_AQ_mux_2[1:1]}),.DIB({vec_in_i_AQ_mux_3[9:9],vec_in_i_AQ_mux_2[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_23.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_23.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_23.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_23.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_21(.DOA({out_Q_i[40:40],out_Q_i[27:27]}),.DOB({vec_out_i_AQ_0[4:4],vec_out_i_AQ_1[3:3]}),.DOC(mat_i_1_I_21_DOC[1:0]),.DOD(mat_i_1_I_21_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_4,vec_in_i_AQ_mux_1[3:3]}),.DIB({vec_in_i_AQ_mux_0_4,vec_in_i_AQ_mux_1[3:3]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_21.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_21.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_21.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_21.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_19(.DOA({out_Q_i[14:14],out_Q_i[0:0]}),.DOB({vec_out_i_AQ_2[2:2],vec_out_i_AQ_3[0:0]}),.DOC(mat_i_1_I_19_DOC[1:0]),.DOD(mat_i_1_I_19_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_2[2:2],vec_in_i_AQ_mux_3[0:0]}),.DIB({vec_in_i_AQ_mux_2[2:2],vec_in_i_AQ_mux_3[0:0]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_19.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_19.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_19.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_19.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_17(.DOA({out_Q_i[6:6],out_Q_i[34:34]}),.DOB({vec_out_i_AQ_3[6:6],vec_out_i_AQ_1[10:10]}),.DOC(mat_i_1_I_17_DOC[1:0]),.DOD(mat_i_1_I_17_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[6:6],vec_in_i_AQ_mux_1[10:10]}),.DIB({vec_in_i_AQ_mux_3[6:6],vec_in_i_AQ_mux_1[10:10]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_17.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_17.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_17.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_17.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_15(.DOA({out_Q_i[42:42],out_Q_i[1:1]}),.DOB({vec_out_i_AQ_0[6:6],vec_out_i_AQ_3[1:1]}),.DOC(mat_i_1_I_15_DOC[1:0]),.DOD(mat_i_1_I_15_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_6,vec_in_i_AQ_mux_3[1:1]}),.DIB({vec_in_i_AQ_mux_0_6,vec_in_i_AQ_mux_3[1:1]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_15.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_15.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_15.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_15.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_13(.DOA({out_Q_i[7:7],out_Q_i[47:47]}),.DOB({vec_out_i_AQ_3[7:7],vec_out_i_AQ_0[11:11]}),.DOC(mat_i_1_I_13_DOC[1:0]),.DOD(mat_i_1_I_13_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[7:7],vec_in_i_AQ_mux_0_11}),.DIB({vec_in_i_AQ_mux_3[7:7],vec_in_i_AQ_mux_0_11}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_13.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_13.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_13.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_13.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_11(.DOA({out_Q_i[30:30],out_Q_i[17:17]}),.DOB({vec_out_i_AQ_1[6:6],vec_out_i_AQ_2[5:5]}),.DOC(mat_i_1_I_11_DOC[1:0]),.DOD(mat_i_1_I_11_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_1[6:6],vec_in_i_AQ_mux_2[5:5]}),.DIB({vec_in_i_AQ_mux_1[6:6],vec_in_i_AQ_mux_2[5:5]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_11.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_11.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_11.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_11.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_9(.DOA({out_Q_i[44:44],out_Q_i[31:31]}),.DOB({vec_out_i_AQ_0[8:8],vec_out_i_AQ_1[7:7]}),.DOC(mat_i_1_I_9_DOC[1:0]),.DOD(mat_i_1_I_9_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_0_8,vec_in_i_AQ_mux_1[7:7]}),.DIB({vec_in_i_AQ_mux_0_8,vec_in_i_AQ_mux_1[7:7]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_9.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_9.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_9.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_9.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_7(.DOA({out_Q_i[3:3],out_Q_i[45:45]}),.DOB({vec_out_i_AQ_3[3:3],vec_out_i_AQ_0[9:9]}),.DOC(mat_i_1_I_7_DOC[1:0]),.DOD(mat_i_1_I_7_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[3:3],vec_in_i_AQ_mux_0_9}),.DIB({vec_in_i_AQ_mux_3[3:3],vec_in_i_AQ_mux_0_9}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_7.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_7.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_7.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_7.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_5(.DOA({out_Q_i[4:4],out_Q_i[28:28]}),.DOB({vec_out_i_AQ_3[4:4],vec_out_i_AQ_1[4:4]}),.DOC(mat_i_1_I_5_DOC[1:0]),.DOD(mat_i_1_I_5_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_3[4:4],vec_in_i_AQ_mux_1[4:4]}),.DIB({vec_in_i_AQ_mux_3[4:4],vec_in_i_AQ_mux_1[4:4]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_5.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_5.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_5.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_5.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_3(.DOA({out_Q_i[15:15],out_Q_i[33:33]}),.DOB({vec_out_i_AQ_2[3:3],vec_out_i_AQ_1[9:9]}),.DOC(mat_i_1_I_3_DOC[1:0]),.DOD(mat_i_1_I_3_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_2[3:3],vec_in_i_AQ_mux_1[9:9]}),.DIB({vec_in_i_AQ_mux_2[3:3],vec_in_i_AQ_mux_1[9:9]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_3.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_3.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_3.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_3.INIT_D=64'h0000000000000000;
  RAM32M mat_i_1_I_1(.DOA({out_Q_i[29:29],out_Q_i[16:16]}),.DOB({vec_out_i_AQ_1[5:5],vec_out_i_AQ_2[4:4]}),.DOC(mat_i_1_I_1_DOC[1:0]),.DOD(mat_i_1_I_1_DOD[1:0]),.ADDRA({GND,GND,GND,col_sel_AQ2_mux_i_m3_lut6_2_O5,col_sel_AQ2_mux_i_m3_lut6_2_O6}),.ADDRB({GND,GND,GND,col_sel_AQ_int[1:0]}),.ADDRC({GND,GND,GND,GND,GND}),.ADDRD({GND,GND,GND,w_col_sel_AQ_mux_i_m3_lut6_2_O5,w_col_sel_AQ_mux_i_m3_lut6_2_O6}),.DIA({vec_in_i_AQ_mux_1[5:5],vec_in_i_AQ_mux_2[4:4]}),.DIB({vec_in_i_AQ_mux_1[5:5],vec_in_i_AQ_mux_2[4:4]}),.DIC({GND,GND}),.DID({GND,GND}),.WCLK(clk),.WE(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam mat_i_1_I_1.INIT_A=64'h0000000000000000;
defparam mat_i_1_I_1.INIT_B=64'h0000000000000000;
defparam mat_i_1_I_1.INIT_C=64'h0000000000000000;
defparam mat_i_1_I_1.INIT_D=64'h0000000000000000;
  LUT6 desc0(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[3:3]),.I3(out_Q_r[15:15]),.I4(out_Q_r[27:27]),.I5(out_Q_r[39:39]),.O(N_645));
defparam desc0.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc1(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[4:4]),.I3(out_Q_r[40:40]),.I4(out_Q_r[16:16]),.I5(out_Q_r[28:28]),.O(N_641));
defparam desc1.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc2(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[4:4]),.I3(vec_out_r_AQ_3[4:4]),.I4(vec_out_r_AQ_1[4:4]),.I5(vec_out_r_AQ_2[4:4]),.O(N_637));
defparam desc2.INIT=64'hFE76BA32DC549810;
  LUT6 desc3(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[11:11]),.I3(out_Q_r[23:23]),.I4(out_Q_r[35:35]),.I5(out_Q_r[47:47]),.O(N_632));
defparam desc3.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc4(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[5:5]),.I3(vec_out_i_AQ_1[5:5]),.I4(vec_out_i_AQ_2[5:5]),.I5(vec_out_i_AQ_3[5:5]),.O(N_628));
defparam desc4.INIT=64'hFEBADC9876325410;
  LUT6 desc5(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[11:11]),.I3(vec_out_r_AQ_1[11:11]),.I4(vec_out_r_AQ_2[11:11]),.I5(vec_out_r_AQ_3[11:11]),.O(N_624));
defparam desc5.INIT=64'hFEBADC9876325410;
  LUT6 desc6(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[7:7]),.I3(vec_out_r_AQ_3[7:7]),.I4(vec_out_r_AQ_1[7:7]),.I5(vec_out_r_AQ_2[7:7]),.O(N_623));
defparam desc6.INIT=64'hFE76BA32DC549810;
  LUT6 desc7(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[0:0]),.I3(vec_out_r_AQ_1[0:0]),.I4(vec_out_r_AQ_2[0:0]),.I5(vec_out_r_AQ_3[0:0]),.O(N_622));
defparam desc7.INIT=64'hFEBADC9876325410;
  LUT6 desc8(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[8:8]),.I3(out_Q_i[32:32]),.I4(out_Q_i[44:44]),.I5(out_Q_i[20:20]),.O(N_612));
defparam desc8.INIT=64'hF7B3E6A2D591C480;
  LUT6 desc9(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[10:10]),.I3(out_Q_r[22:22]),.I4(out_Q_r[46:46]),.I5(out_Q_r[34:34]),.O(N_607));
defparam desc9.INIT=64'hF7D5E6C4B391A280;
  LUT6 desc10(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[9:9]),.I3(out_Q_r[21:21]),.I4(out_Q_r[33:33]),.I5(out_Q_r[45:45]),.O(N_606));
defparam desc10.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc11(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[12:12]),.I3(out_Q_r[24:24]),.I4(out_Q_r[36:36]),.I5(out_Q_r[0:0]),.O(N_605));
defparam desc11.INIT=64'hFDB9ECA875316420;
  LUT6 desc12(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[10:10]),.I3(vec_out_r_AQ_2[10:10]),.I4(vec_out_r_AQ_3[10:10]),.I5(vec_out_r_AQ_1[10:10]),.O(N_597));
defparam desc12.INIT=64'hFEDC7654BA983210;
  LUT6 desc13(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_3[9:9]),.I3(vec_out_r_AQ_0[9:9]),.I4(vec_out_r_AQ_1[9:9]),.I5(vec_out_r_AQ_2[9:9]),.O(N_596));
defparam desc13.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc14(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[6:6]),.I3(vec_out_r_AQ_1[6:6]),.I4(vec_out_r_AQ_3[6:6]),.I5(vec_out_r_AQ_2[6:6]),.O(N_595));
defparam desc14.INIT=64'hFEBA7632DC985410;
  LUT6 desc15(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[10:10]),.I3(out_Q_i[22:22]),.I4(out_Q_i[46:46]),.I5(out_Q_i[34:34]),.O(N_586));
defparam desc15.INIT=64'hF7D5E6C4B391A280;
  LUT6 desc16(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[9:9]),.I3(out_Q_i[21:21]),.I4(out_Q_i[33:33]),.I5(out_Q_i[45:45]),.O(N_585));
defparam desc16.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc17(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[7:7]),.I3(out_Q_i[43:43]),.I4(out_Q_i[19:19]),.I5(out_Q_i[31:31]),.O(N_584));
defparam desc17.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc18(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[6:6]),.I3(out_Q_i[30:30]),.I4(out_Q_i[42:42]),.I5(out_Q_i[18:18]),.O(N_583));
defparam desc18.INIT=64'hF7B3E6A2D591C480;
  LUT6 desc19(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[3:3]),.I3(out_Q_i[15:15]),.I4(out_Q_i[27:27]),.I5(out_Q_i[39:39]),.O(N_582));
defparam desc19.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc20(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[6:6]),.I3(out_Q_r[30:30]),.I4(out_Q_r[42:42]),.I5(out_Q_r[18:18]),.O(N_571));
defparam desc20.INIT=64'hF7B3E6A2D591C480;
  LUT6 desc21(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[7:7]),.I3(vec_out_i_AQ_3[7:7]),.I4(vec_out_i_AQ_1[7:7]),.I5(vec_out_i_AQ_2[7:7]),.O(N_568));
defparam desc21.INIT=64'hFE76BA32DC549810;
  LUT6 desc22(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[6:6]),.I3(vec_out_i_AQ_1[6:6]),.I4(vec_out_i_AQ_3[6:6]),.I5(vec_out_i_AQ_2[6:6]),.O(N_567));
defparam desc22.INIT=64'hFEBA7632DC985410;
  LUT6 desc23(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_2[3:3]),.I3(vec_out_i_AQ_3[3:3]),.I4(vec_out_i_AQ_0[3:3]),.I5(vec_out_i_AQ_1[3:3]),.O(N_566));
defparam desc23.INIT=64'hFD75EC64B931A820;
  LUT6 desc24(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[14:14]),.I3(out_Q_i[26:26]),.I4(out_Q_i[38:38]),.I5(out_Q_i[2:2]),.O(N_555));
defparam desc24.INIT=64'hFDB9ECA875316420;
  LUT6 desc25(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[8:8]),.I3(out_Q_r[32:32]),.I4(out_Q_r[44:44]),.I5(out_Q_r[20:20]),.O(N_552));
defparam desc25.INIT=64'hF7B3E6A2D591C480;
  LUT6 desc26(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[2:2]),.I3(vec_out_i_AQ_1[2:2]),.I4(vec_out_i_AQ_2[2:2]),.I5(vec_out_i_AQ_3[2:2]),.O(N_549));
defparam desc26.INIT=64'hFEBADC9876325410;
  LUT6 desc27(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[14:14]),.I3(out_Q_r[26:26]),.I4(out_Q_r[38:38]),.I5(out_Q_r[2:2]),.O(single_out_r_AQ2_1));
defparam desc27.INIT=64'hFDB9ECA875316420;
  LUT6 desc28(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[5:5]),.I3(vec_out_r_AQ_1[5:5]),.I4(vec_out_r_AQ_2[5:5]),.I5(vec_out_r_AQ_3[5:5]),.O(single_out_r_AQ_4));
defparam desc28.INIT=64'hFEBADC9876325410;
  LUT6 desc29(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_2[3:3]),.I3(vec_out_r_AQ_3[3:3]),.I4(vec_out_r_AQ_0[3:3]),.I5(vec_out_r_AQ_1[3:3]),.O(single_out_r_AQ_2));
defparam desc29.INIT=64'hFD75EC64B931A820;
  LUT6 desc30(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[1:1]),.I3(out_Q_i[13:13]),.I4(out_Q_i[25:25]),.I5(out_Q_i[37:37]),.O(single_out_i_AQ2_1));
defparam desc30.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc31(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[1:1]),.I3(vec_out_i_AQ_1[1:1]),.I4(vec_out_i_AQ_2[1:1]),.I5(vec_out_i_AQ_3[1:1]),.O(single_out_i_AQ_1));
defparam desc31.INIT=64'hFEBADC9876325410;
  LUT6 desc32(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[29:29]),.I3(out_Q_i[41:41]),.I4(out_Q_i[5:5]),.I5(out_Q_i[17:17]),.O(single_out_i_AQ2_5));
defparam desc32.INIT=64'hFBEA7362D9C85140;
  LUT6 desc33(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[7:7]),.I3(out_Q_r[43:43]),.I4(out_Q_r[19:19]),.I5(out_Q_r[31:31]),.O(single_out_r_AQ2_6));
defparam desc33.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc34(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[0:0]),.I3(vec_out_i_AQ_1[0:0]),.I4(vec_out_i_AQ_2[0:0]),.I5(vec_out_i_AQ_3[0:0]),.O(single_out_i_AQ_0));
defparam desc34.INIT=64'hFEBADC9876325410;
  LUT6 desc35(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[4:4]),.I3(out_Q_i[40:40]),.I4(out_Q_i[16:16]),.I5(out_Q_i[28:28]),.O(single_out_i_AQ2_4));
defparam desc35.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc36(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[12:12]),.I3(out_Q_i[24:24]),.I4(out_Q_i[36:36]),.I5(out_Q_i[0:0]),.O(single_out_i_AQ2_0));
defparam desc36.INIT=64'hFDB9ECA875316420;
  LUT6 desc37(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[29:29]),.I3(out_Q_r[41:41]),.I4(out_Q_r[5:5]),.I5(out_Q_r[17:17]),.O(single_out_r_AQ2_4));
defparam desc37.INIT=64'hFBEA7362D9C85140;
  LUT6 desc38(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_r[1:1]),.I3(out_Q_r[13:13]),.I4(out_Q_r[25:25]),.I5(out_Q_r[37:37]),.O(single_out_r_AQ2_0));
defparam desc38.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc39(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[8:8]),.I3(vec_out_i_AQ_1[8:8]),.I4(vec_out_i_AQ_3[8:8]),.I5(vec_out_i_AQ_2[8:8]),.O(single_out_i_AQ_8));
defparam desc39.INIT=64'hFEBA7632DC985410;
  LUT6 desc40(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[10:10]),.I3(vec_out_i_AQ_2[10:10]),.I4(vec_out_i_AQ_3[10:10]),.I5(vec_out_i_AQ_1[10:10]),.O(single_out_i_AQ_10));
defparam desc40.INIT=64'hFEDC7654BA983210;
  LUT6 desc41(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(out_Q_i[11:11]),.I3(out_Q_i[23:23]),.I4(out_Q_i[35:35]),.I5(out_Q_i[47:47]),.O(single_out_i_AQ2_11));
defparam desc41.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc42(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[11:11]),.I3(vec_out_i_AQ_1[11:11]),.I4(vec_out_i_AQ_2[11:11]),.I5(vec_out_i_AQ_3[11:11]),.O(single_out_i_AQ_11));
defparam desc42.INIT=64'hFEBADC9876325410;
  LUT6 desc43(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_3[9:9]),.I3(vec_out_i_AQ_0[9:9]),.I4(vec_out_i_AQ_1[9:9]),.I5(vec_out_i_AQ_2[9:9]),.O(single_out_i_AQ_9));
defparam desc43.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc44(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_i_AQ_0[4:4]),.I3(vec_out_i_AQ_3[4:4]),.I4(vec_out_i_AQ_1[4:4]),.I5(vec_out_i_AQ_2[4:4]),.O(single_out_i_AQ_4));
defparam desc44.INIT=64'hFE76BA32DC549810;
  LUT6 desc45(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[8:8]),.I3(vec_out_r_AQ_1[8:8]),.I4(vec_out_r_AQ_3[8:8]),.I5(vec_out_r_AQ_2[8:8]),.O(single_out_r_AQ_7));
defparam desc45.INIT=64'hFEBA7632DC985410;
  LUT6 desc46(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[2:2]),.I3(vec_out_r_AQ_1[2:2]),.I4(vec_out_r_AQ_2[2:2]),.I5(vec_out_r_AQ_3[2:2]),.O(single_out_r_AQ_1));
defparam desc46.INIT=64'hFEBADC9876325410;
  LUT6 desc47(.I0(row_sel_AQ[1:1]),.I1(row_sel_AQ[0:0]),.I2(vec_out_r_AQ_0[1:1]),.I3(vec_out_r_AQ_1[1:1]),.I4(vec_out_r_AQ_2[1:1]),.I5(vec_out_r_AQ_3[1:1]),.O(single_out_r_AQ_0));
defparam desc47.INIT=64'hFEBADC9876325410;
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
endmodule
module mult_pipe_inj (mult1_out,in_a_r_reg,in_b_r_reg,clk);
output [23:23] mult1_out ;
input [11:0] in_a_r_reg ;
input [11:0] in_b_r_reg ;
input clk ;
wire clk ;
wire [29:0] ACOUT_33 ;
wire [17:0] BCOUT_33 ;
wire [3:0] CARRYOUT_33 ;
wire [22:0] pre_out_P_0 ;
wire [47:24] P_uc_33 ;
wire [47:0] PCOUT_33 ;
wire CARRYCASCOUT_33 ;
wire MULTSIGNOUT_33 ;
wire OVERFLOW_33 ;
wire PATTERNBDETECT_33 ;
wire PATTERNDETECT_33 ;
wire UNDERFLOW_33 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc264(.ACOUT(ACOUT_33[29:0]),.BCOUT(BCOUT_33[17:0]),.CARRYCASCOUT(CARRYCASCOUT_33),.CARRYOUT(CARRYOUT_33[3:0]),.MULTSIGNOUT(MULTSIGNOUT_33),.OVERFLOW(OVERFLOW_33),.P({P_uc_33[47:24],mult1_out[23:23],pre_out_P_0[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_33),.PATTERNDETECT(PATTERNDETECT_33),.PCOUT(PCOUT_33[47:0]),.UNDERFLOW(UNDERFLOW_33),.A({in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(VCC),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc264.ACASCREG=0;
defparam desc264.ADREG=0;
defparam desc264.ALUMODEREG=0;
defparam desc264.AREG=0;
defparam desc264.AUTORESET_PATDET="NO_RESET";
defparam desc264.A_INPUT="DIRECT";
defparam desc264.BCASCREG=0;
defparam desc264.BREG=0;
defparam desc264.B_INPUT="DIRECT";
defparam desc264.CARRYINREG=0;
defparam desc264.CARRYINSELREG=0;
defparam desc264.CREG=1;
defparam desc264.DREG=0;
defparam desc264.INMODEREG=0;
defparam desc264.MREG=1;
defparam desc264.OPMODEREG=0;
defparam desc264.PREG=0;
defparam desc264.USE_DPORT="FALSE";
defparam desc264.USE_MULT="MULTIPLY";
defparam desc264.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_1_inj (mult2_out_23,mult2_out_0,P_uc_34_0,in_a_i_reg,in_b_i_reg,clk);
output mult2_out_23 ;
output [23:0] mult2_out_0 ;
output [47:24] P_uc_34_0 ;
input [11:0] in_a_i_reg ;
input [11:0] in_b_i_reg ;
input clk ;
wire mult2_out_23 ;
wire clk ;
wire [29:0] ACOUT_34 ;
wire [17:0] BCOUT_34 ;
wire [3:0] CARRYOUT_34 ;
wire [22:0] mult2_out ;
wire [47:24] P_uc_34 ;
wire CARRYCASCOUT_34 ;
wire MULTSIGNOUT_34 ;
wire OVERFLOW_34 ;
wire PATTERNBDETECT_34 ;
wire PATTERNDETECT_34 ;
wire UNDERFLOW_34 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc265(.ACOUT(ACOUT_34[29:0]),.BCOUT(BCOUT_34[17:0]),.CARRYCASCOUT(CARRYCASCOUT_34),.CARRYOUT(CARRYOUT_34[3:0]),.MULTSIGNOUT(MULTSIGNOUT_34),.OVERFLOW(OVERFLOW_34),.P({P_uc_34[47:24],mult2_out_23,mult2_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_34),.PATTERNDETECT(PATTERNDETECT_34),.PCOUT({P_uc_34_0[47:24],mult2_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_34),.A({in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc265.ACASCREG=0;
defparam desc265.ADREG=0;
defparam desc265.ALUMODEREG=0;
defparam desc265.AREG=0;
defparam desc265.AUTORESET_PATDET="NO_RESET";
defparam desc265.A_INPUT="DIRECT";
defparam desc265.BCASCREG=0;
defparam desc265.BREG=0;
defparam desc265.B_INPUT="DIRECT";
defparam desc265.CARRYINREG=0;
defparam desc265.CARRYINSELREG=0;
defparam desc265.CREG=1;
defparam desc265.DREG=0;
defparam desc265.INMODEREG=0;
defparam desc265.MREG=0;
defparam desc265.OPMODEREG=0;
defparam desc265.PREG=1;
defparam desc265.USE_DPORT="FALSE";
defparam desc265.USE_MULT="MULTIPLY";
defparam desc265.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_10_inj (mult3_out_23,vec_out_r_AQ_1,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult3_out_23 ;
input [11:0] vec_out_r_AQ_1 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult3_out_23 ;
wire clk ;
wire [29:0] ACOUT_22 ;
wire [17:0] BCOUT_22 ;
wire [3:0] CARRYOUT_22 ;
wire [22:0] mult3_out ;
wire [47:24] P_uc_22 ;
wire [47:0] PCOUT_22 ;
wire CARRYCASCOUT_22 ;
wire MULTSIGNOUT_22 ;
wire OVERFLOW_22 ;
wire PATTERNBDETECT_22 ;
wire PATTERNDETECT_22 ;
wire UNDERFLOW_22 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc532(.ACOUT(ACOUT_22[29:0]),.BCOUT(BCOUT_22[17:0]),.CARRYCASCOUT(CARRYCASCOUT_22),.CARRYOUT(CARRYOUT_22[3:0]),.MULTSIGNOUT(MULTSIGNOUT_22),.OVERFLOW(OVERFLOW_22),.P({P_uc_22[47:24],mult3_out_23,mult3_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_22),.PATTERNDETECT(PATTERNDETECT_22),.PCOUT(PCOUT_22[47:0]),.UNDERFLOW(UNDERFLOW_22),.A({vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc532.ACASCREG=1;
defparam desc532.ADREG=0;
defparam desc532.ALUMODEREG=0;
defparam desc532.AREG=1;
defparam desc532.AUTORESET_PATDET="NO_RESET";
defparam desc532.A_INPUT="DIRECT";
defparam desc532.BCASCREG=1;
defparam desc532.BREG=1;
defparam desc532.B_INPUT="DIRECT";
defparam desc532.CARRYINREG=0;
defparam desc532.CARRYINSELREG=0;
defparam desc532.CREG=1;
defparam desc532.DREG=0;
defparam desc532.INMODEREG=0;
defparam desc532.MREG=0;
defparam desc532.OPMODEREG=0;
defparam desc532.PREG=1;
defparam desc532.USE_DPORT="FALSE";
defparam desc532.USE_MULT="MULTIPLY";
defparam desc532.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_11_inj (mult4_out_23,mult4_out_0,P_uc_23_0,out_inner_prod_r,vec_out_i_AQ_1,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult4_out_23 ;
output [23:0] mult4_out_0 ;
output [47:24] P_uc_23_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_i_AQ_1 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult4_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_23 ;
wire [17:0] BCOUT_23 ;
wire [3:0] CARRYOUT_23 ;
wire [22:0] mult4_out ;
wire [47:24] P_uc_23 ;
wire CARRYCASCOUT_23 ;
wire MULTSIGNOUT_23 ;
wire OVERFLOW_23 ;
wire PATTERNBDETECT_23 ;
wire PATTERNDETECT_23 ;
wire UNDERFLOW_23 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc533(.ACOUT(ACOUT_23[29:0]),.BCOUT(BCOUT_23[17:0]),.CARRYCASCOUT(CARRYCASCOUT_23),.CARRYOUT(CARRYOUT_23[3:0]),.MULTSIGNOUT(MULTSIGNOUT_23),.OVERFLOW(OVERFLOW_23),.P({P_uc_23[47:24],mult4_out_23,mult4_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_23),.PATTERNDETECT(PATTERNDETECT_23),.PCOUT({P_uc_23_0[47:24],mult4_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_23),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc533.ACASCREG=1;
defparam desc533.ADREG=1;
defparam desc533.ALUMODEREG=0;
defparam desc533.AREG=1;
defparam desc533.AUTORESET_PATDET="NO_RESET";
defparam desc533.A_INPUT="DIRECT";
defparam desc533.BCASCREG=2;
defparam desc533.BREG=2;
defparam desc533.B_INPUT="DIRECT";
defparam desc533.CARRYINREG=0;
defparam desc533.CARRYINSELREG=0;
defparam desc533.CREG=1;
defparam desc533.DREG=1;
defparam desc533.INMODEREG=1;
defparam desc533.MREG=0;
defparam desc533.OPMODEREG=0;
defparam desc533.PREG=0;
defparam desc533.USE_DPORT="TRUE";
defparam desc533.USE_MULT="MULTIPLY";
defparam desc533.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_12_inj (mult1_out_23,mult1_out_0,P_uc_16_0,out_inner_prod_r,vec_out_r_AQ_0,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult1_out_23 ;
output [23:0] mult1_out_0 ;
output [47:24] P_uc_16_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_0 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult1_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_16 ;
wire [17:0] BCOUT_16 ;
wire [3:0] CARRYOUT_16 ;
wire [22:0] mult1_out ;
wire [47:24] P_uc_16 ;
wire CARRYCASCOUT_16 ;
wire MULTSIGNOUT_16 ;
wire OVERFLOW_16 ;
wire PATTERNBDETECT_16 ;
wire PATTERNDETECT_16 ;
wire UNDERFLOW_16 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc585(.ACOUT(ACOUT_16[29:0]),.BCOUT(BCOUT_16[17:0]),.CARRYCASCOUT(CARRYCASCOUT_16),.CARRYOUT(CARRYOUT_16[3:0]),.MULTSIGNOUT(MULTSIGNOUT_16),.OVERFLOW(OVERFLOW_16),.P({P_uc_16[47:24],mult1_out_23,mult1_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_16),.PATTERNDETECT(PATTERNDETECT_16),.PCOUT({P_uc_16_0[47:24],mult1_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_16),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc585.ACASCREG=1;
defparam desc585.ADREG=1;
defparam desc585.ALUMODEREG=0;
defparam desc585.AREG=1;
defparam desc585.AUTORESET_PATDET="NO_RESET";
defparam desc585.A_INPUT="DIRECT";
defparam desc585.BCASCREG=2;
defparam desc585.BREG=2;
defparam desc585.B_INPUT="DIRECT";
defparam desc585.CARRYINREG=0;
defparam desc585.CARRYINSELREG=0;
defparam desc585.CREG=1;
defparam desc585.DREG=1;
defparam desc585.INMODEREG=1;
defparam desc585.MREG=0;
defparam desc585.OPMODEREG=0;
defparam desc585.PREG=0;
defparam desc585.USE_DPORT="TRUE";
defparam desc585.USE_MULT="MULTIPLY";
defparam desc585.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_13_inj (mult2_out_23,vec_out_i_AQ_0,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult2_out_23 ;
input [11:0] vec_out_i_AQ_0 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult2_out_23 ;
wire clk ;
wire [29:0] ACOUT_17 ;
wire [17:0] BCOUT_17 ;
wire [3:0] CARRYOUT_17 ;
wire [22:0] mult2_out ;
wire [47:24] P_uc_17 ;
wire [47:0] PCOUT_17 ;
wire CARRYCASCOUT_17 ;
wire MULTSIGNOUT_17 ;
wire OVERFLOW_17 ;
wire PATTERNBDETECT_17 ;
wire PATTERNDETECT_17 ;
wire UNDERFLOW_17 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc586(.ACOUT(ACOUT_17[29:0]),.BCOUT(BCOUT_17[17:0]),.CARRYCASCOUT(CARRYCASCOUT_17),.CARRYOUT(CARRYOUT_17[3:0]),.MULTSIGNOUT(MULTSIGNOUT_17),.OVERFLOW(OVERFLOW_17),.P({P_uc_17[47:24],mult2_out_23,mult2_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_17),.PATTERNDETECT(PATTERNDETECT_17),.PCOUT(PCOUT_17[47:0]),.UNDERFLOW(UNDERFLOW_17),.A({vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc586.ACASCREG=1;
defparam desc586.ADREG=0;
defparam desc586.ALUMODEREG=0;
defparam desc586.AREG=1;
defparam desc586.AUTORESET_PATDET="NO_RESET";
defparam desc586.A_INPUT="DIRECT";
defparam desc586.BCASCREG=1;
defparam desc586.BREG=1;
defparam desc586.B_INPUT="DIRECT";
defparam desc586.CARRYINREG=0;
defparam desc586.CARRYINSELREG=0;
defparam desc586.CREG=1;
defparam desc586.DREG=0;
defparam desc586.INMODEREG=0;
defparam desc586.MREG=0;
defparam desc586.OPMODEREG=0;
defparam desc586.PREG=1;
defparam desc586.USE_DPORT="FALSE";
defparam desc586.USE_MULT="MULTIPLY";
defparam desc586.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_14_inj (mult3_out_23,vec_out_r_AQ_0,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult3_out_23 ;
input [11:0] vec_out_r_AQ_0 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult3_out_23 ;
wire clk ;
wire [29:0] ACOUT_18 ;
wire [17:0] BCOUT_18 ;
wire [3:0] CARRYOUT_18 ;
wire [22:0] mult3_out ;
wire [47:24] P_uc_18 ;
wire [47:0] PCOUT_18 ;
wire CARRYCASCOUT_18 ;
wire MULTSIGNOUT_18 ;
wire OVERFLOW_18 ;
wire PATTERNBDETECT_18 ;
wire PATTERNDETECT_18 ;
wire UNDERFLOW_18 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc587(.ACOUT(ACOUT_18[29:0]),.BCOUT(BCOUT_18[17:0]),.CARRYCASCOUT(CARRYCASCOUT_18),.CARRYOUT(CARRYOUT_18[3:0]),.MULTSIGNOUT(MULTSIGNOUT_18),.OVERFLOW(OVERFLOW_18),.P({P_uc_18[47:24],mult3_out_23,mult3_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_18),.PATTERNDETECT(PATTERNDETECT_18),.PCOUT(PCOUT_18[47:0]),.UNDERFLOW(UNDERFLOW_18),.A({vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:11],vec_out_r_AQ_0[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc587.ACASCREG=1;
defparam desc587.ADREG=0;
defparam desc587.ALUMODEREG=0;
defparam desc587.AREG=1;
defparam desc587.AUTORESET_PATDET="NO_RESET";
defparam desc587.A_INPUT="DIRECT";
defparam desc587.BCASCREG=1;
defparam desc587.BREG=1;
defparam desc587.B_INPUT="DIRECT";
defparam desc587.CARRYINREG=0;
defparam desc587.CARRYINSELREG=0;
defparam desc587.CREG=1;
defparam desc587.DREG=0;
defparam desc587.INMODEREG=0;
defparam desc587.MREG=0;
defparam desc587.OPMODEREG=0;
defparam desc587.PREG=1;
defparam desc587.USE_DPORT="FALSE";
defparam desc587.USE_MULT="MULTIPLY";
defparam desc587.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_15_inj (mult4_out_23,mult4_out_0,P_uc_19_0,out_inner_prod_r,vec_out_i_AQ_0,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult4_out_23 ;
output [23:0] mult4_out_0 ;
output [47:24] P_uc_19_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_i_AQ_0 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult4_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_19 ;
wire [17:0] BCOUT_19 ;
wire [3:0] CARRYOUT_19 ;
wire [22:0] mult4_out ;
wire [47:24] P_uc_19 ;
wire CARRYCASCOUT_19 ;
wire MULTSIGNOUT_19 ;
wire OVERFLOW_19 ;
wire PATTERNBDETECT_19 ;
wire PATTERNDETECT_19 ;
wire UNDERFLOW_19 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc588(.ACOUT(ACOUT_19[29:0]),.BCOUT(BCOUT_19[17:0]),.CARRYCASCOUT(CARRYCASCOUT_19),.CARRYOUT(CARRYOUT_19[3:0]),.MULTSIGNOUT(MULTSIGNOUT_19),.OVERFLOW(OVERFLOW_19),.P({P_uc_19[47:24],mult4_out_23,mult4_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_19),.PATTERNDETECT(PATTERNDETECT_19),.PCOUT({P_uc_19_0[47:24],mult4_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_19),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:11],vec_out_i_AQ_0[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc588.ACASCREG=1;
defparam desc588.ADREG=1;
defparam desc588.ALUMODEREG=0;
defparam desc588.AREG=1;
defparam desc588.AUTORESET_PATDET="NO_RESET";
defparam desc588.A_INPUT="DIRECT";
defparam desc588.BCASCREG=2;
defparam desc588.BREG=2;
defparam desc588.B_INPUT="DIRECT";
defparam desc588.CARRYINREG=0;
defparam desc588.CARRYINSELREG=0;
defparam desc588.CREG=1;
defparam desc588.DREG=1;
defparam desc588.INMODEREG=1;
defparam desc588.MREG=0;
defparam desc588.OPMODEREG=0;
defparam desc588.PREG=0;
defparam desc588.USE_DPORT="TRUE";
defparam desc588.USE_MULT="MULTIPLY";
defparam desc588.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_16_inj (mult1_out_23,mult1_out_0,P_uc_28_0,out_inner_prod_r,vec_out_r_AQ_3,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult1_out_23 ;
output [23:0] mult1_out_0 ;
output [47:24] P_uc_28_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_3 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult1_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_28 ;
wire [17:0] BCOUT_28 ;
wire [3:0] CARRYOUT_28 ;
wire [22:0] mult1_out ;
wire [47:24] P_uc_28 ;
wire CARRYCASCOUT_28 ;
wire MULTSIGNOUT_28 ;
wire OVERFLOW_28 ;
wire PATTERNBDETECT_28 ;
wire PATTERNDETECT_28 ;
wire UNDERFLOW_28 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc640(.ACOUT(ACOUT_28[29:0]),.BCOUT(BCOUT_28[17:0]),.CARRYCASCOUT(CARRYCASCOUT_28),.CARRYOUT(CARRYOUT_28[3:0]),.MULTSIGNOUT(MULTSIGNOUT_28),.OVERFLOW(OVERFLOW_28),.P({P_uc_28[47:24],mult1_out_23,mult1_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_28),.PATTERNDETECT(PATTERNDETECT_28),.PCOUT({P_uc_28_0[47:24],mult1_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_28),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc640.ACASCREG=1;
defparam desc640.ADREG=1;
defparam desc640.ALUMODEREG=0;
defparam desc640.AREG=1;
defparam desc640.AUTORESET_PATDET="NO_RESET";
defparam desc640.A_INPUT="DIRECT";
defparam desc640.BCASCREG=2;
defparam desc640.BREG=2;
defparam desc640.B_INPUT="DIRECT";
defparam desc640.CARRYINREG=0;
defparam desc640.CARRYINSELREG=0;
defparam desc640.CREG=1;
defparam desc640.DREG=1;
defparam desc640.INMODEREG=1;
defparam desc640.MREG=0;
defparam desc640.OPMODEREG=0;
defparam desc640.PREG=0;
defparam desc640.USE_DPORT="TRUE";
defparam desc640.USE_MULT="MULTIPLY";
defparam desc640.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_17_inj (mult2_out_23,vec_out_i_AQ_3,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult2_out_23 ;
input [11:0] vec_out_i_AQ_3 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult2_out_23 ;
wire clk ;
wire [29:0] ACOUT_29 ;
wire [17:0] BCOUT_29 ;
wire [3:0] CARRYOUT_29 ;
wire [22:0] mult2_out ;
wire [47:24] P_uc_29 ;
wire [47:0] PCOUT_29 ;
wire CARRYCASCOUT_29 ;
wire MULTSIGNOUT_29 ;
wire OVERFLOW_29 ;
wire PATTERNBDETECT_29 ;
wire PATTERNDETECT_29 ;
wire UNDERFLOW_29 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc641(.ACOUT(ACOUT_29[29:0]),.BCOUT(BCOUT_29[17:0]),.CARRYCASCOUT(CARRYCASCOUT_29),.CARRYOUT(CARRYOUT_29[3:0]),.MULTSIGNOUT(MULTSIGNOUT_29),.OVERFLOW(OVERFLOW_29),.P({P_uc_29[47:24],mult2_out_23,mult2_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_29),.PATTERNDETECT(PATTERNDETECT_29),.PCOUT(PCOUT_29[47:0]),.UNDERFLOW(UNDERFLOW_29),.A({vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc641.ACASCREG=1;
defparam desc641.ADREG=0;
defparam desc641.ALUMODEREG=0;
defparam desc641.AREG=1;
defparam desc641.AUTORESET_PATDET="NO_RESET";
defparam desc641.A_INPUT="DIRECT";
defparam desc641.BCASCREG=1;
defparam desc641.BREG=1;
defparam desc641.B_INPUT="DIRECT";
defparam desc641.CARRYINREG=0;
defparam desc641.CARRYINSELREG=0;
defparam desc641.CREG=1;
defparam desc641.DREG=0;
defparam desc641.INMODEREG=0;
defparam desc641.MREG=0;
defparam desc641.OPMODEREG=0;
defparam desc641.PREG=1;
defparam desc641.USE_DPORT="FALSE";
defparam desc641.USE_MULT="MULTIPLY";
defparam desc641.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_18_inj (mult3_out_23,vec_out_r_AQ_3,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult3_out_23 ;
input [11:0] vec_out_r_AQ_3 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult3_out_23 ;
wire clk ;
wire [29:0] ACOUT_30 ;
wire [17:0] BCOUT_30 ;
wire [3:0] CARRYOUT_30 ;
wire [22:0] mult3_out ;
wire [47:24] P_uc_30 ;
wire [47:0] PCOUT_30 ;
wire CARRYCASCOUT_30 ;
wire MULTSIGNOUT_30 ;
wire OVERFLOW_30 ;
wire PATTERNBDETECT_30 ;
wire PATTERNDETECT_30 ;
wire UNDERFLOW_30 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc642(.ACOUT(ACOUT_30[29:0]),.BCOUT(BCOUT_30[17:0]),.CARRYCASCOUT(CARRYCASCOUT_30),.CARRYOUT(CARRYOUT_30[3:0]),.MULTSIGNOUT(MULTSIGNOUT_30),.OVERFLOW(OVERFLOW_30),.P({P_uc_30[47:24],mult3_out_23,mult3_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_30),.PATTERNDETECT(PATTERNDETECT_30),.PCOUT(PCOUT_30[47:0]),.UNDERFLOW(UNDERFLOW_30),.A({vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:11],vec_out_r_AQ_3[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc642.ACASCREG=1;
defparam desc642.ADREG=0;
defparam desc642.ALUMODEREG=0;
defparam desc642.AREG=1;
defparam desc642.AUTORESET_PATDET="NO_RESET";
defparam desc642.A_INPUT="DIRECT";
defparam desc642.BCASCREG=1;
defparam desc642.BREG=1;
defparam desc642.B_INPUT="DIRECT";
defparam desc642.CARRYINREG=0;
defparam desc642.CARRYINSELREG=0;
defparam desc642.CREG=1;
defparam desc642.DREG=0;
defparam desc642.INMODEREG=0;
defparam desc642.MREG=0;
defparam desc642.OPMODEREG=0;
defparam desc642.PREG=1;
defparam desc642.USE_DPORT="FALSE";
defparam desc642.USE_MULT="MULTIPLY";
defparam desc642.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_19_inj (mult4_out_23,mult4_out_0,P_uc_31_0,out_inner_prod_r,vec_out_i_AQ_3,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult4_out_23 ;
output [23:0] mult4_out_0 ;
output [47:24] P_uc_31_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_i_AQ_3 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult4_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_31 ;
wire [17:0] BCOUT_31 ;
wire [3:0] CARRYOUT_31 ;
wire [22:0] mult4_out ;
wire [47:24] P_uc_31 ;
wire CARRYCASCOUT_31 ;
wire MULTSIGNOUT_31 ;
wire OVERFLOW_31 ;
wire PATTERNBDETECT_31 ;
wire PATTERNDETECT_31 ;
wire UNDERFLOW_31 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc643(.ACOUT(ACOUT_31[29:0]),.BCOUT(BCOUT_31[17:0]),.CARRYCASCOUT(CARRYCASCOUT_31),.CARRYOUT(CARRYOUT_31[3:0]),.MULTSIGNOUT(MULTSIGNOUT_31),.OVERFLOW(OVERFLOW_31),.P({P_uc_31[47:24],mult4_out_23,mult4_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_31),.PATTERNDETECT(PATTERNDETECT_31),.PCOUT({P_uc_31_0[47:24],mult4_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_31),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:11],vec_out_i_AQ_3[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc643.ACASCREG=1;
defparam desc643.ADREG=1;
defparam desc643.ALUMODEREG=0;
defparam desc643.AREG=1;
defparam desc643.AUTORESET_PATDET="NO_RESET";
defparam desc643.A_INPUT="DIRECT";
defparam desc643.BCASCREG=2;
defparam desc643.BREG=2;
defparam desc643.B_INPUT="DIRECT";
defparam desc643.CARRYINREG=0;
defparam desc643.CARRYINSELREG=0;
defparam desc643.CREG=1;
defparam desc643.DREG=1;
defparam desc643.INMODEREG=1;
defparam desc643.MREG=0;
defparam desc643.OPMODEREG=0;
defparam desc643.PREG=0;
defparam desc643.USE_DPORT="TRUE";
defparam desc643.USE_MULT="MULTIPLY";
defparam desc643.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_2_inj (mult3_out_23,mult3_out_0,P_uc_35_0,in_a_r_reg,in_b_i_reg,clk);
output mult3_out_23 ;
output [23:0] mult3_out_0 ;
output [47:24] P_uc_35_0 ;
input [11:0] in_a_r_reg ;
input [11:0] in_b_i_reg ;
input clk ;
wire mult3_out_23 ;
wire clk ;
wire [29:0] ACOUT_35 ;
wire [17:0] BCOUT_35 ;
wire [3:0] CARRYOUT_35 ;
wire [22:0] mult3_out ;
wire [47:24] P_uc_35 ;
wire CARRYCASCOUT_35 ;
wire MULTSIGNOUT_35 ;
wire OVERFLOW_35 ;
wire PATTERNBDETECT_35 ;
wire PATTERNDETECT_35 ;
wire UNDERFLOW_35 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc266(.ACOUT(ACOUT_35[29:0]),.BCOUT(BCOUT_35[17:0]),.CARRYCASCOUT(CARRYCASCOUT_35),.CARRYOUT(CARRYOUT_35[3:0]),.MULTSIGNOUT(MULTSIGNOUT_35),.OVERFLOW(OVERFLOW_35),.P({P_uc_35[47:24],mult3_out_23,mult3_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_35),.PATTERNDETECT(PATTERNDETECT_35),.PCOUT({P_uc_35_0[47:24],mult3_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_35),.A({in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:11],in_a_r_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:11],in_b_i_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc266.ACASCREG=0;
defparam desc266.ADREG=0;
defparam desc266.ALUMODEREG=0;
defparam desc266.AREG=0;
defparam desc266.AUTORESET_PATDET="NO_RESET";
defparam desc266.A_INPUT="DIRECT";
defparam desc266.BCASCREG=0;
defparam desc266.BREG=0;
defparam desc266.B_INPUT="DIRECT";
defparam desc266.CARRYINREG=0;
defparam desc266.CARRYINSELREG=0;
defparam desc266.CREG=1;
defparam desc266.DREG=0;
defparam desc266.INMODEREG=0;
defparam desc266.MREG=0;
defparam desc266.OPMODEREG=0;
defparam desc266.PREG=1;
defparam desc266.USE_DPORT="FALSE";
defparam desc266.USE_MULT="MULTIPLY";
defparam desc266.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_3_inj (mult4_out,in_a_i_reg,in_b_r_reg,clk);
output [23:23] mult4_out ;
input [11:0] in_a_i_reg ;
input [11:0] in_b_r_reg ;
input clk ;
wire clk ;
wire [29:0] ACOUT_36 ;
wire [17:0] BCOUT_36 ;
wire [3:0] CARRYOUT_36 ;
wire [22:0] pre_out_P ;
wire [47:24] P_uc_36 ;
wire [47:0] PCOUT_36 ;
wire CARRYCASCOUT_36 ;
wire MULTSIGNOUT_36 ;
wire OVERFLOW_36 ;
wire PATTERNBDETECT_36 ;
wire PATTERNDETECT_36 ;
wire UNDERFLOW_36 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc267(.ACOUT(ACOUT_36[29:0]),.BCOUT(BCOUT_36[17:0]),.CARRYCASCOUT(CARRYCASCOUT_36),.CARRYOUT(CARRYOUT_36[3:0]),.MULTSIGNOUT(MULTSIGNOUT_36),.OVERFLOW(OVERFLOW_36),.P({P_uc_36[47:24],mult4_out[23:23],pre_out_P[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_36),.PATTERNDETECT(PATTERNDETECT_36),.PCOUT(PCOUT_36[47:0]),.UNDERFLOW(UNDERFLOW_36),.A({in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:11],in_a_i_reg[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:11],in_b_r_reg[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(VCC),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc267.ACASCREG=0;
defparam desc267.ADREG=0;
defparam desc267.ALUMODEREG=0;
defparam desc267.AREG=0;
defparam desc267.AUTORESET_PATDET="NO_RESET";
defparam desc267.A_INPUT="DIRECT";
defparam desc267.BCASCREG=0;
defparam desc267.BREG=0;
defparam desc267.B_INPUT="DIRECT";
defparam desc267.CARRYINREG=0;
defparam desc267.CARRYINSELREG=0;
defparam desc267.CREG=1;
defparam desc267.DREG=0;
defparam desc267.INMODEREG=0;
defparam desc267.MREG=1;
defparam desc267.OPMODEREG=0;
defparam desc267.PREG=0;
defparam desc267.USE_DPORT="FALSE";
defparam desc267.USE_MULT="MULTIPLY";
defparam desc267.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_4_inj (mult1_out_23,mult1_out_0,P_uc_24_0,out_inner_prod_r,vec_out_r_AQ_2,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult1_out_23 ;
output [23:0] mult1_out_0 ;
output [47:24] P_uc_24_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_2 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult1_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_24 ;
wire [17:0] BCOUT_24 ;
wire [3:0] CARRYOUT_24 ;
wire [22:0] mult1_out ;
wire [47:24] P_uc_24 ;
wire CARRYCASCOUT_24 ;
wire MULTSIGNOUT_24 ;
wire OVERFLOW_24 ;
wire PATTERNBDETECT_24 ;
wire PATTERNDETECT_24 ;
wire UNDERFLOW_24 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc475(.ACOUT(ACOUT_24[29:0]),.BCOUT(BCOUT_24[17:0]),.CARRYCASCOUT(CARRYCASCOUT_24),.CARRYOUT(CARRYOUT_24[3:0]),.MULTSIGNOUT(MULTSIGNOUT_24),.OVERFLOW(OVERFLOW_24),.P({P_uc_24[47:24],mult1_out_23,mult1_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_24),.PATTERNDETECT(PATTERNDETECT_24),.PCOUT({P_uc_24_0[47:24],mult1_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_24),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc475.ACASCREG=1;
defparam desc475.ADREG=1;
defparam desc475.ALUMODEREG=0;
defparam desc475.AREG=1;
defparam desc475.AUTORESET_PATDET="NO_RESET";
defparam desc475.A_INPUT="DIRECT";
defparam desc475.BCASCREG=2;
defparam desc475.BREG=2;
defparam desc475.B_INPUT="DIRECT";
defparam desc475.CARRYINREG=0;
defparam desc475.CARRYINSELREG=0;
defparam desc475.CREG=1;
defparam desc475.DREG=1;
defparam desc475.INMODEREG=1;
defparam desc475.MREG=0;
defparam desc475.OPMODEREG=0;
defparam desc475.PREG=0;
defparam desc475.USE_DPORT="TRUE";
defparam desc475.USE_MULT="MULTIPLY";
defparam desc475.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_5_inj (mult2_out_23,vec_out_i_AQ_2,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult2_out_23 ;
input [11:0] vec_out_i_AQ_2 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult2_out_23 ;
wire clk ;
wire [29:0] ACOUT_25 ;
wire [17:0] BCOUT_25 ;
wire [3:0] CARRYOUT_25 ;
wire [22:0] mult2_out ;
wire [47:24] P_uc_25 ;
wire [47:0] PCOUT_25 ;
wire CARRYCASCOUT_25 ;
wire MULTSIGNOUT_25 ;
wire OVERFLOW_25 ;
wire PATTERNBDETECT_25 ;
wire PATTERNDETECT_25 ;
wire UNDERFLOW_25 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc476(.ACOUT(ACOUT_25[29:0]),.BCOUT(BCOUT_25[17:0]),.CARRYCASCOUT(CARRYCASCOUT_25),.CARRYOUT(CARRYOUT_25[3:0]),.MULTSIGNOUT(MULTSIGNOUT_25),.OVERFLOW(OVERFLOW_25),.P({P_uc_25[47:24],mult2_out_23,mult2_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_25),.PATTERNDETECT(PATTERNDETECT_25),.PCOUT(PCOUT_25[47:0]),.UNDERFLOW(UNDERFLOW_25),.A({vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc476.ACASCREG=1;
defparam desc476.ADREG=0;
defparam desc476.ALUMODEREG=0;
defparam desc476.AREG=1;
defparam desc476.AUTORESET_PATDET="NO_RESET";
defparam desc476.A_INPUT="DIRECT";
defparam desc476.BCASCREG=1;
defparam desc476.BREG=1;
defparam desc476.B_INPUT="DIRECT";
defparam desc476.CARRYINREG=0;
defparam desc476.CARRYINSELREG=0;
defparam desc476.CREG=1;
defparam desc476.DREG=0;
defparam desc476.INMODEREG=0;
defparam desc476.MREG=0;
defparam desc476.OPMODEREG=0;
defparam desc476.PREG=1;
defparam desc476.USE_DPORT="FALSE";
defparam desc476.USE_MULT="MULTIPLY";
defparam desc476.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_6_inj (mult3_out_23,vec_out_r_AQ_2,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult3_out_23 ;
input [11:0] vec_out_r_AQ_2 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult3_out_23 ;
wire clk ;
wire [29:0] ACOUT_26 ;
wire [17:0] BCOUT_26 ;
wire [3:0] CARRYOUT_26 ;
wire [22:0] mult3_out ;
wire [47:24] P_uc_26 ;
wire [47:0] PCOUT_26 ;
wire CARRYCASCOUT_26 ;
wire MULTSIGNOUT_26 ;
wire OVERFLOW_26 ;
wire PATTERNBDETECT_26 ;
wire PATTERNDETECT_26 ;
wire UNDERFLOW_26 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc477(.ACOUT(ACOUT_26[29:0]),.BCOUT(BCOUT_26[17:0]),.CARRYCASCOUT(CARRYCASCOUT_26),.CARRYOUT(CARRYOUT_26[3:0]),.MULTSIGNOUT(MULTSIGNOUT_26),.OVERFLOW(OVERFLOW_26),.P({P_uc_26[47:24],mult3_out_23,mult3_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_26),.PATTERNDETECT(PATTERNDETECT_26),.PCOUT(PCOUT_26[47:0]),.UNDERFLOW(UNDERFLOW_26),.A({vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:11],vec_out_r_AQ_2[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc477.ACASCREG=1;
defparam desc477.ADREG=0;
defparam desc477.ALUMODEREG=0;
defparam desc477.AREG=1;
defparam desc477.AUTORESET_PATDET="NO_RESET";
defparam desc477.A_INPUT="DIRECT";
defparam desc477.BCASCREG=1;
defparam desc477.BREG=1;
defparam desc477.B_INPUT="DIRECT";
defparam desc477.CARRYINREG=0;
defparam desc477.CARRYINSELREG=0;
defparam desc477.CREG=1;
defparam desc477.DREG=0;
defparam desc477.INMODEREG=0;
defparam desc477.MREG=0;
defparam desc477.OPMODEREG=0;
defparam desc477.PREG=1;
defparam desc477.USE_DPORT="FALSE";
defparam desc477.USE_MULT="MULTIPLY";
defparam desc477.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_7_inj (mult4_out_23,mult4_out_0,P_uc_27_0,out_inner_prod_r,vec_out_i_AQ_2,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult4_out_23 ;
output [23:0] mult4_out_0 ;
output [47:24] P_uc_27_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_i_AQ_2 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult4_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_27 ;
wire [17:0] BCOUT_27 ;
wire [3:0] CARRYOUT_27 ;
wire [22:0] mult4_out ;
wire [47:24] P_uc_27 ;
wire CARRYCASCOUT_27 ;
wire MULTSIGNOUT_27 ;
wire OVERFLOW_27 ;
wire PATTERNBDETECT_27 ;
wire PATTERNDETECT_27 ;
wire UNDERFLOW_27 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc478(.ACOUT(ACOUT_27[29:0]),.BCOUT(BCOUT_27[17:0]),.CARRYCASCOUT(CARRYCASCOUT_27),.CARRYOUT(CARRYOUT_27[3:0]),.MULTSIGNOUT(MULTSIGNOUT_27),.OVERFLOW(OVERFLOW_27),.P({P_uc_27[47:24],mult4_out_23,mult4_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_27),.PATTERNDETECT(PATTERNDETECT_27),.PCOUT({P_uc_27_0[47:24],mult4_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_27),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:11],vec_out_i_AQ_2[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc478.ACASCREG=1;
defparam desc478.ADREG=1;
defparam desc478.ALUMODEREG=0;
defparam desc478.AREG=1;
defparam desc478.AUTORESET_PATDET="NO_RESET";
defparam desc478.A_INPUT="DIRECT";
defparam desc478.BCASCREG=2;
defparam desc478.BREG=2;
defparam desc478.B_INPUT="DIRECT";
defparam desc478.CARRYINREG=0;
defparam desc478.CARRYINSELREG=0;
defparam desc478.CREG=1;
defparam desc478.DREG=1;
defparam desc478.INMODEREG=1;
defparam desc478.MREG=0;
defparam desc478.OPMODEREG=0;
defparam desc478.PREG=0;
defparam desc478.USE_DPORT="TRUE";
defparam desc478.USE_MULT="MULTIPLY";
defparam desc478.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_8_inj (mult1_out_23,mult1_out_0,P_uc_20_0,out_inner_prod_r,vec_out_r_AQ_1,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,in_b_vec_mult_sel,clk,N_425_i,N_428_i,N_431_i,N_434_i);
output mult1_out_23 ;
output [23:0] mult1_out_0 ;
output [47:24] P_uc_20_0 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_1 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input in_b_vec_mult_sel ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire mult1_out_23 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [29:0] ACOUT_20 ;
wire [17:0] BCOUT_20 ;
wire [3:0] CARRYOUT_20 ;
wire [22:0] mult1_out ;
wire [47:24] P_uc_20 ;
wire CARRYCASCOUT_20 ;
wire MULTSIGNOUT_20 ;
wire OVERFLOW_20 ;
wire PATTERNBDETECT_20 ;
wire PATTERNDETECT_20 ;
wire UNDERFLOW_20 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc530(.ACOUT(ACOUT_20[29:0]),.BCOUT(BCOUT_20[17:0]),.CARRYCASCOUT(CARRYCASCOUT_20),.CARRYOUT(CARRYOUT_20[3:0]),.MULTSIGNOUT(MULTSIGNOUT_20),.OVERFLOW(OVERFLOW_20),.P({P_uc_20[47:24],mult1_out_23,mult1_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_20),.PATTERNDETECT(PATTERNDETECT_20),.PCOUT({P_uc_20_0[47:24],mult1_out_0[23:0]}),.UNDERFLOW(UNDERFLOW_20),.A({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:11],vec_out_r_AQ_1[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(VCC),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk),.D({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.INMODE({GND,GND,in_b_vec_mult_sel,in_b_vec_mult_sel,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc530.ACASCREG=1;
defparam desc530.ADREG=1;
defparam desc530.ALUMODEREG=0;
defparam desc530.AREG=1;
defparam desc530.AUTORESET_PATDET="NO_RESET";
defparam desc530.A_INPUT="DIRECT";
defparam desc530.BCASCREG=2;
defparam desc530.BREG=2;
defparam desc530.B_INPUT="DIRECT";
defparam desc530.CARRYINREG=0;
defparam desc530.CARRYINSELREG=0;
defparam desc530.CREG=1;
defparam desc530.DREG=1;
defparam desc530.INMODEREG=1;
defparam desc530.MREG=0;
defparam desc530.OPMODEREG=0;
defparam desc530.PREG=0;
defparam desc530.USE_DPORT="TRUE";
defparam desc530.USE_MULT="MULTIPLY";
defparam desc530.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_pipe_9_inj (mult2_out_23,vec_out_i_AQ_1,out_inner_prod_i,in_b_vec_mult_sel,clk);
output mult2_out_23 ;
input [11:0] vec_out_i_AQ_1 ;
input [11:0] out_inner_prod_i ;
input in_b_vec_mult_sel ;
input clk ;
wire mult2_out_23 ;
wire clk ;
wire [29:0] ACOUT_21 ;
wire [17:0] BCOUT_21 ;
wire [3:0] CARRYOUT_21 ;
wire [22:0] mult2_out ;
wire [47:24] P_uc_21 ;
wire [47:0] PCOUT_21 ;
wire CARRYCASCOUT_21 ;
wire MULTSIGNOUT_21 ;
wire OVERFLOW_21 ;
wire PATTERNBDETECT_21 ;
wire PATTERNDETECT_21 ;
wire UNDERFLOW_21 ;
wire VCC ;
wire GND ;
// instances
  DSP48E1 desc531(.ACOUT(ACOUT_21[29:0]),.BCOUT(BCOUT_21[17:0]),.CARRYCASCOUT(CARRYCASCOUT_21),.CARRYOUT(CARRYOUT_21[3:0]),.MULTSIGNOUT(MULTSIGNOUT_21),.OVERFLOW(OVERFLOW_21),.P({P_uc_21[47:24],mult2_out_23,mult2_out[22:0]}),.PATTERNBDETECT(PATTERNBDETECT_21),.PATTERNDETECT(PATTERNDETECT_21),.PCOUT(PCOUT_21[47:0]),.UNDERFLOW(UNDERFLOW_21),.A({vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:11],vec_out_i_AQ_1[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:11],out_inner_prod_i[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(in_b_vec_mult_sel),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc531.ACASCREG=1;
defparam desc531.ADREG=0;
defparam desc531.ALUMODEREG=0;
defparam desc531.AREG=1;
defparam desc531.AUTORESET_PATDET="NO_RESET";
defparam desc531.A_INPUT="DIRECT";
defparam desc531.BCASCREG=1;
defparam desc531.BREG=1;
defparam desc531.B_INPUT="DIRECT";
defparam desc531.CARRYINREG=0;
defparam desc531.CARRYINSELREG=0;
defparam desc531.CREG=1;
defparam desc531.DREG=0;
defparam desc531.INMODEREG=0;
defparam desc531.MREG=0;
defparam desc531.OPMODEREG=0;
defparam desc531.PREG=1;
defparam desc531.USE_DPORT="FALSE";
defparam desc531.USE_MULT="MULTIPLY";
defparam desc531.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module mult_with_reg_inj (un8_rnd_out,un8_rnd_out_P_19,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,out_inner_prod_r,pre_out_19,pre_out_20,pre_out_21,pre_out_22,pre_out_reg,N_425_i,N_428_i,N_431_i,N_434_i,N_512_i,clk,PATTERNDETECT_32);
output [10:0] un8_rnd_out ;
output un8_rnd_out_P_19 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input [11:0] out_inner_prod_r ;
output pre_out_19 ;
output pre_out_20 ;
output pre_out_21 ;
output pre_out_22 ;
output [23:23] pre_out_reg ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
input N_512_i ;
input clk ;
output PATTERNDETECT_32 ;
wire un8_rnd_out_P_19 ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire pre_out_19 ;
wire pre_out_20 ;
wire pre_out_21 ;
wire pre_out_22 ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire N_512_i ;
wire clk ;
wire PATTERNDETECT_32 ;
wire [29:0] ACOUT_12 ;
wire [17:0] BCOUT_12 ;
wire [3:0] CARRYOUT_12 ;
wire [6:0] un8_rnd_out_P ;
wire [23:20] P_uc_2 ;
wire [47:24] P_uc_12 ;
wire [47:0] PCOUT_12 ;
wire [29:0] ACOUT_32 ;
wire [17:0] BCOUT_32 ;
wire [3:0] CARRYOUT_32 ;
wire [18:0] pre_out ;
wire [47:24] P_uc_32 ;
wire [47:0] PCOUT_32 ;
wire CARRYCASCOUT_12 ;
wire MULTSIGNOUT_12 ;
wire OVERFLOW_12 ;
wire N_3 ;
wire PATTERNBDETECT_12 ;
wire PATTERNDETECT_12 ;
wire UNDERFLOW_12 ;
wire VCC ;
wire GND ;
wire CARRYCASCOUT_32 ;
wire MULTSIGNOUT_32 ;
wire OVERFLOW_32 ;
wire PATTERNBDETECT_32 ;
wire UNDERFLOW_32 ;
// instances
  DSP48E1 desc843(.ACOUT(ACOUT_12[29:0]),.BCOUT(BCOUT_12[17:0]),.CARRYCASCOUT(CARRYCASCOUT_12),.CARRYOUT(CARRYOUT_12[3:0]),.MULTSIGNOUT(MULTSIGNOUT_12),.OVERFLOW(OVERFLOW_12),.P({P_uc_12[47:24],P_uc_2[23:20],un8_rnd_out_P_19,un8_rnd_out[10:0],N_3,un8_rnd_out_P[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_12),.PATTERNDETECT(PATTERNDETECT_12),.PCOUT(PCOUT_12[47:0]),.UNDERFLOW(UNDERFLOW_12),.A({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,GND,GND,GND,GND,GND,GND,GND}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(N_512_i),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,VCC,VCC,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc843.ACASCREG=2;
defparam desc843.ADREG=0;
defparam desc843.ALUMODEREG=0;
defparam desc843.AREG=2;
defparam desc843.AUTORESET_PATDET="NO_RESET";
defparam desc843.A_INPUT="DIRECT";
defparam desc843.BCASCREG=1;
defparam desc843.BREG=1;
defparam desc843.B_INPUT="DIRECT";
defparam desc843.CARRYINREG=0;
defparam desc843.CARRYINSELREG=0;
defparam desc843.CREG=0;
defparam desc843.DREG=0;
defparam desc843.INMODEREG=0;
defparam desc843.MREG=0;
defparam desc843.OPMODEREG=0;
defparam desc843.PREG=0;
defparam desc843.USE_DPORT="FALSE";
defparam desc843.USE_MULT="MULTIPLY";
defparam desc843.USE_SIMD="ONE48";
  DSP48E1 desc844(.ACOUT(ACOUT_32[29:0]),.BCOUT(BCOUT_32[17:0]),.CARRYCASCOUT(CARRYCASCOUT_32),.CARRYOUT(CARRYOUT_32[3:0]),.MULTSIGNOUT(MULTSIGNOUT_32),.OVERFLOW(OVERFLOW_32),.P({P_uc_32[47:24],pre_out_reg[23:23],pre_out_22,pre_out_21,pre_out_20,pre_out_19,pre_out[18:0]}),.PATTERNBDETECT(PATTERNBDETECT_32),.PATTERNDETECT(PATTERNDETECT_32),.PCOUT(PCOUT_32[47:0]),.UNDERFLOW(UNDERFLOW_32),.A({out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_11,out_inv_sqrt_10,out_inv_sqrt_9,out_inv_sqrt_8,out_inv_sqrt_7,N_434_i,N_431_i,N_428_i,N_425_i,out_inv_sqrt_2,out_inv_sqrt_1,out_inv_sqrt_0}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(N_512_i),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc844.ACASCREG=2;
defparam desc844.ADREG=0;
defparam desc844.ALUMODEREG=0;
defparam desc844.AREG=2;
defparam desc844.AUTORESET_PATDET="NO_RESET";
defparam desc844.A_INPUT="DIRECT";
defparam desc844.BCASCREG=1;
defparam desc844.BREG=1;
defparam desc844.B_INPUT="DIRECT";
defparam desc844.CARRYINREG=0;
defparam desc844.CARRYINSELREG=0;
defparam desc844.CREG=1;
defparam desc844.DREG=0;
defparam desc844.INMODEREG=0;
defparam desc844.MASK=48'b111111111111111111111111011111111111111111111111;
defparam desc844.MREG=0;
defparam desc844.OPMODEREG=0;
defparam desc844.PATTERN=48'b111111111111111111111111111111111111111111111111;
defparam desc844.PREG=0;
defparam desc844.SEL_MASK="MASK";
defparam desc844.USE_DPORT="FALSE";
defparam desc844.USE_MULT="MULTIPLY";
defparam desc844.USE_PATTERN_DETECT="PATDET";
defparam desc844.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module multiplier_inj (mult1_out,pre_output);
output [11:0] mult1_out ;
input [11:0] pre_output ;
wire [23:0] pre_out ;
wire [18:8] un8_rnd_out_P ;
wire [19:19] un8_rnd_out_P_0 ;
wire [29:0] ACOUT_9 ;
wire [17:0] BCOUT_9 ;
wire [3:0] CARRYOUT_9 ;
wire [6:0] un8_rnd_out_P_1 ;
wire [23:20] P_uc ;
wire [47:24] P_uc_9 ;
wire [47:0] PCOUT_9 ;
wire [29:0] ACOUT_13 ;
wire [17:0] BCOUT_13 ;
wire [3:0] CARRYOUT_13 ;
wire [47:24] P_uc_13 ;
wire [47:0] PCOUT_13 ;
wire un5_output_3_0 ;
wire PATTERNDETECT_13 ;
wire CARRYCASCOUT_9 ;
wire MULTSIGNOUT_9 ;
wire OVERFLOW_9 ;
wire N_15 ;
wire PATTERNBDETECT_9 ;
wire PATTERNDETECT_9 ;
wire UNDERFLOW_9 ;
wire VCC ;
wire GND ;
wire CARRYCASCOUT_13 ;
wire MULTSIGNOUT_13 ;
wire OVERFLOW_13 ;
wire PATTERNBDETECT_13 ;
wire UNDERFLOW_13 ;
// instances
  LUT2 desc910(.I0(pre_out[21:21]),.I1(pre_out[22:22]),.O(un5_output_3_0));
defparam desc910.INIT=4'h8;
  LUT6 desc911(.I0(un8_rnd_out_P[8:8]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[0:0]));
defparam desc911.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc912(.I0(un8_rnd_out_P[9:9]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[1:1]));
defparam desc912.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc913(.I0(un8_rnd_out_P[10:10]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[2:2]));
defparam desc913.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc914(.I0(un8_rnd_out_P[11:11]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[3:3]));
defparam desc914.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc915(.I0(un8_rnd_out_P[12:12]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[4:4]));
defparam desc915.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc916(.I0(un8_rnd_out_P[13:13]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[5:5]));
defparam desc916.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc917(.I0(un8_rnd_out_P[14:14]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[6:6]));
defparam desc917.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc918(.I0(un8_rnd_out_P[15:15]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[7:7]));
defparam desc918.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc919(.I0(un8_rnd_out_P[16:16]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[8:8]));
defparam desc919.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc920(.I0(un8_rnd_out_P[17:17]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[9:9]));
defparam desc920.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc921(.I0(un8_rnd_out_P[18:18]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[10:10]));
defparam desc921.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc922(.I0(un8_rnd_out_P_0[19:19]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_13),.O(mult1_out[11:11]));
defparam desc922.INIT=64'hBFAAFFAABF00FF00;
  DSP48E1 desc923(.ACOUT(ACOUT_9[29:0]),.BCOUT(BCOUT_9[17:0]),.CARRYCASCOUT(CARRYCASCOUT_9),.CARRYOUT(CARRYOUT_9[3:0]),.MULTSIGNOUT(MULTSIGNOUT_9),.OVERFLOW(OVERFLOW_9),.P({P_uc_9[47:24],P_uc[23:20],un8_rnd_out_P_0[19:19],un8_rnd_out_P[18:8],N_15,un8_rnd_out_P_1[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_9),.PATTERNDETECT(PATTERNDETECT_9),.PCOUT(PCOUT_9[47:0]),.UNDERFLOW(UNDERFLOW_9),.A({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,GND,GND,GND,GND,GND,GND,GND}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(GND),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,VCC,VCC,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc923.ACASCREG=0;
defparam desc923.ADREG=0;
defparam desc923.ALUMODEREG=0;
defparam desc923.AREG=0;
defparam desc923.AUTORESET_PATDET="NO_RESET";
defparam desc923.A_INPUT="DIRECT";
defparam desc923.BCASCREG=0;
defparam desc923.BREG=0;
defparam desc923.B_INPUT="DIRECT";
defparam desc923.CARRYINREG=0;
defparam desc923.CARRYINSELREG=0;
defparam desc923.CREG=0;
defparam desc923.DREG=0;
defparam desc923.INMODEREG=0;
defparam desc923.MREG=0;
defparam desc923.OPMODEREG=0;
defparam desc923.PREG=0;
defparam desc923.USE_DPORT="FALSE";
defparam desc923.USE_MULT="MULTIPLY";
defparam desc923.USE_SIMD="ONE48";
  DSP48E1 desc924(.ACOUT(ACOUT_13[29:0]),.BCOUT(BCOUT_13[17:0]),.CARRYCASCOUT(CARRYCASCOUT_13),.CARRYOUT(CARRYOUT_13[3:0]),.MULTSIGNOUT(MULTSIGNOUT_13),.OVERFLOW(OVERFLOW_13),.P({P_uc_13[47:24],pre_out[23:0]}),.PATTERNBDETECT(PATTERNBDETECT_13),.PATTERNDETECT(PATTERNDETECT_13),.PCOUT(PCOUT_13[47:0]),.UNDERFLOW(UNDERFLOW_13),.A({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(GND),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc924.ACASCREG=0;
defparam desc924.ADREG=0;
defparam desc924.ALUMODEREG=0;
defparam desc924.AREG=0;
defparam desc924.AUTORESET_PATDET="NO_RESET";
defparam desc924.A_INPUT="DIRECT";
defparam desc924.BCASCREG=0;
defparam desc924.BREG=0;
defparam desc924.B_INPUT="DIRECT";
defparam desc924.CARRYINREG=0;
defparam desc924.CARRYINSELREG=0;
defparam desc924.CREG=1;
defparam desc924.DREG=0;
defparam desc924.INMODEREG=0;
defparam desc924.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc924.MREG=0;
defparam desc924.OPMODEREG=0;
defparam desc924.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc924.PREG=0;
defparam desc924.SEL_MASK="MASK";
defparam desc924.USE_DPORT="FALSE";
defparam desc924.USE_MULT="MULTIPLY";
defparam desc924.USE_PATTERN_DETECT="PATDET";
defparam desc924.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module multiplier_1_inj (mult2_out,pre_output,out_inner_prod_r,start_inv_sqrt,clk);
output [11:0] mult2_out ;
input [11:0] pre_output ;
input [11:0] out_inner_prod_r ;
input start_inv_sqrt ;
input clk ;
wire start_inv_sqrt ;
wire clk ;
wire [23:0] pre_out ;
wire [18:0] un8_rnd_out_P_0 ;
wire [19:19] un8_rnd_out_P_1 ;
wire [29:0] ACOUT_10 ;
wire [17:0] BCOUT_10 ;
wire [3:0] CARRYOUT_10 ;
wire [23:20] P_uc_0 ;
wire [47:24] P_uc_10 ;
wire [47:0] PCOUT_10 ;
wire [29:0] ACOUT_14 ;
wire [17:0] BCOUT_14 ;
wire [3:0] CARRYOUT_14 ;
wire [47:24] P_uc_14 ;
wire [47:0] PCOUT_14 ;
wire un5_output_3_0 ;
wire PATTERNDETECT_14 ;
wire CARRYCASCOUT_10 ;
wire MULTSIGNOUT_10 ;
wire OVERFLOW_10 ;
wire N_3 ;
wire PATTERNBDETECT_10 ;
wire PATTERNDETECT_10 ;
wire UNDERFLOW_10 ;
wire VCC ;
wire GND ;
wire CARRYCASCOUT_14 ;
wire MULTSIGNOUT_14 ;
wire OVERFLOW_14 ;
wire PATTERNBDETECT_14 ;
wire UNDERFLOW_14 ;
// instances
  LUT2 desc925(.I0(pre_out[21:21]),.I1(pre_out[22:22]),.O(un5_output_3_0));
defparam desc925.INIT=4'h8;
  LUT6 desc926(.I0(un8_rnd_out_P_0[8:8]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[0:0]));
defparam desc926.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc927(.I0(un8_rnd_out_P_0[9:9]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[1:1]));
defparam desc927.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc928(.I0(un8_rnd_out_P_0[10:10]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[2:2]));
defparam desc928.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc929(.I0(un8_rnd_out_P_0[11:11]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[3:3]));
defparam desc929.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc930(.I0(un8_rnd_out_P_0[12:12]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[4:4]));
defparam desc930.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc931(.I0(un8_rnd_out_P_0[13:13]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[5:5]));
defparam desc931.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc932(.I0(un8_rnd_out_P_0[14:14]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[6:6]));
defparam desc932.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc933(.I0(un8_rnd_out_P_0[15:15]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[7:7]));
defparam desc933.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc934(.I0(un8_rnd_out_P_0[16:16]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[8:8]));
defparam desc934.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc935(.I0(un8_rnd_out_P_0[17:17]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[9:9]));
defparam desc935.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc936(.I0(un8_rnd_out_P_0[18:18]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[10:10]));
defparam desc936.INIT=64'h80AA00AA80FF00FF;
  LUT6 desc937(.I0(un8_rnd_out_P_1[19:19]),.I1(pre_out[19:19]),.I2(pre_out[20:20]),.I3(pre_out[23:23]),.I4(un5_output_3_0),.I5(PATTERNDETECT_14),.O(mult2_out[11:11]));
defparam desc937.INIT=64'hBFAAFFAABF00FF00;
  DSP48E1 desc938(.ACOUT(ACOUT_10[29:0]),.BCOUT(BCOUT_10[17:0]),.CARRYCASCOUT(CARRYCASCOUT_10),.CARRYOUT(CARRYOUT_10[3:0]),.MULTSIGNOUT(MULTSIGNOUT_10),.OVERFLOW(OVERFLOW_10),.P({P_uc_10[47:24],P_uc_0[23:20],un8_rnd_out_P_1[19:19],un8_rnd_out_P_0[18:8],N_3,un8_rnd_out_P_0[6:0]}),.PATTERNBDETECT(PATTERNBDETECT_10),.PATTERNDETECT(PATTERNDETECT_10),.PCOUT(PCOUT_10[47:0]),.UNDERFLOW(UNDERFLOW_10),.A({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,GND,GND,GND,GND,GND,GND,GND}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(start_inv_sqrt),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,VCC,VCC,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc938.ACASCREG=0;
defparam desc938.ADREG=0;
defparam desc938.ALUMODEREG=0;
defparam desc938.AREG=0;
defparam desc938.AUTORESET_PATDET="NO_RESET";
defparam desc938.A_INPUT="DIRECT";
defparam desc938.BCASCREG=1;
defparam desc938.BREG=1;
defparam desc938.B_INPUT="DIRECT";
defparam desc938.CARRYINREG=0;
defparam desc938.CARRYINSELREG=0;
defparam desc938.CREG=0;
defparam desc938.DREG=0;
defparam desc938.INMODEREG=0;
defparam desc938.MREG=0;
defparam desc938.OPMODEREG=0;
defparam desc938.PREG=0;
defparam desc938.USE_DPORT="FALSE";
defparam desc938.USE_MULT="MULTIPLY";
defparam desc938.USE_SIMD="ONE48";
  DSP48E1 desc939(.ACOUT(ACOUT_14[29:0]),.BCOUT(BCOUT_14[17:0]),.CARRYCASCOUT(CARRYCASCOUT_14),.CARRYOUT(CARRYOUT_14[3:0]),.MULTSIGNOUT(MULTSIGNOUT_14),.OVERFLOW(OVERFLOW_14),.P({P_uc_14[47:24],pre_out[23:0]}),.PATTERNBDETECT(PATTERNBDETECT_14),.PATTERNDETECT(PATTERNDETECT_14),.PCOUT(PCOUT_14[47:0]),.UNDERFLOW(UNDERFLOW_14),.A({pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:11],pre_output[11:0]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:11],out_inner_prod_r[11:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(start_inv_sqrt),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(GND),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc939.ACASCREG=0;
defparam desc939.ADREG=0;
defparam desc939.ALUMODEREG=0;
defparam desc939.AREG=0;
defparam desc939.AUTORESET_PATDET="NO_RESET";
defparam desc939.A_INPUT="DIRECT";
defparam desc939.BCASCREG=1;
defparam desc939.BREG=1;
defparam desc939.B_INPUT="DIRECT";
defparam desc939.CARRYINREG=0;
defparam desc939.CARRYINSELREG=0;
defparam desc939.CREG=1;
defparam desc939.DREG=0;
defparam desc939.INMODEREG=0;
defparam desc939.MASK=48'b111111111111111111111111100001111111111111111111;
defparam desc939.MREG=0;
defparam desc939.OPMODEREG=0;
defparam desc939.PATTERN=48'b111111111111111111111111100001111111111111111111;
defparam desc939.PREG=0;
defparam desc939.SEL_MASK="MASK";
defparam desc939.USE_DPORT="FALSE";
defparam desc939.USE_MULT="MULTIPLY";
defparam desc939.USE_PATTERN_DETECT="PATDET";
defparam desc939.USE_SIMD="ONE48";
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module qr_decomp_inj (out_Q_r,out_Q_i,col_sel_R,out_R_i,out_R_r,col_sel_AQ,in_A_r,in_A_i,clk,rst,wr_A_QR,start_QR,done_QR,red_mat_reg_0,p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_,p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_,p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_,p_desc951_p_O_FDEinv_sqrt_,p_desc952_p_O_FDEinv_sqrt_,p_desc953_p_O_FDEinv_sqrt_,p_desc954_p_O_FDEinv_sqrt_,p_desc955_p_O_FDEinv_sqrt_,p_desc956_p_O_FDEinv_sqrt_,p_desc957_p_O_FDEinv_sqrt_,p_desc958_p_O_FDEinv_sqrt_,p_desc959_p_O_FDEinv_sqrt_,p_desc960_p_O_FDEinv_sqrt_,p_desc961_p_O_FDEinv_sqrt_,p_desc962_p_O_FDEinv_sqrt_,p_desc48_p_O_FDEr_mat_regs_,p_desc49_p_O_FDEr_mat_regs_,p_desc50_p_O_FDEr_mat_regs_,p_desc51_p_O_FDEr_mat_regs_,p_desc52_p_O_FDEr_mat_regs_,p_desc53_p_O_FDEr_mat_regs_,p_desc54_p_O_FDEr_mat_regs_,p_desc55_p_O_FDEr_mat_regs_,p_desc56_p_O_FDEr_mat_regs_,p_desc57_p_O_FDEr_mat_regs_,p_desc58_p_O_FDEr_mat_regs_,p_desc59_p_O_FDEr_mat_regs_,p_desc60_p_O_FDEr_mat_regs_,p_desc61_p_O_FDEr_mat_regs_,p_desc62_p_O_FDEr_mat_regs_,p_desc63_p_O_FDEr_mat_regs_,p_desc64_p_O_FDEr_mat_regs_,p_desc65_p_O_FDEr_mat_regs_,p_desc66_p_O_FDEr_mat_regs_,p_desc67_p_O_FDEr_mat_regs_,p_desc68_p_O_FDEr_mat_regs_,p_desc69_p_O_FDEr_mat_regs_,p_desc70_p_O_FDEr_mat_regs_,p_desc71_p_O_FDEr_mat_regs_,p_desc72_p_O_FDEr_mat_regs_,p_desc73_p_O_FDEr_mat_regs_,p_desc74_p_O_FDEr_mat_regs_,p_desc75_p_O_FDEr_mat_regs_,p_desc76_p_O_FDEr_mat_regs_,p_desc77_p_O_FDEr_mat_regs_,p_desc78_p_O_FDEr_mat_regs_,p_desc79_p_O_FDEr_mat_regs_,p_desc80_p_O_FDEr_mat_regs_,p_desc81_p_O_FDEr_mat_regs_,p_desc82_p_O_FDEr_mat_regs_,p_desc83_p_O_FDEr_mat_regs_,p_desc84_p_O_FDEr_mat_regs_,p_desc85_p_O_FDEr_mat_regs_,p_desc86_p_O_FDEr_mat_regs_,p_desc87_p_O_FDEr_mat_regs_,p_desc88_p_O_FDEr_mat_regs_,p_desc89_p_O_FDEr_mat_regs_,p_desc90_p_O_FDEr_mat_regs_,p_desc91_p_O_FDEr_mat_regs_,p_desc92_p_O_FDEr_mat_regs_,p_desc93_p_O_FDEr_mat_regs_,p_desc94_p_O_FDEr_mat_regs_,p_desc95_p_O_FDEr_mat_regs_,p_desc96_p_O_FDEr_mat_regs_,p_desc97_p_O_FDEr_mat_regs_,p_desc98_p_O_FDEr_mat_regs_,p_desc99_p_O_FDEr_mat_regs_,p_desc100_p_O_FDEr_mat_regs_,p_desc101_p_O_FDEr_mat_regs_,p_desc102_p_O_FDEr_mat_regs_,p_desc103_p_O_FDEr_mat_regs_,p_desc104_p_O_FDEr_mat_regs_,p_desc105_p_O_FDEr_mat_regs_,p_desc106_p_O_FDEr_mat_regs_,p_desc107_p_O_FDEr_mat_regs_,p_desc108_p_O_FDEr_mat_regs_,p_desc109_p_O_FDEr_mat_regs_,p_desc110_p_O_FDEr_mat_regs_,p_desc111_p_O_FDEr_mat_regs_,p_desc112_p_O_FDEr_mat_regs_,p_desc113_p_O_FDEr_mat_regs_,p_desc114_p_O_FDEr_mat_regs_,p_desc115_p_O_FDEr_mat_regs_,p_desc116_p_O_FDEr_mat_regs_,p_desc117_p_O_FDEr_mat_regs_,p_desc118_p_O_FDEr_mat_regs_,p_desc119_p_O_FDEr_mat_regs_,p_desc120_p_O_FDEr_mat_regs_,p_desc121_p_O_FDEr_mat_regs_,p_desc122_p_O_FDEr_mat_regs_,p_desc123_p_O_FDEr_mat_regs_,p_desc124_p_O_FDEr_mat_regs_,p_desc125_p_O_FDEr_mat_regs_,p_desc126_p_O_FDEr_mat_regs_,p_desc127_p_O_FDEr_mat_regs_,p_desc128_p_O_FDEr_mat_regs_,p_desc129_p_O_FDEr_mat_regs_,p_desc130_p_O_FDEr_mat_regs_,p_desc131_p_O_FDEr_mat_regs_,p_desc132_p_O_FDEr_mat_regs_,p_desc133_p_O_FDEr_mat_regs_,p_desc134_p_O_FDEr_mat_regs_,p_desc135_p_O_FDEr_mat_regs_,p_desc136_p_O_FDEr_mat_regs_,p_desc137_p_O_FDEr_mat_regs_,p_desc138_p_O_FDEr_mat_regs_,p_desc139_p_O_FDEr_mat_regs_,p_desc140_p_O_FDEr_mat_regs_,p_desc141_p_O_FDEr_mat_regs_,p_desc142_p_O_FDEr_mat_regs_,p_desc143_p_O_FDEr_mat_regs_,p_desc144_p_O_FDEr_mat_regs_,p_desc145_p_O_FDEr_mat_regs_,p_desc146_p_O_FDEr_mat_regs_,p_desc147_p_O_FDEr_mat_regs_,p_desc148_p_O_FDEr_mat_regs_,p_desc149_p_O_FDEr_mat_regs_,p_desc150_p_O_FDEr_mat_regs_,p_desc151_p_O_FDEr_mat_regs_,p_desc152_p_O_FDEr_mat_regs_,p_desc153_p_O_FDEr_mat_regs_,p_desc154_p_O_FDEr_mat_regs_,p_desc155_p_O_FDEr_mat_regs_,p_desc156_p_O_FDEr_mat_regs_,p_desc157_p_O_FDEr_mat_regs_,p_desc158_p_O_FDEr_mat_regs_,p_desc159_p_O_FDEr_mat_regs_,p_desc160_p_O_FDEr_mat_regs_,p_desc161_p_O_FDEr_mat_regs_,p_desc162_p_O_FDEr_mat_regs_,p_desc163_p_O_FDEr_mat_regs_,p_desc164_p_O_FDEr_mat_regs_,p_desc165_p_O_FDEr_mat_regs_,p_desc166_p_O_FDEr_mat_regs_,p_desc167_p_O_FDEr_mat_regs_,p_desc168_p_O_FDEr_mat_regs_,p_desc169_p_O_FDEr_mat_regs_,p_desc170_p_O_FDEr_mat_regs_,p_desc171_p_O_FDEr_mat_regs_,p_desc172_p_O_FDEr_mat_regs_,p_desc173_p_O_FDEr_mat_regs_,p_desc174_p_O_FDEr_mat_regs_,p_desc175_p_O_FDEr_mat_regs_,p_desc176_p_O_FDEr_mat_regs_,p_desc177_p_O_FDEr_mat_regs_,p_desc178_p_O_FDEr_mat_regs_,p_desc179_p_O_FDEr_mat_regs_,p_desc180_p_O_FDEr_mat_regs_,p_desc181_p_O_FDEr_mat_regs_,p_desc182_p_O_FDEr_mat_regs_,p_desc183_p_O_FDEr_mat_regs_,p_desc184_p_O_FDEr_mat_regs_,p_desc185_p_O_FDEr_mat_regs_,p_desc186_p_O_FDEr_mat_regs_,p_desc187_p_O_FDEr_mat_regs_,p_desc188_p_O_FDEr_mat_regs_,p_desc189_p_O_FDEr_mat_regs_,p_desc190_p_O_FDEr_mat_regs_,p_desc191_p_O_FDEr_mat_regs_,p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_,p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_,p_desc739_p_O_FDEvec_sub_,p_desc740_p_O_FDEvec_sub_,p_desc741_p_O_FDEvec_sub_,p_desc742_p_O_FDEvec_sub_,p_desc743_p_O_FDEvec_sub_,p_desc744_p_O_FDEvec_sub_,p_desc745_p_O_FDEvec_sub_,p_desc746_p_O_FDEvec_sub_,p_desc747_p_O_FDEvec_sub_,p_desc748_p_O_FDEvec_sub_,p_desc749_p_O_FDEvec_sub_,p_desc750_p_O_FDEvec_sub_,p_desc751_p_O_FDEvec_sub_,p_desc752_p_O_FDEvec_sub_,p_desc753_p_O_FDEvec_sub_,p_desc754_p_O_FDEvec_sub_,p_desc755_p_O_FDEvec_sub_,p_desc756_p_O_FDEvec_sub_,p_desc757_p_O_FDEvec_sub_,p_desc758_p_O_FDEvec_sub_,p_desc759_p_O_FDEvec_sub_,p_desc760_p_O_FDEvec_sub_,p_desc761_p_O_FDEvec_sub_,p_desc762_p_O_FDEvec_sub_,p_desc763_p_O_FDEvec_sub_,p_desc764_p_O_FDEvec_sub_,p_desc765_p_O_FDEvec_sub_,p_desc766_p_O_FDEvec_sub_,p_desc767_p_O_FDEvec_sub_,p_desc768_p_O_FDEvec_sub_,p_desc769_p_O_FDEvec_sub_,p_desc770_p_O_FDEvec_sub_,p_desc771_p_O_FDEvec_sub_,p_desc772_p_O_FDEvec_sub_,p_desc773_p_O_FDEvec_sub_,p_desc774_p_O_FDEvec_sub_,p_desc775_p_O_FDEvec_sub_,p_desc776_p_O_FDEvec_sub_,p_desc777_p_O_FDEvec_sub_,p_desc778_p_O_FDEvec_sub_,p_desc779_p_O_FDEvec_sub_,p_desc780_p_O_FDEvec_sub_,p_desc781_p_O_FDEvec_sub_,p_desc782_p_O_FDEvec_sub_,p_desc783_p_O_FDEvec_sub_,p_desc784_p_O_FDEvec_sub_,p_desc785_p_O_FDEvec_sub_,p_desc786_p_O_FDEvec_sub_,p_desc787_p_O_FDEvec_sub_,p_desc788_p_O_FDEvec_sub_,p_desc789_p_O_FDEvec_sub_,p_desc790_p_O_FDEvec_sub_,p_desc791_p_O_FDEvec_sub_,p_desc792_p_O_FDEvec_sub_,p_desc793_p_O_FDEvec_sub_,p_desc794_p_O_FDEvec_sub_,p_desc795_p_O_FDEvec_sub_,p_desc796_p_O_FDEvec_sub_,p_desc797_p_O_FDEvec_sub_,p_desc798_p_O_FDEvec_sub_,p_desc799_p_O_FDEvec_sub_,p_desc800_p_O_FDEvec_sub_,p_desc801_p_O_FDEvec_sub_,p_desc802_p_O_FDEvec_sub_,p_desc803_p_O_FDEvec_sub_,p_desc804_p_O_FDEvec_sub_,p_desc805_p_O_FDEvec_sub_,p_desc806_p_O_FDEvec_sub_,p_desc807_p_O_FDEvec_sub_,p_desc808_p_O_FDEvec_sub_,p_desc809_p_O_FDEvec_sub_,p_desc810_p_O_FDEvec_sub_,p_desc811_p_O_FDEvec_sub_,p_desc812_p_O_FDEvec_sub_,p_desc813_p_O_FDEvec_sub_,p_desc814_p_O_FDEvec_sub_,p_desc815_p_O_FDEvec_sub_,p_desc816_p_O_FDEvec_sub_,p_desc817_p_O_FDEvec_sub_,p_desc818_p_O_FDEvec_sub_,p_desc819_p_O_FDEvec_sub_,p_desc820_p_O_FDEvec_sub_,p_desc821_p_O_FDEvec_sub_,p_desc822_p_O_FDEvec_sub_,p_desc823_p_O_FDEvec_sub_,p_desc824_p_O_FDEvec_sub_,p_desc825_p_O_FDEvec_sub_,p_desc826_p_O_FDEvec_sub_,p_desc827_p_O_FDEvec_sub_,p_desc828_p_O_FDEvec_sub_,p_desc829_p_O_FDEvec_sub_,p_desc830_p_O_FDEvec_sub_,p_desc831_p_O_FDEvec_sub_,p_desc832_p_O_FDEvec_sub_,p_desc833_p_O_FDEvec_sub_,p_desc834_p_O_FDEvec_sub_,p_output_reg_pipe_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_,p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_,p_desc318_p_O_FDCinner_prod_,p_desc319_p_O_FDCinner_prod_,p_desc320_p_O_FDCinner_prod_,p_desc321_p_O_FDCinner_prod_,p_desc322_p_O_FDCinner_prod_,p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_,p_done_Z_p_O_FDCinner_prod_,p_acc_enable_Z_p_O_FDCinner_prod_,p_desc325_p_O_FDCinner_prod_,p_desc326_p_O_FDCinner_prod_,p_desc327_p_O_FDCinner_prod_,p_desc328_p_O_FDCinner_prod_,p_desc329_p_O_FDCinner_prod_,p_desc330_p_O_FDCinner_prod_,p_desc331_p_O_FDCinner_prod_,p_desc332_p_O_FDCinner_prod_,p_desc333_p_O_FDCinner_prod_,p_desc334_p_O_FDCinner_prod_,p_desc335_p_O_FDCinner_prod_,p_desc336_p_O_FDCinner_prod_,p_desc337_p_O_FDCinner_prod_,p_desc338_p_O_FDCinner_prod_,p_desc339_p_O_FDCinner_prod_,p_desc340_p_O_FDCinner_prod_,p_desc341_p_O_FDCinner_prod_,p_desc342_p_O_FDCinner_prod_,p_desc343_p_O_FDCinner_prod_,p_desc344_p_O_FDCinner_prod_,p_desc345_p_O_FDCinner_prod_,p_desc346_p_O_FDCinner_prod_,p_desc347_p_O_FDCinner_prod_,p_desc348_p_O_FDCinner_prod_,p_desc349_p_O_FDCinner_prod_,p_desc350_p_O_FDCinner_prod_,p_desc375_p_O_FDCinner_prod_,p_desc376_p_O_FDCinner_prod_,p_desc377_p_O_FDCinner_prod_,p_desc378_p_O_FDCinner_prod_,p_desc379_p_O_FDCinner_prod_,p_desc380_p_O_FDCinner_prod_,p_desc381_p_O_FDCinner_prod_,p_desc382_p_O_FDCinner_prod_,p_desc383_p_O_FDCinner_prod_,p_desc384_p_O_FDCinner_prod_,p_desc385_p_O_FDCinner_prod_,p_desc386_p_O_FDCinner_prod_,p_desc387_p_O_FDCinner_prod_,p_desc388_p_O_FDCinner_prod_,p_desc389_p_O_FDCinner_prod_,p_desc390_p_O_FDCinner_prod_,p_desc391_p_O_FDCinner_prod_,p_desc392_p_O_FDCinner_prod_,p_desc393_p_O_FDCinner_prod_,p_desc394_p_O_FDCinner_prod_,p_desc395_p_O_FDCinner_prod_,p_desc396_p_O_FDCinner_prod_,p_desc397_p_O_FDCinner_prod_,p_desc398_p_O_FDCinner_prod_,p_done_Z_p_O_FDCinv_sqrt_,p_desc946_p_O_FDCinv_sqrt_,p_desc947_p_O_FDCinv_sqrt_,p_desc948_p_O_FDCinv_sqrt_,p_desc949_p_O_FDCinv_sqrt_,p_desc950_p_O_FDCinv_sqrt_,p_desc1255_p_O_FDCqr_decomp_ctl_,p_desc1256_p_O_FDCqr_decomp_ctl_,p_desc1257_p_O_FDCqr_decomp_ctl_,p_desc1258_p_O_FDCqr_decomp_ctl_,p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_,p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_,p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_,p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_,p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_,p_desc1274_p_O_FDCqr_decomp_ctl_,p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_,p_done_Z_p_O_FDCqr_decomp_ctl_,p_desc1275_p_O_FDCqr_decomp_ctl_,p_desc1276_p_O_FDCqr_decomp_ctl_,p_desc1277_p_O_FDCqr_decomp_ctl_,p_desc1278_p_O_FDCqr_decomp_ctl_,p_desc1279_p_O_FDCqr_decomp_ctl_,p_desc1281_p_O_FDCqr_decomp_ctl_,p_desc1282_p_O_FDCqr_decomp_ctl_,p_desc1283_p_O_FDCqr_decomp_ctl_,p_desc1284_p_O_FDCqr_decomp_ctl_,p_desc1285_p_O_FDCqr_decomp_ctl_,p_desc1286_p_O_FDCqr_decomp_ctl_,p_desc1287_p_O_FDCqr_decomp_ctl_,p_desc1288_p_O_FDCqr_decomp_ctl_,p_acc_clear_Z_p_O_FDPinner_prod_,p_desc1265_p_O_FDPqr_decomp_ctl_,p_desc1268_p_O_FDPqr_decomp_ctl_,p_desc1280_p_O_FDPqr_decomp_ctl_,p_desc324_p_O_FDCEinner_prod_,p_desc351_p_O_FDCEinner_prod_,p_desc352_p_O_FDCEinner_prod_,p_desc353_p_O_FDCEinner_prod_,p_desc354_p_O_FDCEinner_prod_,p_desc355_p_O_FDCEinner_prod_,p_desc356_p_O_FDCEinner_prod_,p_desc357_p_O_FDCEinner_prod_,p_desc358_p_O_FDCEinner_prod_,p_desc359_p_O_FDCEinner_prod_,p_desc360_p_O_FDCEinner_prod_,p_desc361_p_O_FDCEinner_prod_,p_desc362_p_O_FDCEinner_prod_,p_desc363_p_O_FDCEinner_prod_,p_desc364_p_O_FDCEinner_prod_,p_desc365_p_O_FDCEinner_prod_,p_desc366_p_O_FDCEinner_prod_,p_desc367_p_O_FDCEinner_prod_,p_desc368_p_O_FDCEinner_prod_,p_desc369_p_O_FDCEinner_prod_,p_desc370_p_O_FDCEinner_prod_,p_desc371_p_O_FDCEinner_prod_,p_desc372_p_O_FDCEinner_prod_,p_desc373_p_O_FDCEinner_prod_,p_desc374_p_O_FDCEinner_prod_,p_desc1263_p_O_FDCEqr_decomp_ctl_,p_desc1264_p_O_FDCEqr_decomp_ctl_,p_desc1266_p_O_FDCEqr_decomp_ctl_,p_desc1267_p_O_FDCEqr_decomp_ctl_,p_desc1269_p_O_FDCEqr_decomp_ctl_,p_desc1270_p_O_FDCEqr_decomp_ctl_,p_desc1271_p_O_FDCEqr_decomp_ctl_,p_desc1272_p_O_FDCEqr_decomp_ctl_,p_desc1273_p_O_FDCEqr_decomp_ctl_);
output [47:0] out_Q_r ;
output [47:0] out_Q_i ;
input [1:0] col_sel_R ;
output [47:12] out_R_i ;
output [47:0] out_R_r ;
input [1:0] col_sel_AQ ;
input [47:0] in_A_r ;
input [47:0] in_A_i ;
input clk ;
input rst ;
input wr_A_QR ;
input start_QR ;
output done_QR ;
input red_mat_reg_0 ;
wire clk ;
wire rst ;
wire wr_A_QR ;
wire start_QR ;
wire done_QR ;
wire red_mat_reg_0 ;
wire col_sel_AQ2_mux_i_m3_lut6_2_O6 ;
wire col_sel_AQ2_mux_i_m3_lut6_2_O5 ;
wire [1:0] col_sel_AQ_int ;
wire w_col_sel_AQ_mux_i_m3_lut6_2_O6 ;
wire w_col_sel_AQ_mux_i_m3_lut6_2_O5 ;
wire [11:0] vec_out_r_AQ_0 ;
wire [11:1] vec_in_r_AQ_mux_0 ;
wire [11:0] vec_out_r_AQ_3 ;
wire [11:0] vec_in_r_AQ_mux_3 ;
wire [11:0] vec_out_r_AQ_2 ;
wire [11:0] vec_out_r_AQ_1 ;
wire [11:0] vec_in_r_AQ_mux_2 ;
wire [11:0] vec_in_r_AQ_mux_1 ;
wire [11:0] vec_out_i_AQ_0 ;
wire [11:0] vec_in_i_AQ_mux_0 ;
wire [11:0] vec_out_i_AQ_3 ;
wire [11:0] vec_in_i_AQ_mux_3 ;
wire [11:0] vec_out_i_AQ_2 ;
wire [11:0] vec_out_i_AQ_1 ;
wire [11:0] vec_in_i_AQ_mux_2 ;
wire [11:0] vec_in_i_AQ_mux_1 ;
wire [1:0] row_sel_AQ ;
wire [7:1] single_out_r_AQ2 ;
wire [11:0] single_out_i_AQ2 ;
wire [11:0] single_out_i_AQ ;
wire [8:1] single_out_r_AQ ;
wire [1:0] row_sel_R ;
wire col_sel_R_mux_i_m3_lut6_2_O6 ;
wire col_sel_R_mux_i_m3_lut6_2_O5 ;
wire [11:11] single_in_r_R_mux ;
wire wr_en_AQ_sel ;
wire [1:0] col_sel_R_int ;
wire [11:0] out_inner_prod_i ;
wire [11:0] out_inner_prod_r ;
wire in_a_inner_prod_sel ;
wire in_b_inner_prod_sel ;
wire [10:0] output_iv ;
wire [10:1] output_iv_0 ;
wire [11:11] out_r_vec_sub_0 ;
wire [11:11] out_i_vec_sub_0 ;
wire in_b_vec_mult_sel ;
wire [11:0] out_i_vec_mult_2 ;
wire [11:0] out_r_vec_mult_2 ;
wire [11:0] out_inv_sqrt ;
wire [11:0] out_i_vec_mult_1 ;
wire [11:0] out_r_vec_mult_1 ;
wire [11:0] out_i_vec_mult_0 ;
wire [11:0] out_r_vec_mult_0 ;
wire [11:0] out_i_vec_mult_3 ;
wire [11:0] out_r_vec_mult_3 ;
wire [11:11] in_a_r_reg_3 ;
wire [11:11] in_a_r_reg_2 ;
wire [11:11] in_a_r_reg_1 ;
wire [11:0] in_a_r_reg_0 ;
wire [11:11] in_a_i_reg_3 ;
wire [11:11] in_a_i_reg_2 ;
wire [11:11] in_a_i_reg_1 ;
wire [11:11] in_a_i_reg_0 ;
wire [22:1] pre_out ;
wire [10:0] pre_out_i_m ;
wire [11:1] pre_out_0 ;
wire [6:0] pre_out_i_m_0 ;
wire [11:1] pre_out_1 ;
wire [11:1] pre_out_2 ;
wire pre_out_i_m_1 ;
wire [11:2] pre_out_3 ;
wire [11:11] pre_out_4 ;
wire pre_out_i_m_2 ;
wire pre_out_i_m_3 ;
wire pre_out_i_m_4 ;
wire [11:11] pre_out_5 ;
wire [11:11] pre_out_6 ;
wire [10:0] un8_rnd_out ;
wire [19:19] un8_rnd_out_P ;
wire [23:23] pre_out_reg ;
wire single_in_R_sel ;
wire single_in_R_sel_0 ;
wire [1:0] w_col_sel_AQ_int ;
wire [1:0] col_sel_AQ2_int ;
wire [8:3] state ;
wire wr_en_AQ_sel_0 ;
wire [1:0] vec_in_AQ_sel ;
wire wr_en_AQ_mux_i_m3_lut6_2_O6 ;
wire N_507 ;
wire N_508 ;
wire N_505 ;
wire N_506 ;
wire N_645 ;
wire N_641 ;
wire N_637 ;
wire N_632 ;
wire N_628 ;
wire N_624 ;
wire N_623 ;
wire N_622 ;
wire N_612 ;
wire N_607 ;
wire N_606 ;
wire N_605 ;
wire N_597 ;
wire N_596 ;
wire N_595 ;
wire N_586 ;
wire N_585 ;
wire N_584 ;
wire N_583 ;
wire N_582 ;
wire N_571 ;
wire N_568 ;
wire N_567 ;
wire N_566 ;
wire N_555 ;
wire N_552 ;
wire N_549 ;
wire wr_en_R ;
wire N_28_i ;
wire N_30_i ;
wire N_32_i ;
wire N_34_i ;
wire N_383_i ;
wire N_384_i ;
wire N_385_i ;
wire N_386_i ;
wire N_387_i ;
wire N_388_i ;
wire N_389_i ;
wire N_390_i ;
wire N_391_i ;
wire N_392_i ;
wire N_393_i ;
wire N_394_i ;
wire N_395_i ;
wire N_396_i ;
wire N_397_i ;
wire N_398_i ;
wire N_399_i ;
wire N_400_i ;
wire N_401_i ;
wire start_inner_prod ;
wire red_mat_reg ;
wire done_inner_prod ;
wire N_501 ;
wire N_500 ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire w_in_a_vec_sub ;
wire un5_output ;
wire un5_output_0 ;
wire un5_output_1 ;
wire un5_output_2 ;
wire un5_output_3 ;
wire un5_output_4 ;
wire N_512_i ;
wire PATTERNDETECT_32 ;
wire done_inv_sqrt ;
wire start_inv_sqrt ;
wire wr_en_AQ_int ;
wire GND ;
wire VCC ;
input p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_ ;
input p_desc951_p_O_FDEinv_sqrt_ ;
input p_desc952_p_O_FDEinv_sqrt_ ;
input p_desc953_p_O_FDEinv_sqrt_ ;
input p_desc954_p_O_FDEinv_sqrt_ ;
input p_desc955_p_O_FDEinv_sqrt_ ;
input p_desc956_p_O_FDEinv_sqrt_ ;
input p_desc957_p_O_FDEinv_sqrt_ ;
input p_desc958_p_O_FDEinv_sqrt_ ;
input p_desc959_p_O_FDEinv_sqrt_ ;
input p_desc960_p_O_FDEinv_sqrt_ ;
input p_desc961_p_O_FDEinv_sqrt_ ;
input p_desc962_p_O_FDEinv_sqrt_ ;
input p_desc48_p_O_FDEr_mat_regs_ ;
input p_desc49_p_O_FDEr_mat_regs_ ;
input p_desc50_p_O_FDEr_mat_regs_ ;
input p_desc51_p_O_FDEr_mat_regs_ ;
input p_desc52_p_O_FDEr_mat_regs_ ;
input p_desc53_p_O_FDEr_mat_regs_ ;
input p_desc54_p_O_FDEr_mat_regs_ ;
input p_desc55_p_O_FDEr_mat_regs_ ;
input p_desc56_p_O_FDEr_mat_regs_ ;
input p_desc57_p_O_FDEr_mat_regs_ ;
input p_desc58_p_O_FDEr_mat_regs_ ;
input p_desc59_p_O_FDEr_mat_regs_ ;
input p_desc60_p_O_FDEr_mat_regs_ ;
input p_desc61_p_O_FDEr_mat_regs_ ;
input p_desc62_p_O_FDEr_mat_regs_ ;
input p_desc63_p_O_FDEr_mat_regs_ ;
input p_desc64_p_O_FDEr_mat_regs_ ;
input p_desc65_p_O_FDEr_mat_regs_ ;
input p_desc66_p_O_FDEr_mat_regs_ ;
input p_desc67_p_O_FDEr_mat_regs_ ;
input p_desc68_p_O_FDEr_mat_regs_ ;
input p_desc69_p_O_FDEr_mat_regs_ ;
input p_desc70_p_O_FDEr_mat_regs_ ;
input p_desc71_p_O_FDEr_mat_regs_ ;
input p_desc72_p_O_FDEr_mat_regs_ ;
input p_desc73_p_O_FDEr_mat_regs_ ;
input p_desc74_p_O_FDEr_mat_regs_ ;
input p_desc75_p_O_FDEr_mat_regs_ ;
input p_desc76_p_O_FDEr_mat_regs_ ;
input p_desc77_p_O_FDEr_mat_regs_ ;
input p_desc78_p_O_FDEr_mat_regs_ ;
input p_desc79_p_O_FDEr_mat_regs_ ;
input p_desc80_p_O_FDEr_mat_regs_ ;
input p_desc81_p_O_FDEr_mat_regs_ ;
input p_desc82_p_O_FDEr_mat_regs_ ;
input p_desc83_p_O_FDEr_mat_regs_ ;
input p_desc84_p_O_FDEr_mat_regs_ ;
input p_desc85_p_O_FDEr_mat_regs_ ;
input p_desc86_p_O_FDEr_mat_regs_ ;
input p_desc87_p_O_FDEr_mat_regs_ ;
input p_desc88_p_O_FDEr_mat_regs_ ;
input p_desc89_p_O_FDEr_mat_regs_ ;
input p_desc90_p_O_FDEr_mat_regs_ ;
input p_desc91_p_O_FDEr_mat_regs_ ;
input p_desc92_p_O_FDEr_mat_regs_ ;
input p_desc93_p_O_FDEr_mat_regs_ ;
input p_desc94_p_O_FDEr_mat_regs_ ;
input p_desc95_p_O_FDEr_mat_regs_ ;
input p_desc96_p_O_FDEr_mat_regs_ ;
input p_desc97_p_O_FDEr_mat_regs_ ;
input p_desc98_p_O_FDEr_mat_regs_ ;
input p_desc99_p_O_FDEr_mat_regs_ ;
input p_desc100_p_O_FDEr_mat_regs_ ;
input p_desc101_p_O_FDEr_mat_regs_ ;
input p_desc102_p_O_FDEr_mat_regs_ ;
input p_desc103_p_O_FDEr_mat_regs_ ;
input p_desc104_p_O_FDEr_mat_regs_ ;
input p_desc105_p_O_FDEr_mat_regs_ ;
input p_desc106_p_O_FDEr_mat_regs_ ;
input p_desc107_p_O_FDEr_mat_regs_ ;
input p_desc108_p_O_FDEr_mat_regs_ ;
input p_desc109_p_O_FDEr_mat_regs_ ;
input p_desc110_p_O_FDEr_mat_regs_ ;
input p_desc111_p_O_FDEr_mat_regs_ ;
input p_desc112_p_O_FDEr_mat_regs_ ;
input p_desc113_p_O_FDEr_mat_regs_ ;
input p_desc114_p_O_FDEr_mat_regs_ ;
input p_desc115_p_O_FDEr_mat_regs_ ;
input p_desc116_p_O_FDEr_mat_regs_ ;
input p_desc117_p_O_FDEr_mat_regs_ ;
input p_desc118_p_O_FDEr_mat_regs_ ;
input p_desc119_p_O_FDEr_mat_regs_ ;
input p_desc120_p_O_FDEr_mat_regs_ ;
input p_desc121_p_O_FDEr_mat_regs_ ;
input p_desc122_p_O_FDEr_mat_regs_ ;
input p_desc123_p_O_FDEr_mat_regs_ ;
input p_desc124_p_O_FDEr_mat_regs_ ;
input p_desc125_p_O_FDEr_mat_regs_ ;
input p_desc126_p_O_FDEr_mat_regs_ ;
input p_desc127_p_O_FDEr_mat_regs_ ;
input p_desc128_p_O_FDEr_mat_regs_ ;
input p_desc129_p_O_FDEr_mat_regs_ ;
input p_desc130_p_O_FDEr_mat_regs_ ;
input p_desc131_p_O_FDEr_mat_regs_ ;
input p_desc132_p_O_FDEr_mat_regs_ ;
input p_desc133_p_O_FDEr_mat_regs_ ;
input p_desc134_p_O_FDEr_mat_regs_ ;
input p_desc135_p_O_FDEr_mat_regs_ ;
input p_desc136_p_O_FDEr_mat_regs_ ;
input p_desc137_p_O_FDEr_mat_regs_ ;
input p_desc138_p_O_FDEr_mat_regs_ ;
input p_desc139_p_O_FDEr_mat_regs_ ;
input p_desc140_p_O_FDEr_mat_regs_ ;
input p_desc141_p_O_FDEr_mat_regs_ ;
input p_desc142_p_O_FDEr_mat_regs_ ;
input p_desc143_p_O_FDEr_mat_regs_ ;
input p_desc144_p_O_FDEr_mat_regs_ ;
input p_desc145_p_O_FDEr_mat_regs_ ;
input p_desc146_p_O_FDEr_mat_regs_ ;
input p_desc147_p_O_FDEr_mat_regs_ ;
input p_desc148_p_O_FDEr_mat_regs_ ;
input p_desc149_p_O_FDEr_mat_regs_ ;
input p_desc150_p_O_FDEr_mat_regs_ ;
input p_desc151_p_O_FDEr_mat_regs_ ;
input p_desc152_p_O_FDEr_mat_regs_ ;
input p_desc153_p_O_FDEr_mat_regs_ ;
input p_desc154_p_O_FDEr_mat_regs_ ;
input p_desc155_p_O_FDEr_mat_regs_ ;
input p_desc156_p_O_FDEr_mat_regs_ ;
input p_desc157_p_O_FDEr_mat_regs_ ;
input p_desc158_p_O_FDEr_mat_regs_ ;
input p_desc159_p_O_FDEr_mat_regs_ ;
input p_desc160_p_O_FDEr_mat_regs_ ;
input p_desc161_p_O_FDEr_mat_regs_ ;
input p_desc162_p_O_FDEr_mat_regs_ ;
input p_desc163_p_O_FDEr_mat_regs_ ;
input p_desc164_p_O_FDEr_mat_regs_ ;
input p_desc165_p_O_FDEr_mat_regs_ ;
input p_desc166_p_O_FDEr_mat_regs_ ;
input p_desc167_p_O_FDEr_mat_regs_ ;
input p_desc168_p_O_FDEr_mat_regs_ ;
input p_desc169_p_O_FDEr_mat_regs_ ;
input p_desc170_p_O_FDEr_mat_regs_ ;
input p_desc171_p_O_FDEr_mat_regs_ ;
input p_desc172_p_O_FDEr_mat_regs_ ;
input p_desc173_p_O_FDEr_mat_regs_ ;
input p_desc174_p_O_FDEr_mat_regs_ ;
input p_desc175_p_O_FDEr_mat_regs_ ;
input p_desc176_p_O_FDEr_mat_regs_ ;
input p_desc177_p_O_FDEr_mat_regs_ ;
input p_desc178_p_O_FDEr_mat_regs_ ;
input p_desc179_p_O_FDEr_mat_regs_ ;
input p_desc180_p_O_FDEr_mat_regs_ ;
input p_desc181_p_O_FDEr_mat_regs_ ;
input p_desc182_p_O_FDEr_mat_regs_ ;
input p_desc183_p_O_FDEr_mat_regs_ ;
input p_desc184_p_O_FDEr_mat_regs_ ;
input p_desc185_p_O_FDEr_mat_regs_ ;
input p_desc186_p_O_FDEr_mat_regs_ ;
input p_desc187_p_O_FDEr_mat_regs_ ;
input p_desc188_p_O_FDEr_mat_regs_ ;
input p_desc189_p_O_FDEr_mat_regs_ ;
input p_desc190_p_O_FDEr_mat_regs_ ;
input p_desc191_p_O_FDEr_mat_regs_ ;
input p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_ ;
input p_desc739_p_O_FDEvec_sub_ ;
input p_desc740_p_O_FDEvec_sub_ ;
input p_desc741_p_O_FDEvec_sub_ ;
input p_desc742_p_O_FDEvec_sub_ ;
input p_desc743_p_O_FDEvec_sub_ ;
input p_desc744_p_O_FDEvec_sub_ ;
input p_desc745_p_O_FDEvec_sub_ ;
input p_desc746_p_O_FDEvec_sub_ ;
input p_desc747_p_O_FDEvec_sub_ ;
input p_desc748_p_O_FDEvec_sub_ ;
input p_desc749_p_O_FDEvec_sub_ ;
input p_desc750_p_O_FDEvec_sub_ ;
input p_desc751_p_O_FDEvec_sub_ ;
input p_desc752_p_O_FDEvec_sub_ ;
input p_desc753_p_O_FDEvec_sub_ ;
input p_desc754_p_O_FDEvec_sub_ ;
input p_desc755_p_O_FDEvec_sub_ ;
input p_desc756_p_O_FDEvec_sub_ ;
input p_desc757_p_O_FDEvec_sub_ ;
input p_desc758_p_O_FDEvec_sub_ ;
input p_desc759_p_O_FDEvec_sub_ ;
input p_desc760_p_O_FDEvec_sub_ ;
input p_desc761_p_O_FDEvec_sub_ ;
input p_desc762_p_O_FDEvec_sub_ ;
input p_desc763_p_O_FDEvec_sub_ ;
input p_desc764_p_O_FDEvec_sub_ ;
input p_desc765_p_O_FDEvec_sub_ ;
input p_desc766_p_O_FDEvec_sub_ ;
input p_desc767_p_O_FDEvec_sub_ ;
input p_desc768_p_O_FDEvec_sub_ ;
input p_desc769_p_O_FDEvec_sub_ ;
input p_desc770_p_O_FDEvec_sub_ ;
input p_desc771_p_O_FDEvec_sub_ ;
input p_desc772_p_O_FDEvec_sub_ ;
input p_desc773_p_O_FDEvec_sub_ ;
input p_desc774_p_O_FDEvec_sub_ ;
input p_desc775_p_O_FDEvec_sub_ ;
input p_desc776_p_O_FDEvec_sub_ ;
input p_desc777_p_O_FDEvec_sub_ ;
input p_desc778_p_O_FDEvec_sub_ ;
input p_desc779_p_O_FDEvec_sub_ ;
input p_desc780_p_O_FDEvec_sub_ ;
input p_desc781_p_O_FDEvec_sub_ ;
input p_desc782_p_O_FDEvec_sub_ ;
input p_desc783_p_O_FDEvec_sub_ ;
input p_desc784_p_O_FDEvec_sub_ ;
input p_desc785_p_O_FDEvec_sub_ ;
input p_desc786_p_O_FDEvec_sub_ ;
input p_desc787_p_O_FDEvec_sub_ ;
input p_desc788_p_O_FDEvec_sub_ ;
input p_desc789_p_O_FDEvec_sub_ ;
input p_desc790_p_O_FDEvec_sub_ ;
input p_desc791_p_O_FDEvec_sub_ ;
input p_desc792_p_O_FDEvec_sub_ ;
input p_desc793_p_O_FDEvec_sub_ ;
input p_desc794_p_O_FDEvec_sub_ ;
input p_desc795_p_O_FDEvec_sub_ ;
input p_desc796_p_O_FDEvec_sub_ ;
input p_desc797_p_O_FDEvec_sub_ ;
input p_desc798_p_O_FDEvec_sub_ ;
input p_desc799_p_O_FDEvec_sub_ ;
input p_desc800_p_O_FDEvec_sub_ ;
input p_desc801_p_O_FDEvec_sub_ ;
input p_desc802_p_O_FDEvec_sub_ ;
input p_desc803_p_O_FDEvec_sub_ ;
input p_desc804_p_O_FDEvec_sub_ ;
input p_desc805_p_O_FDEvec_sub_ ;
input p_desc806_p_O_FDEvec_sub_ ;
input p_desc807_p_O_FDEvec_sub_ ;
input p_desc808_p_O_FDEvec_sub_ ;
input p_desc809_p_O_FDEvec_sub_ ;
input p_desc810_p_O_FDEvec_sub_ ;
input p_desc811_p_O_FDEvec_sub_ ;
input p_desc812_p_O_FDEvec_sub_ ;
input p_desc813_p_O_FDEvec_sub_ ;
input p_desc814_p_O_FDEvec_sub_ ;
input p_desc815_p_O_FDEvec_sub_ ;
input p_desc816_p_O_FDEvec_sub_ ;
input p_desc817_p_O_FDEvec_sub_ ;
input p_desc818_p_O_FDEvec_sub_ ;
input p_desc819_p_O_FDEvec_sub_ ;
input p_desc820_p_O_FDEvec_sub_ ;
input p_desc821_p_O_FDEvec_sub_ ;
input p_desc822_p_O_FDEvec_sub_ ;
input p_desc823_p_O_FDEvec_sub_ ;
input p_desc824_p_O_FDEvec_sub_ ;
input p_desc825_p_O_FDEvec_sub_ ;
input p_desc826_p_O_FDEvec_sub_ ;
input p_desc827_p_O_FDEvec_sub_ ;
input p_desc828_p_O_FDEvec_sub_ ;
input p_desc829_p_O_FDEvec_sub_ ;
input p_desc830_p_O_FDEvec_sub_ ;
input p_desc831_p_O_FDEvec_sub_ ;
input p_desc832_p_O_FDEvec_sub_ ;
input p_desc833_p_O_FDEvec_sub_ ;
input p_desc834_p_O_FDEvec_sub_ ;
input p_output_reg_pipe_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_ ;
input p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_ ;
input p_desc318_p_O_FDCinner_prod_ ;
input p_desc319_p_O_FDCinner_prod_ ;
input p_desc320_p_O_FDCinner_prod_ ;
input p_desc321_p_O_FDCinner_prod_ ;
input p_desc322_p_O_FDCinner_prod_ ;
input p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_ ;
input p_done_Z_p_O_FDCinner_prod_ ;
input p_acc_enable_Z_p_O_FDCinner_prod_ ;
input p_desc325_p_O_FDCinner_prod_ ;
input p_desc326_p_O_FDCinner_prod_ ;
input p_desc327_p_O_FDCinner_prod_ ;
input p_desc328_p_O_FDCinner_prod_ ;
input p_desc329_p_O_FDCinner_prod_ ;
input p_desc330_p_O_FDCinner_prod_ ;
input p_desc331_p_O_FDCinner_prod_ ;
input p_desc332_p_O_FDCinner_prod_ ;
input p_desc333_p_O_FDCinner_prod_ ;
input p_desc334_p_O_FDCinner_prod_ ;
input p_desc335_p_O_FDCinner_prod_ ;
input p_desc336_p_O_FDCinner_prod_ ;
input p_desc337_p_O_FDCinner_prod_ ;
input p_desc338_p_O_FDCinner_prod_ ;
input p_desc339_p_O_FDCinner_prod_ ;
input p_desc340_p_O_FDCinner_prod_ ;
input p_desc341_p_O_FDCinner_prod_ ;
input p_desc342_p_O_FDCinner_prod_ ;
input p_desc343_p_O_FDCinner_prod_ ;
input p_desc344_p_O_FDCinner_prod_ ;
input p_desc345_p_O_FDCinner_prod_ ;
input p_desc346_p_O_FDCinner_prod_ ;
input p_desc347_p_O_FDCinner_prod_ ;
input p_desc348_p_O_FDCinner_prod_ ;
input p_desc349_p_O_FDCinner_prod_ ;
input p_desc350_p_O_FDCinner_prod_ ;
input p_desc375_p_O_FDCinner_prod_ ;
input p_desc376_p_O_FDCinner_prod_ ;
input p_desc377_p_O_FDCinner_prod_ ;
input p_desc378_p_O_FDCinner_prod_ ;
input p_desc379_p_O_FDCinner_prod_ ;
input p_desc380_p_O_FDCinner_prod_ ;
input p_desc381_p_O_FDCinner_prod_ ;
input p_desc382_p_O_FDCinner_prod_ ;
input p_desc383_p_O_FDCinner_prod_ ;
input p_desc384_p_O_FDCinner_prod_ ;
input p_desc385_p_O_FDCinner_prod_ ;
input p_desc386_p_O_FDCinner_prod_ ;
input p_desc387_p_O_FDCinner_prod_ ;
input p_desc388_p_O_FDCinner_prod_ ;
input p_desc389_p_O_FDCinner_prod_ ;
input p_desc390_p_O_FDCinner_prod_ ;
input p_desc391_p_O_FDCinner_prod_ ;
input p_desc392_p_O_FDCinner_prod_ ;
input p_desc393_p_O_FDCinner_prod_ ;
input p_desc394_p_O_FDCinner_prod_ ;
input p_desc395_p_O_FDCinner_prod_ ;
input p_desc396_p_O_FDCinner_prod_ ;
input p_desc397_p_O_FDCinner_prod_ ;
input p_desc398_p_O_FDCinner_prod_ ;
input p_done_Z_p_O_FDCinv_sqrt_ ;
input p_desc946_p_O_FDCinv_sqrt_ ;
input p_desc947_p_O_FDCinv_sqrt_ ;
input p_desc948_p_O_FDCinv_sqrt_ ;
input p_desc949_p_O_FDCinv_sqrt_ ;
input p_desc950_p_O_FDCinv_sqrt_ ;
input p_desc1255_p_O_FDCqr_decomp_ctl_ ;
input p_desc1256_p_O_FDCqr_decomp_ctl_ ;
input p_desc1257_p_O_FDCqr_decomp_ctl_ ;
input p_desc1258_p_O_FDCqr_decomp_ctl_ ;
input p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_ ;
input p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_ ;
input p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_ ;
input p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_ ;
input p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_ ;
input p_desc1274_p_O_FDCqr_decomp_ctl_ ;
input p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_ ;
input p_done_Z_p_O_FDCqr_decomp_ctl_ ;
input p_desc1275_p_O_FDCqr_decomp_ctl_ ;
input p_desc1276_p_O_FDCqr_decomp_ctl_ ;
input p_desc1277_p_O_FDCqr_decomp_ctl_ ;
input p_desc1278_p_O_FDCqr_decomp_ctl_ ;
input p_desc1279_p_O_FDCqr_decomp_ctl_ ;
input p_desc1281_p_O_FDCqr_decomp_ctl_ ;
input p_desc1282_p_O_FDCqr_decomp_ctl_ ;
input p_desc1283_p_O_FDCqr_decomp_ctl_ ;
input p_desc1284_p_O_FDCqr_decomp_ctl_ ;
input p_desc1285_p_O_FDCqr_decomp_ctl_ ;
input p_desc1286_p_O_FDCqr_decomp_ctl_ ;
input p_desc1287_p_O_FDCqr_decomp_ctl_ ;
input p_desc1288_p_O_FDCqr_decomp_ctl_ ;
input p_acc_clear_Z_p_O_FDPinner_prod_ ;
input p_desc1265_p_O_FDPqr_decomp_ctl_ ;
input p_desc1268_p_O_FDPqr_decomp_ctl_ ;
input p_desc1280_p_O_FDPqr_decomp_ctl_ ;
input p_desc324_p_O_FDCEinner_prod_ ;
input p_desc351_p_O_FDCEinner_prod_ ;
input p_desc352_p_O_FDCEinner_prod_ ;
input p_desc353_p_O_FDCEinner_prod_ ;
input p_desc354_p_O_FDCEinner_prod_ ;
input p_desc355_p_O_FDCEinner_prod_ ;
input p_desc356_p_O_FDCEinner_prod_ ;
input p_desc357_p_O_FDCEinner_prod_ ;
input p_desc358_p_O_FDCEinner_prod_ ;
input p_desc359_p_O_FDCEinner_prod_ ;
input p_desc360_p_O_FDCEinner_prod_ ;
input p_desc361_p_O_FDCEinner_prod_ ;
input p_desc362_p_O_FDCEinner_prod_ ;
input p_desc363_p_O_FDCEinner_prod_ ;
input p_desc364_p_O_FDCEinner_prod_ ;
input p_desc365_p_O_FDCEinner_prod_ ;
input p_desc366_p_O_FDCEinner_prod_ ;
input p_desc367_p_O_FDCEinner_prod_ ;
input p_desc368_p_O_FDCEinner_prod_ ;
input p_desc369_p_O_FDCEinner_prod_ ;
input p_desc370_p_O_FDCEinner_prod_ ;
input p_desc371_p_O_FDCEinner_prod_ ;
input p_desc372_p_O_FDCEinner_prod_ ;
input p_desc373_p_O_FDCEinner_prod_ ;
input p_desc374_p_O_FDCEinner_prod_ ;
input p_desc1263_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1264_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1266_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1267_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1269_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1270_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1271_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1272_p_O_FDCEqr_decomp_ctl_ ;
input p_desc1273_p_O_FDCEqr_decomp_ctl_ ;
// instances
  mat_regs_inj A_Q_mat(.col_sel_AQ2_mux_i_m3_lut6_2_O6(col_sel_AQ2_mux_i_m3_lut6_2_O6),.col_sel_AQ2_mux_i_m3_lut6_2_O5(col_sel_AQ2_mux_i_m3_lut6_2_O5),.col_sel_AQ_int(col_sel_AQ_int[1:0]),.w_col_sel_AQ_mux_i_m3_lut6_2_O6(w_col_sel_AQ_mux_i_m3_lut6_2_O6),.w_col_sel_AQ_mux_i_m3_lut6_2_O5(w_col_sel_AQ_mux_i_m3_lut6_2_O5),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.vec_in_r_AQ_mux_0_4(vec_in_r_AQ_mux_0[5:5]),.vec_in_r_AQ_mux_0_9(vec_in_r_AQ_mux_0[10:10]),.vec_in_r_AQ_mux_0_6(vec_in_r_AQ_mux_0[7:7]),.vec_in_r_AQ_mux_0_0(vec_in_r_AQ_mux_0[1:1]),.vec_in_r_AQ_mux_0_1(vec_in_r_AQ_mux_0[2:2]),.vec_in_r_AQ_mux_0_2(vec_in_r_AQ_mux_0[3:3]),.vec_in_r_AQ_mux_0_3(vec_in_r_AQ_mux_0[4:4]),.vec_in_r_AQ_mux_0_10(vec_in_r_AQ_mux_0[11:11]),.vec_in_r_AQ_mux_0_7(vec_in_r_AQ_mux_0[8:8]),.vec_in_r_AQ_mux_0_8(vec_in_r_AQ_mux_0[9:9]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.vec_in_r_AQ_mux_3(vec_in_r_AQ_mux_3[11:0]),.out_Q_r(out_Q_r[47:0]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.vec_in_r_AQ_mux_2(vec_in_r_AQ_mux_2[11:0]),.vec_in_r_AQ_mux_1(vec_in_r_AQ_mux_1[11:0]),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.vec_in_i_AQ_mux_0_5(vec_in_i_AQ_mux_0[5:5]),.vec_in_i_AQ_mux_0_10(vec_in_i_AQ_mux_0[10:10]),.vec_in_i_AQ_mux_0_7(vec_in_i_AQ_mux_0[7:7]),.vec_in_i_AQ_mux_0_0(vec_in_i_AQ_mux_0[0:0]),.vec_in_i_AQ_mux_0_1(vec_in_i_AQ_mux_0[1:1]),.vec_in_i_AQ_mux_0_4(vec_in_i_AQ_mux_0[4:4]),.vec_in_i_AQ_mux_0_6(vec_in_i_AQ_mux_0[6:6]),.vec_in_i_AQ_mux_0_11(vec_in_i_AQ_mux_0[11:11]),.vec_in_i_AQ_mux_0_8(vec_in_i_AQ_mux_0[8:8]),.vec_in_i_AQ_mux_0_9(vec_in_i_AQ_mux_0[9:9]),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.vec_in_i_AQ_mux_3(vec_in_i_AQ_mux_3[11:0]),.out_Q_i(out_Q_i[47:0]),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.vec_in_i_AQ_mux_2(vec_in_i_AQ_mux_2[11:0]),.vec_in_i_AQ_mux_1(vec_in_i_AQ_mux_1[11:0]),.row_sel_AQ(row_sel_AQ[1:0]),.single_out_r_AQ2_1(single_out_r_AQ2[2:2]),.single_out_r_AQ2_6(single_out_r_AQ2[7:7]),.single_out_r_AQ2_4(single_out_r_AQ2[5:5]),.single_out_r_AQ2_0(single_out_r_AQ2[1:1]),.single_out_i_AQ2_1(single_out_i_AQ2[1:1]),.single_out_i_AQ2_5(single_out_i_AQ2[5:5]),.single_out_i_AQ2_4(single_out_i_AQ2[4:4]),.single_out_i_AQ2_0(single_out_i_AQ2[0:0]),.single_out_i_AQ2_11(single_out_i_AQ2[11:11]),.single_out_i_AQ_1(single_out_i_AQ[1:1]),.single_out_i_AQ_0(single_out_i_AQ[0:0]),.single_out_i_AQ_8(single_out_i_AQ[8:8]),.single_out_i_AQ_10(single_out_i_AQ[10:10]),.single_out_i_AQ_11(single_out_i_AQ[11:11]),.single_out_i_AQ_9(single_out_i_AQ[9:9]),.single_out_i_AQ_4(single_out_i_AQ[4:4]),.single_out_r_AQ_4(single_out_r_AQ[5:5]),.single_out_r_AQ_2(single_out_r_AQ[3:3]),.single_out_r_AQ_7(single_out_r_AQ[8:8]),.single_out_r_AQ_1(single_out_r_AQ[2:2]),.single_out_r_AQ_0(single_out_r_AQ[1:1]),.clk(clk),.wr_en_AQ_mux_i_m3_lut6_2_O6(wr_en_AQ_mux_i_m3_lut6_2_O6),.N_507(N_507),.N_508(N_508),.N_505(N_505),.N_506(N_506),.N_645(N_645),.N_641(N_641),.N_637(N_637),.N_632(N_632),.N_628(N_628),.N_624(N_624),.N_623(N_623),.N_622(N_622),.N_612(N_612),.N_607(N_607),.N_606(N_606),.N_605(N_605),.N_597(N_597),.N_596(N_596),.N_595(N_595),.N_586(N_586),.N_585(N_585),.N_584(N_584),.N_583(N_583),.N_582(N_582),.N_571(N_571),.N_568(N_568),.N_567(N_567),.N_566(N_566),.N_555(N_555),.N_552(N_552),.N_549(N_549));
  r_mat_regs_inj R_mat(.row_sel_R(row_sel_R[1:0]),.col_sel_R_mux_i_m3_lut6_2_O6(col_sel_R_mux_i_m3_lut6_2_O6),.col_sel_R_mux_i_m3_lut6_2_O5(col_sel_R_mux_i_m3_lut6_2_O5),.single_in_r_R_mux(single_in_r_R_mux[11:11]),.wr_en_AQ_sel(wr_en_AQ_sel),.col_sel_R(col_sel_R[1:0]),.col_sel_R_int(col_sel_R_int[1:0]),.out_R_i(out_R_i[47:12]),.out_R_r(out_R_r[47:0]),.wr_en_R(wr_en_R),.N_28_i(N_28_i),.clk(clk),.N_30_i(N_30_i),.N_32_i(N_32_i),.N_34_i(N_34_i),.N_383_i(N_383_i),.N_384_i(N_384_i),.N_385_i(N_385_i),.N_386_i(N_386_i),.N_387_i(N_387_i),.N_388_i(N_388_i),.N_389_i(N_389_i),.N_390_i(N_390_i),.N_391_i(N_391_i),.N_392_i(N_392_i),.N_393_i(N_393_i),.N_394_i(N_394_i),.N_395_i(N_395_i),.N_396_i(N_396_i),.N_397_i(N_397_i),.N_398_i(N_398_i),.N_399_i(N_399_i),.N_400_i(N_400_i),.N_401_i(N_401_i),.p_desc48_p_O_FDE(p_desc48_p_O_FDEr_mat_regs_),.p_desc49_p_O_FDE(p_desc49_p_O_FDEr_mat_regs_),.p_desc50_p_O_FDE(p_desc50_p_O_FDEr_mat_regs_),.p_desc51_p_O_FDE(p_desc51_p_O_FDEr_mat_regs_),.p_desc52_p_O_FDE(p_desc52_p_O_FDEr_mat_regs_),.p_desc53_p_O_FDE(p_desc53_p_O_FDEr_mat_regs_),.p_desc54_p_O_FDE(p_desc54_p_O_FDEr_mat_regs_),.p_desc55_p_O_FDE(p_desc55_p_O_FDEr_mat_regs_),.p_desc56_p_O_FDE(p_desc56_p_O_FDEr_mat_regs_),.p_desc57_p_O_FDE(p_desc57_p_O_FDEr_mat_regs_),.p_desc58_p_O_FDE(p_desc58_p_O_FDEr_mat_regs_),.p_desc59_p_O_FDE(p_desc59_p_O_FDEr_mat_regs_),.p_desc60_p_O_FDE(p_desc60_p_O_FDEr_mat_regs_),.p_desc61_p_O_FDE(p_desc61_p_O_FDEr_mat_regs_),.p_desc62_p_O_FDE(p_desc62_p_O_FDEr_mat_regs_),.p_desc63_p_O_FDE(p_desc63_p_O_FDEr_mat_regs_),.p_desc64_p_O_FDE(p_desc64_p_O_FDEr_mat_regs_),.p_desc65_p_O_FDE(p_desc65_p_O_FDEr_mat_regs_),.p_desc66_p_O_FDE(p_desc66_p_O_FDEr_mat_regs_),.p_desc67_p_O_FDE(p_desc67_p_O_FDEr_mat_regs_),.p_desc68_p_O_FDE(p_desc68_p_O_FDEr_mat_regs_),.p_desc69_p_O_FDE(p_desc69_p_O_FDEr_mat_regs_),.p_desc70_p_O_FDE(p_desc70_p_O_FDEr_mat_regs_),.p_desc71_p_O_FDE(p_desc71_p_O_FDEr_mat_regs_),.p_desc72_p_O_FDE(p_desc72_p_O_FDEr_mat_regs_),.p_desc73_p_O_FDE(p_desc73_p_O_FDEr_mat_regs_),.p_desc74_p_O_FDE(p_desc74_p_O_FDEr_mat_regs_),.p_desc75_p_O_FDE(p_desc75_p_O_FDEr_mat_regs_),.p_desc76_p_O_FDE(p_desc76_p_O_FDEr_mat_regs_),.p_desc77_p_O_FDE(p_desc77_p_O_FDEr_mat_regs_),.p_desc78_p_O_FDE(p_desc78_p_O_FDEr_mat_regs_),.p_desc79_p_O_FDE(p_desc79_p_O_FDEr_mat_regs_),.p_desc80_p_O_FDE(p_desc80_p_O_FDEr_mat_regs_),.p_desc81_p_O_FDE(p_desc81_p_O_FDEr_mat_regs_),.p_desc82_p_O_FDE(p_desc82_p_O_FDEr_mat_regs_),.p_desc83_p_O_FDE(p_desc83_p_O_FDEr_mat_regs_),.p_desc84_p_O_FDE(p_desc84_p_O_FDEr_mat_regs_),.p_desc85_p_O_FDE(p_desc85_p_O_FDEr_mat_regs_),.p_desc86_p_O_FDE(p_desc86_p_O_FDEr_mat_regs_),.p_desc87_p_O_FDE(p_desc87_p_O_FDEr_mat_regs_),.p_desc88_p_O_FDE(p_desc88_p_O_FDEr_mat_regs_),.p_desc89_p_O_FDE(p_desc89_p_O_FDEr_mat_regs_),.p_desc90_p_O_FDE(p_desc90_p_O_FDEr_mat_regs_),.p_desc91_p_O_FDE(p_desc91_p_O_FDEr_mat_regs_),.p_desc92_p_O_FDE(p_desc92_p_O_FDEr_mat_regs_),.p_desc93_p_O_FDE(p_desc93_p_O_FDEr_mat_regs_),.p_desc94_p_O_FDE(p_desc94_p_O_FDEr_mat_regs_),.p_desc95_p_O_FDE(p_desc95_p_O_FDEr_mat_regs_),.p_desc96_p_O_FDE(p_desc96_p_O_FDEr_mat_regs_),.p_desc97_p_O_FDE(p_desc97_p_O_FDEr_mat_regs_),.p_desc98_p_O_FDE(p_desc98_p_O_FDEr_mat_regs_),.p_desc99_p_O_FDE(p_desc99_p_O_FDEr_mat_regs_),.p_desc100_p_O_FDE(p_desc100_p_O_FDEr_mat_regs_),.p_desc101_p_O_FDE(p_desc101_p_O_FDEr_mat_regs_),.p_desc102_p_O_FDE(p_desc102_p_O_FDEr_mat_regs_),.p_desc103_p_O_FDE(p_desc103_p_O_FDEr_mat_regs_),.p_desc104_p_O_FDE(p_desc104_p_O_FDEr_mat_regs_),.p_desc105_p_O_FDE(p_desc105_p_O_FDEr_mat_regs_),.p_desc106_p_O_FDE(p_desc106_p_O_FDEr_mat_regs_),.p_desc107_p_O_FDE(p_desc107_p_O_FDEr_mat_regs_),.p_desc108_p_O_FDE(p_desc108_p_O_FDEr_mat_regs_),.p_desc109_p_O_FDE(p_desc109_p_O_FDEr_mat_regs_),.p_desc110_p_O_FDE(p_desc110_p_O_FDEr_mat_regs_),.p_desc111_p_O_FDE(p_desc111_p_O_FDEr_mat_regs_),.p_desc112_p_O_FDE(p_desc112_p_O_FDEr_mat_regs_),.p_desc113_p_O_FDE(p_desc113_p_O_FDEr_mat_regs_),.p_desc114_p_O_FDE(p_desc114_p_O_FDEr_mat_regs_),.p_desc115_p_O_FDE(p_desc115_p_O_FDEr_mat_regs_),.p_desc116_p_O_FDE(p_desc116_p_O_FDEr_mat_regs_),.p_desc117_p_O_FDE(p_desc117_p_O_FDEr_mat_regs_),.p_desc118_p_O_FDE(p_desc118_p_O_FDEr_mat_regs_),.p_desc119_p_O_FDE(p_desc119_p_O_FDEr_mat_regs_),.p_desc120_p_O_FDE(p_desc120_p_O_FDEr_mat_regs_),.p_desc121_p_O_FDE(p_desc121_p_O_FDEr_mat_regs_),.p_desc122_p_O_FDE(p_desc122_p_O_FDEr_mat_regs_),.p_desc123_p_O_FDE(p_desc123_p_O_FDEr_mat_regs_),.p_desc124_p_O_FDE(p_desc124_p_O_FDEr_mat_regs_),.p_desc125_p_O_FDE(p_desc125_p_O_FDEr_mat_regs_),.p_desc126_p_O_FDE(p_desc126_p_O_FDEr_mat_regs_),.p_desc127_p_O_FDE(p_desc127_p_O_FDEr_mat_regs_),.p_desc128_p_O_FDE(p_desc128_p_O_FDEr_mat_regs_),.p_desc129_p_O_FDE(p_desc129_p_O_FDEr_mat_regs_),.p_desc130_p_O_FDE(p_desc130_p_O_FDEr_mat_regs_),.p_desc131_p_O_FDE(p_desc131_p_O_FDEr_mat_regs_),.p_desc132_p_O_FDE(p_desc132_p_O_FDEr_mat_regs_),.p_desc133_p_O_FDE(p_desc133_p_O_FDEr_mat_regs_),.p_desc134_p_O_FDE(p_desc134_p_O_FDEr_mat_regs_),.p_desc135_p_O_FDE(p_desc135_p_O_FDEr_mat_regs_),.p_desc136_p_O_FDE(p_desc136_p_O_FDEr_mat_regs_),.p_desc137_p_O_FDE(p_desc137_p_O_FDEr_mat_regs_),.p_desc138_p_O_FDE(p_desc138_p_O_FDEr_mat_regs_),.p_desc139_p_O_FDE(p_desc139_p_O_FDEr_mat_regs_),.p_desc140_p_O_FDE(p_desc140_p_O_FDEr_mat_regs_),.p_desc141_p_O_FDE(p_desc141_p_O_FDEr_mat_regs_),.p_desc142_p_O_FDE(p_desc142_p_O_FDEr_mat_regs_),.p_desc143_p_O_FDE(p_desc143_p_O_FDEr_mat_regs_),.p_desc144_p_O_FDE(p_desc144_p_O_FDEr_mat_regs_),.p_desc145_p_O_FDE(p_desc145_p_O_FDEr_mat_regs_),.p_desc146_p_O_FDE(p_desc146_p_O_FDEr_mat_regs_),.p_desc147_p_O_FDE(p_desc147_p_O_FDEr_mat_regs_),.p_desc148_p_O_FDE(p_desc148_p_O_FDEr_mat_regs_),.p_desc149_p_O_FDE(p_desc149_p_O_FDEr_mat_regs_),.p_desc150_p_O_FDE(p_desc150_p_O_FDEr_mat_regs_),.p_desc151_p_O_FDE(p_desc151_p_O_FDEr_mat_regs_),.p_desc152_p_O_FDE(p_desc152_p_O_FDEr_mat_regs_),.p_desc153_p_O_FDE(p_desc153_p_O_FDEr_mat_regs_),.p_desc154_p_O_FDE(p_desc154_p_O_FDEr_mat_regs_),.p_desc155_p_O_FDE(p_desc155_p_O_FDEr_mat_regs_),.p_desc156_p_O_FDE(p_desc156_p_O_FDEr_mat_regs_),.p_desc157_p_O_FDE(p_desc157_p_O_FDEr_mat_regs_),.p_desc158_p_O_FDE(p_desc158_p_O_FDEr_mat_regs_),.p_desc159_p_O_FDE(p_desc159_p_O_FDEr_mat_regs_),.p_desc160_p_O_FDE(p_desc160_p_O_FDEr_mat_regs_),.p_desc161_p_O_FDE(p_desc161_p_O_FDEr_mat_regs_),.p_desc162_p_O_FDE(p_desc162_p_O_FDEr_mat_regs_),.p_desc163_p_O_FDE(p_desc163_p_O_FDEr_mat_regs_),.p_desc164_p_O_FDE(p_desc164_p_O_FDEr_mat_regs_),.p_desc165_p_O_FDE(p_desc165_p_O_FDEr_mat_regs_),.p_desc166_p_O_FDE(p_desc166_p_O_FDEr_mat_regs_),.p_desc167_p_O_FDE(p_desc167_p_O_FDEr_mat_regs_),.p_desc168_p_O_FDE(p_desc168_p_O_FDEr_mat_regs_),.p_desc169_p_O_FDE(p_desc169_p_O_FDEr_mat_regs_),.p_desc170_p_O_FDE(p_desc170_p_O_FDEr_mat_regs_),.p_desc171_p_O_FDE(p_desc171_p_O_FDEr_mat_regs_),.p_desc172_p_O_FDE(p_desc172_p_O_FDEr_mat_regs_),.p_desc173_p_O_FDE(p_desc173_p_O_FDEr_mat_regs_),.p_desc174_p_O_FDE(p_desc174_p_O_FDEr_mat_regs_),.p_desc175_p_O_FDE(p_desc175_p_O_FDEr_mat_regs_),.p_desc176_p_O_FDE(p_desc176_p_O_FDEr_mat_regs_),.p_desc177_p_O_FDE(p_desc177_p_O_FDEr_mat_regs_),.p_desc178_p_O_FDE(p_desc178_p_O_FDEr_mat_regs_),.p_desc179_p_O_FDE(p_desc179_p_O_FDEr_mat_regs_),.p_desc180_p_O_FDE(p_desc180_p_O_FDEr_mat_regs_),.p_desc181_p_O_FDE(p_desc181_p_O_FDEr_mat_regs_),.p_desc182_p_O_FDE(p_desc182_p_O_FDEr_mat_regs_),.p_desc183_p_O_FDE(p_desc183_p_O_FDEr_mat_regs_),.p_desc184_p_O_FDE(p_desc184_p_O_FDEr_mat_regs_),.p_desc185_p_O_FDE(p_desc185_p_O_FDEr_mat_regs_),.p_desc186_p_O_FDE(p_desc186_p_O_FDEr_mat_regs_),.p_desc187_p_O_FDE(p_desc187_p_O_FDEr_mat_regs_),.p_desc188_p_O_FDE(p_desc188_p_O_FDEr_mat_regs_),.p_desc189_p_O_FDE(p_desc189_p_O_FDEr_mat_regs_),.p_desc190_p_O_FDE(p_desc190_p_O_FDEr_mat_regs_),.p_desc191_p_O_FDE(p_desc191_p_O_FDEr_mat_regs_));
  inner_prod_inj inner_prod_inst(.out_inner_prod_i(out_inner_prod_i[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.in_a_inner_prod_sel(in_a_inner_prod_sel),.single_out_r_AQ_7(single_out_r_AQ[8:8]),.single_out_r_AQ_0(single_out_r_AQ[1:1]),.single_out_r_AQ_1(single_out_r_AQ[2:2]),.single_out_r_AQ_4(single_out_r_AQ[5:5]),.single_out_r_AQ_2(single_out_r_AQ[3:3]),.in_b_inner_prod_sel(in_b_inner_prod_sel),.vec_in_r_AQ_mux_0_6(vec_in_r_AQ_mux_0[7:7]),.vec_in_r_AQ_mux_0_7(vec_in_r_AQ_mux_0[8:8]),.vec_in_r_AQ_mux_0_0(vec_in_r_AQ_mux_0[1:1]),.vec_in_r_AQ_mux_0_9(vec_in_r_AQ_mux_0[10:10]),.vec_in_r_AQ_mux_0_1(vec_in_r_AQ_mux_0[2:2]),.vec_in_r_AQ_mux_0_8(vec_in_r_AQ_mux_0[9:9]),.vec_in_r_AQ_mux_0_4(vec_in_r_AQ_mux_0[5:5]),.vec_in_r_AQ_mux_0_3(vec_in_r_AQ_mux_0[4:4]),.vec_in_r_AQ_mux_0_2(vec_in_r_AQ_mux_0[3:3]),.vec_in_r_AQ_mux_0_10(vec_in_r_AQ_mux_0[11:11]),.vec_in_i_AQ_mux_0_7(vec_in_i_AQ_mux_0[7:7]),.vec_in_i_AQ_mux_0_1(vec_in_i_AQ_mux_0[1:1]),.vec_in_i_AQ_mux_0_0(vec_in_i_AQ_mux_0[0:0]),.vec_in_i_AQ_mux_0_6(vec_in_i_AQ_mux_0[6:6]),.vec_in_i_AQ_mux_0_8(vec_in_i_AQ_mux_0[8:8]),.vec_in_i_AQ_mux_0_10(vec_in_i_AQ_mux_0[10:10]),.vec_in_i_AQ_mux_0_5(vec_in_i_AQ_mux_0[5:5]),.vec_in_i_AQ_mux_0_9(vec_in_i_AQ_mux_0[9:9]),.vec_in_i_AQ_mux_0_4(vec_in_i_AQ_mux_0[4:4]),.vec_in_i_AQ_mux_0_11(vec_in_i_AQ_mux_0[11:11]),.single_out_i_AQ_1(single_out_i_AQ[1:1]),.single_out_i_AQ_0(single_out_i_AQ[0:0]),.single_out_i_AQ_8(single_out_i_AQ[8:8]),.single_out_i_AQ_10(single_out_i_AQ[10:10]),.single_out_i_AQ_9(single_out_i_AQ[9:9]),.single_out_i_AQ_4(single_out_i_AQ[4:4]),.single_out_i_AQ_11(single_out_i_AQ[11:11]),.output_iv(output_iv[10:0]),.single_out_r_AQ2_4(single_out_r_AQ2[5:5]),.single_out_r_AQ2_0(single_out_r_AQ2[1:1]),.single_out_r_AQ2_1(single_out_r_AQ2[2:2]),.single_out_r_AQ2_6(single_out_r_AQ2[7:7]),.output_iv_0_4(output_iv_0[5:5]),.output_iv_0_7(output_iv_0[8:8]),.output_iv_0_0(output_iv_0[1:1]),.output_iv_0_9(output_iv_0[10:10]),.output_iv_0_1(output_iv_0[2:2]),.output_iv_0_6(output_iv_0[7:7]),.output_iv_0_3(output_iv_0[4:4]),.output_iv_0_2(output_iv_0[3:3]),.output_iv_0_8(output_iv_0[9:9]),.out_r_vec_sub_0(out_r_vec_sub_0[11:11]),.out_i_vec_sub_0(out_i_vec_sub_0[11:11]),.single_out_i_AQ2_0(single_out_i_AQ2[0:0]),.single_out_i_AQ2_5(single_out_i_AQ2[5:5]),.single_out_i_AQ2_4(single_out_i_AQ2[4:4]),.single_out_i_AQ2_1(single_out_i_AQ2[1:1]),.single_out_i_AQ2_11(single_out_i_AQ2[11:11]),.start_inner_prod(start_inner_prod),.red_mat_reg(red_mat_reg),.clk(clk),.rst(rst),.done_inner_prod(done_inner_prod),.N_623(N_623),.N_568(N_568),.N_622(N_622),.N_507(N_507),.N_549(N_549),.N_505(N_505),.N_597(N_597),.N_567(N_567),.N_596(N_596),.N_628(N_628),.N_637(N_637),.N_566(N_566),.N_506(N_506),.N_585(N_585),.N_584(N_584),.N_612(N_612),.N_583(N_583),.N_595(N_595),.N_508(N_508),.N_501(N_501),.N_605(N_605),.N_624(N_624),.N_607(N_607),.N_552(N_552),.N_555(N_555),.N_586(N_586),.N_645(N_645),.N_641(N_641),.N_582(N_582),.N_606(N_606),.N_632(N_632),.N_500(N_500),.N_571(N_571),.p_desc318_p_O_FDC(p_desc318_p_O_FDCinner_prod_),.p_desc319_p_O_FDC(p_desc319_p_O_FDCinner_prod_),.p_desc320_p_O_FDC(p_desc320_p_O_FDCinner_prod_),.p_desc321_p_O_FDC(p_desc321_p_O_FDCinner_prod_),.p_desc322_p_O_FDC(p_desc322_p_O_FDCinner_prod_),.p_in_reg_enable_fsm_Z_p_O_FDC(p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_),.p_done_Z_p_O_FDC(p_done_Z_p_O_FDCinner_prod_),.p_acc_enable_Z_p_O_FDC(p_acc_enable_Z_p_O_FDCinner_prod_),.p_desc325_p_O_FDC(p_desc325_p_O_FDCinner_prod_),.p_desc326_p_O_FDC(p_desc326_p_O_FDCinner_prod_),.p_desc327_p_O_FDC(p_desc327_p_O_FDCinner_prod_),.p_desc328_p_O_FDC(p_desc328_p_O_FDCinner_prod_),.p_desc329_p_O_FDC(p_desc329_p_O_FDCinner_prod_),.p_desc330_p_O_FDC(p_desc330_p_O_FDCinner_prod_),.p_desc331_p_O_FDC(p_desc331_p_O_FDCinner_prod_),.p_desc332_p_O_FDC(p_desc332_p_O_FDCinner_prod_),.p_desc333_p_O_FDC(p_desc333_p_O_FDCinner_prod_),.p_desc334_p_O_FDC(p_desc334_p_O_FDCinner_prod_),.p_desc335_p_O_FDC(p_desc335_p_O_FDCinner_prod_),.p_desc336_p_O_FDC(p_desc336_p_O_FDCinner_prod_),.p_desc337_p_O_FDC(p_desc337_p_O_FDCinner_prod_),.p_desc338_p_O_FDC(p_desc338_p_O_FDCinner_prod_),.p_desc339_p_O_FDC(p_desc339_p_O_FDCinner_prod_),.p_desc340_p_O_FDC(p_desc340_p_O_FDCinner_prod_),.p_desc341_p_O_FDC(p_desc341_p_O_FDCinner_prod_),.p_desc342_p_O_FDC(p_desc342_p_O_FDCinner_prod_),.p_desc343_p_O_FDC(p_desc343_p_O_FDCinner_prod_),.p_desc344_p_O_FDC(p_desc344_p_O_FDCinner_prod_),.p_desc345_p_O_FDC(p_desc345_p_O_FDCinner_prod_),.p_desc346_p_O_FDC(p_desc346_p_O_FDCinner_prod_),.p_desc347_p_O_FDC(p_desc347_p_O_FDCinner_prod_),.p_desc348_p_O_FDC(p_desc348_p_O_FDCinner_prod_),.p_desc349_p_O_FDC(p_desc349_p_O_FDCinner_prod_),.p_desc350_p_O_FDC(p_desc350_p_O_FDCinner_prod_),.p_desc375_p_O_FDC(p_desc375_p_O_FDCinner_prod_),.p_desc376_p_O_FDC(p_desc376_p_O_FDCinner_prod_),.p_desc377_p_O_FDC(p_desc377_p_O_FDCinner_prod_),.p_desc378_p_O_FDC(p_desc378_p_O_FDCinner_prod_),.p_desc379_p_O_FDC(p_desc379_p_O_FDCinner_prod_),.p_desc380_p_O_FDC(p_desc380_p_O_FDCinner_prod_),.p_desc381_p_O_FDC(p_desc381_p_O_FDCinner_prod_),.p_desc382_p_O_FDC(p_desc382_p_O_FDCinner_prod_),.p_desc383_p_O_FDC(p_desc383_p_O_FDCinner_prod_),.p_desc384_p_O_FDC(p_desc384_p_O_FDCinner_prod_),.p_desc385_p_O_FDC(p_desc385_p_O_FDCinner_prod_),.p_desc386_p_O_FDC(p_desc386_p_O_FDCinner_prod_),.p_desc387_p_O_FDC(p_desc387_p_O_FDCinner_prod_),.p_desc388_p_O_FDC(p_desc388_p_O_FDCinner_prod_),.p_desc389_p_O_FDC(p_desc389_p_O_FDCinner_prod_),.p_desc390_p_O_FDC(p_desc390_p_O_FDCinner_prod_),.p_desc391_p_O_FDC(p_desc391_p_O_FDCinner_prod_),.p_desc392_p_O_FDC(p_desc392_p_O_FDCinner_prod_),.p_desc393_p_O_FDC(p_desc393_p_O_FDCinner_prod_),.p_desc394_p_O_FDC(p_desc394_p_O_FDCinner_prod_),.p_desc395_p_O_FDC(p_desc395_p_O_FDCinner_prod_),.p_desc396_p_O_FDC(p_desc396_p_O_FDCinner_prod_),.p_desc397_p_O_FDC(p_desc397_p_O_FDCinner_prod_),.p_desc398_p_O_FDC(p_desc398_p_O_FDCinner_prod_),.p_acc_clear_Z_p_O_FDP(p_acc_clear_Z_p_O_FDPinner_prod_),.p_desc324_p_O_FDCE(p_desc324_p_O_FDCEinner_prod_),.p_desc351_p_O_FDCE(p_desc351_p_O_FDCEinner_prod_),.p_desc352_p_O_FDCE(p_desc352_p_O_FDCEinner_prod_),.p_desc353_p_O_FDCE(p_desc353_p_O_FDCEinner_prod_),.p_desc354_p_O_FDCE(p_desc354_p_O_FDCEinner_prod_),.p_desc355_p_O_FDCE(p_desc355_p_O_FDCEinner_prod_),.p_desc356_p_O_FDCE(p_desc356_p_O_FDCEinner_prod_),.p_desc357_p_O_FDCE(p_desc357_p_O_FDCEinner_prod_),.p_desc358_p_O_FDCE(p_desc358_p_O_FDCEinner_prod_),.p_desc359_p_O_FDCE(p_desc359_p_O_FDCEinner_prod_),.p_desc360_p_O_FDCE(p_desc360_p_O_FDCEinner_prod_),.p_desc361_p_O_FDCE(p_desc361_p_O_FDCEinner_prod_),.p_desc362_p_O_FDCE(p_desc362_p_O_FDCEinner_prod_),.p_desc363_p_O_FDCE(p_desc363_p_O_FDCEinner_prod_),.p_desc364_p_O_FDCE(p_desc364_p_O_FDCEinner_prod_),.p_desc365_p_O_FDCE(p_desc365_p_O_FDCEinner_prod_),.p_desc366_p_O_FDCE(p_desc366_p_O_FDCEinner_prod_),.p_desc367_p_O_FDCE(p_desc367_p_O_FDCEinner_prod_),.p_desc368_p_O_FDCE(p_desc368_p_O_FDCEinner_prod_),.p_desc369_p_O_FDCE(p_desc369_p_O_FDCEinner_prod_),.p_desc370_p_O_FDCE(p_desc370_p_O_FDCEinner_prod_),.p_desc371_p_O_FDCE(p_desc371_p_O_FDCEinner_prod_),.p_desc372_p_O_FDCE(p_desc372_p_O_FDCEinner_prod_),.p_desc373_p_O_FDCE(p_desc373_p_O_FDCEinner_prod_),.p_desc374_p_O_FDCE(p_desc374_p_O_FDCEinner_prod_));
  vec_mult_inj vec_mult_inst(.in_b_vec_mult_sel(in_b_vec_mult_sel),.out_inner_prod_i(out_inner_prod_i[11:0]),.out_i_vec_mult_2(out_i_vec_mult_2[11:0]),.out_r_vec_mult_2(out_r_vec_mult_2[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.out_inv_sqrt_0(out_inv_sqrt[0:0]),.out_inv_sqrt_1(out_inv_sqrt[1:1]),.out_inv_sqrt_2(out_inv_sqrt[2:2]),.out_inv_sqrt_7(out_inv_sqrt[7:7]),.out_inv_sqrt_8(out_inv_sqrt[8:8]),.out_inv_sqrt_9(out_inv_sqrt[9:9]),.out_inv_sqrt_10(out_inv_sqrt[10:10]),.out_inv_sqrt_11(out_inv_sqrt[11:11]),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.out_i_vec_mult_1(out_i_vec_mult_1[11:0]),.out_r_vec_mult_1(out_r_vec_mult_1[11:0]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.out_i_vec_mult_0(out_i_vec_mult_0[11:0]),.out_r_vec_mult_0(out_r_vec_mult_0[11:0]),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.out_i_vec_mult_3(out_i_vec_mult_3[11:0]),.out_r_vec_mult_3(out_r_vec_mult_3[11:0]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  vec_sub_inj vec_sub_inst(.in_a_r_reg_3_11(in_a_r_reg_3[11:11]),.in_a_r_reg_2_11(in_a_r_reg_2[11:11]),.in_a_r_reg_1_11(in_a_r_reg_1[11:11]),.in_a_r_reg_0_0(in_a_r_reg_0[0:0]),.in_a_r_reg_0_11(in_a_r_reg_0[11:11]),.out_Q_r(out_Q_r[47:0]),.in_a_i_reg_3_11(in_a_i_reg_3[11:11]),.in_a_i_reg_2_11(in_a_i_reg_2[11:11]),.in_a_i_reg_1_11(in_a_i_reg_1[11:11]),.in_a_i_reg_0_11(in_a_i_reg_0[11:11]),.out_Q_i(out_Q_i[47:0]),.out_r_vec_mult_0(out_r_vec_mult_0[11:0]),.out_r_vec_mult_1(out_r_vec_mult_1[11:0]),.out_r_vec_mult_2(out_r_vec_mult_2[11:0]),.pre_out(pre_out[11:1]),.out_r_vec_mult_3(out_r_vec_mult_3[11:0]),.pre_out_i_m_1(pre_out_i_m[0:0]),.pre_out_0(pre_out_0[11:1]),.output_iv({output_iv[10:10],output_iv_0[9:7],output_iv[6:5],output_iv_0[4:4],output_iv[3:3],output_iv_0[2:2],output_iv[1:0]}),.output_iv_0_0(output_iv_0[1:1]),.output_iv_0_1(output_iv[2:2]),.output_iv_0_2(output_iv_0[3:3]),.output_iv_0_3(output_iv[4:4]),.output_iv_0_4(output_iv_0[5:5]),.output_iv_0_6(output_iv[7:7]),.output_iv_0_7(output_iv[8:8]),.output_iv_0_8(output_iv[9:9]),.output_iv_0_9(output_iv_0[10:10]),.out_i_vec_sub_0(out_i_vec_sub_0[11:11]),.out_i_vec_mult_0(out_i_vec_mult_0[11:0]),.pre_out_i_m_2(pre_out_i_m_0[0:0]),.out_i_vec_mult_1(out_i_vec_mult_1[11:0]),.pre_out_1(pre_out_1[11:1]),.pre_out_4(pre_out_2[11:11]),.pre_out_i_m_3(pre_out_i_m_1),.out_i_vec_mult_2(out_i_vec_mult_2[11:0]),.pre_out_2({pre_out_3[11:11],pre_out_2[10:1]}),.pre_out_5(pre_out_4[11:11]),.out_i_vec_mult_3(out_i_vec_mult_3[11:0]),.pre_out_i_m({pre_out_i_m[10:1],pre_out_i_m_2}),.pre_out_i_m_0_0(pre_out_i_m_3),.pre_out_i_m_0_1(pre_out_i_m_0[1:1]),.pre_out_i_m_0_6(pre_out_i_m_0[6:6]),.pre_out_i_m_0_4(pre_out_i_m_0[4:4]),.pre_out_i_m_4(pre_out_i_m_4),.pre_out_6(pre_out_5[11:11]),.pre_out_3_9(pre_out_6[11:11]),.pre_out_3_0(pre_out_3[2:2]),.pre_out_3_1(pre_out_3[3:3]),.pre_out_3_3(pre_out_3[5:5]),.pre_out_3_5(pre_out_3[7:7]),.pre_out_3_7(pre_out_3[9:9]),.pre_out_3_8(pre_out_3[10:10]),.pre_out_3_6(pre_out_3[8:8]),.clk(clk),.w_in_a_vec_sub(w_in_a_vec_sub),.N_500(N_500),.un5_output(un5_output),.un5_output_0(un5_output_0),.un5_output_1(un5_output_1),.un5_output_2(un5_output_2),.un5_output_3(un5_output_3),.un5_output_4(un5_output_4),.p_desc739_p_O_FDE(p_desc739_p_O_FDEvec_sub_),.p_desc740_p_O_FDE(p_desc740_p_O_FDEvec_sub_),.p_desc741_p_O_FDE(p_desc741_p_O_FDEvec_sub_),.p_desc742_p_O_FDE(p_desc742_p_O_FDEvec_sub_),.p_desc743_p_O_FDE(p_desc743_p_O_FDEvec_sub_),.p_desc744_p_O_FDE(p_desc744_p_O_FDEvec_sub_),.p_desc745_p_O_FDE(p_desc745_p_O_FDEvec_sub_),.p_desc746_p_O_FDE(p_desc746_p_O_FDEvec_sub_),.p_desc747_p_O_FDE(p_desc747_p_O_FDEvec_sub_),.p_desc748_p_O_FDE(p_desc748_p_O_FDEvec_sub_),.p_desc749_p_O_FDE(p_desc749_p_O_FDEvec_sub_),.p_desc750_p_O_FDE(p_desc750_p_O_FDEvec_sub_),.p_desc751_p_O_FDE(p_desc751_p_O_FDEvec_sub_),.p_desc752_p_O_FDE(p_desc752_p_O_FDEvec_sub_),.p_desc753_p_O_FDE(p_desc753_p_O_FDEvec_sub_),.p_desc754_p_O_FDE(p_desc754_p_O_FDEvec_sub_),.p_desc755_p_O_FDE(p_desc755_p_O_FDEvec_sub_),.p_desc756_p_O_FDE(p_desc756_p_O_FDEvec_sub_),.p_desc757_p_O_FDE(p_desc757_p_O_FDEvec_sub_),.p_desc758_p_O_FDE(p_desc758_p_O_FDEvec_sub_),.p_desc759_p_O_FDE(p_desc759_p_O_FDEvec_sub_),.p_desc760_p_O_FDE(p_desc760_p_O_FDEvec_sub_),.p_desc761_p_O_FDE(p_desc761_p_O_FDEvec_sub_),.p_desc762_p_O_FDE(p_desc762_p_O_FDEvec_sub_),.p_desc763_p_O_FDE(p_desc763_p_O_FDEvec_sub_),.p_desc764_p_O_FDE(p_desc764_p_O_FDEvec_sub_),.p_desc765_p_O_FDE(p_desc765_p_O_FDEvec_sub_),.p_desc766_p_O_FDE(p_desc766_p_O_FDEvec_sub_),.p_desc767_p_O_FDE(p_desc767_p_O_FDEvec_sub_),.p_desc768_p_O_FDE(p_desc768_p_O_FDEvec_sub_),.p_desc769_p_O_FDE(p_desc769_p_O_FDEvec_sub_),.p_desc770_p_O_FDE(p_desc770_p_O_FDEvec_sub_),.p_desc771_p_O_FDE(p_desc771_p_O_FDEvec_sub_),.p_desc772_p_O_FDE(p_desc772_p_O_FDEvec_sub_),.p_desc773_p_O_FDE(p_desc773_p_O_FDEvec_sub_),.p_desc774_p_O_FDE(p_desc774_p_O_FDEvec_sub_),.p_desc775_p_O_FDE(p_desc775_p_O_FDEvec_sub_),.p_desc776_p_O_FDE(p_desc776_p_O_FDEvec_sub_),.p_desc777_p_O_FDE(p_desc777_p_O_FDEvec_sub_),.p_desc778_p_O_FDE(p_desc778_p_O_FDEvec_sub_),.p_desc779_p_O_FDE(p_desc779_p_O_FDEvec_sub_),.p_desc780_p_O_FDE(p_desc780_p_O_FDEvec_sub_),.p_desc781_p_O_FDE(p_desc781_p_O_FDEvec_sub_),.p_desc782_p_O_FDE(p_desc782_p_O_FDEvec_sub_),.p_desc783_p_O_FDE(p_desc783_p_O_FDEvec_sub_),.p_desc784_p_O_FDE(p_desc784_p_O_FDEvec_sub_),.p_desc785_p_O_FDE(p_desc785_p_O_FDEvec_sub_),.p_desc786_p_O_FDE(p_desc786_p_O_FDEvec_sub_),.p_desc787_p_O_FDE(p_desc787_p_O_FDEvec_sub_),.p_desc788_p_O_FDE(p_desc788_p_O_FDEvec_sub_),.p_desc789_p_O_FDE(p_desc789_p_O_FDEvec_sub_),.p_desc790_p_O_FDE(p_desc790_p_O_FDEvec_sub_),.p_desc791_p_O_FDE(p_desc791_p_O_FDEvec_sub_),.p_desc792_p_O_FDE(p_desc792_p_O_FDEvec_sub_),.p_desc793_p_O_FDE(p_desc793_p_O_FDEvec_sub_),.p_desc794_p_O_FDE(p_desc794_p_O_FDEvec_sub_),.p_desc795_p_O_FDE(p_desc795_p_O_FDEvec_sub_),.p_desc796_p_O_FDE(p_desc796_p_O_FDEvec_sub_),.p_desc797_p_O_FDE(p_desc797_p_O_FDEvec_sub_),.p_desc798_p_O_FDE(p_desc798_p_O_FDEvec_sub_),.p_desc799_p_O_FDE(p_desc799_p_O_FDEvec_sub_),.p_desc800_p_O_FDE(p_desc800_p_O_FDEvec_sub_),.p_desc801_p_O_FDE(p_desc801_p_O_FDEvec_sub_),.p_desc802_p_O_FDE(p_desc802_p_O_FDEvec_sub_),.p_desc803_p_O_FDE(p_desc803_p_O_FDEvec_sub_),.p_desc804_p_O_FDE(p_desc804_p_O_FDEvec_sub_),.p_desc805_p_O_FDE(p_desc805_p_O_FDEvec_sub_),.p_desc806_p_O_FDE(p_desc806_p_O_FDEvec_sub_),.p_desc807_p_O_FDE(p_desc807_p_O_FDEvec_sub_),.p_desc808_p_O_FDE(p_desc808_p_O_FDEvec_sub_),.p_desc809_p_O_FDE(p_desc809_p_O_FDEvec_sub_),.p_desc810_p_O_FDE(p_desc810_p_O_FDEvec_sub_),.p_desc811_p_O_FDE(p_desc811_p_O_FDEvec_sub_),.p_desc812_p_O_FDE(p_desc812_p_O_FDEvec_sub_),.p_desc813_p_O_FDE(p_desc813_p_O_FDEvec_sub_),.p_desc814_p_O_FDE(p_desc814_p_O_FDEvec_sub_),.p_desc815_p_O_FDE(p_desc815_p_O_FDEvec_sub_),.p_desc816_p_O_FDE(p_desc816_p_O_FDEvec_sub_),.p_desc817_p_O_FDE(p_desc817_p_O_FDEvec_sub_),.p_desc818_p_O_FDE(p_desc818_p_O_FDEvec_sub_),.p_desc819_p_O_FDE(p_desc819_p_O_FDEvec_sub_),.p_desc820_p_O_FDE(p_desc820_p_O_FDEvec_sub_),.p_desc821_p_O_FDE(p_desc821_p_O_FDEvec_sub_),.p_desc822_p_O_FDE(p_desc822_p_O_FDEvec_sub_),.p_desc823_p_O_FDE(p_desc823_p_O_FDEvec_sub_),.p_desc824_p_O_FDE(p_desc824_p_O_FDEvec_sub_),.p_desc825_p_O_FDE(p_desc825_p_O_FDEvec_sub_),.p_desc826_p_O_FDE(p_desc826_p_O_FDEvec_sub_),.p_desc827_p_O_FDE(p_desc827_p_O_FDEvec_sub_),.p_desc828_p_O_FDE(p_desc828_p_O_FDEvec_sub_),.p_desc829_p_O_FDE(p_desc829_p_O_FDEvec_sub_),.p_desc830_p_O_FDE(p_desc830_p_O_FDEvec_sub_),.p_desc831_p_O_FDE(p_desc831_p_O_FDEvec_sub_),.p_desc832_p_O_FDE(p_desc832_p_O_FDEvec_sub_),.p_desc833_p_O_FDE(p_desc833_p_O_FDEvec_sub_),.p_desc834_p_O_FDE(p_desc834_p_O_FDEvec_sub_));
  mult_with_reg_inj r_mult(.un8_rnd_out(un8_rnd_out[10:0]),.un8_rnd_out_P_19(un8_rnd_out_P[19:19]),.out_inv_sqrt_0(out_inv_sqrt[0:0]),.out_inv_sqrt_1(out_inv_sqrt[1:1]),.out_inv_sqrt_2(out_inv_sqrt[2:2]),.out_inv_sqrt_7(out_inv_sqrt[7:7]),.out_inv_sqrt_8(out_inv_sqrt[8:8]),.out_inv_sqrt_9(out_inv_sqrt[9:9]),.out_inv_sqrt_10(out_inv_sqrt[10:10]),.out_inv_sqrt_11(out_inv_sqrt[11:11]),.out_inner_prod_r(out_inner_prod_r[11:0]),.pre_out_19(pre_out[19:19]),.pre_out_20(pre_out[20:20]),.pre_out_21(pre_out[21:21]),.pre_out_22(pre_out[22:22]),.pre_out_reg(pre_out_reg[23:23]),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i),.N_512_i(N_512_i),.clk(clk),.PATTERNDETECT_32(PATTERNDETECT_32));
  inv_sqrt_inj inv_sqrt_inst(.out_inner_prod_r(out_inner_prod_r[11:0]),.out_inv_sqrt_9(out_inv_sqrt[9:9]),.out_inv_sqrt_10(out_inv_sqrt[10:10]),.out_inv_sqrt_8(out_inv_sqrt[8:8]),.out_inv_sqrt_7(out_inv_sqrt[7:7]),.out_inv_sqrt_2(out_inv_sqrt[2:2]),.out_inv_sqrt_1(out_inv_sqrt[1:1]),.out_inv_sqrt_11(out_inv_sqrt[11:11]),.out_inv_sqrt_0(out_inv_sqrt[0:0]),.done_inv_sqrt(done_inv_sqrt),.clk(clk),.rst(rst),.start_inv_sqrt(start_inv_sqrt),.N_434_i(N_434_i),.N_431_i(N_431_i),.N_428_i(N_428_i),.N_425_i(N_425_i),.p_output_reg_pipe_13_Z_p_O_FDshifterZ0_(p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_),.p_output_reg_pipe_12_Z_p_O_FDshifterZ0_(p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_),.p_output_reg_pipe_Z_p_O_FDshifterZ0_(p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_),.p_desc951_p_O_FDE(p_desc951_p_O_FDEinv_sqrt_),.p_desc952_p_O_FDE(p_desc952_p_O_FDEinv_sqrt_),.p_desc953_p_O_FDE(p_desc953_p_O_FDEinv_sqrt_),.p_desc954_p_O_FDE(p_desc954_p_O_FDEinv_sqrt_),.p_desc955_p_O_FDE(p_desc955_p_O_FDEinv_sqrt_),.p_desc956_p_O_FDE(p_desc956_p_O_FDEinv_sqrt_),.p_desc957_p_O_FDE(p_desc957_p_O_FDEinv_sqrt_),.p_desc958_p_O_FDE(p_desc958_p_O_FDEinv_sqrt_),.p_desc959_p_O_FDE(p_desc959_p_O_FDEinv_sqrt_),.p_desc960_p_O_FDE(p_desc960_p_O_FDEinv_sqrt_),.p_desc961_p_O_FDE(p_desc961_p_O_FDEinv_sqrt_),.p_desc962_p_O_FDE(p_desc962_p_O_FDEinv_sqrt_),.p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_(p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_),.p_output_reg_pipe_Z_p_O_FDRE(p_output_reg_pipe_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_3_Z_p_O_FDRE(p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_6_Z_p_O_FDRE(p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_9_Z_p_O_FDRE(p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_12_Z_p_O_FDRE(p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_15_Z_p_O_FDRE(p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_16_Z_p_O_FDRE(p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_17_Z_p_O_FDRE(p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_18_Z_p_O_FDRE(p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_),.p_output_reg_pipe_21_Z_p_O_FDRE(p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_),.p_done_Z_p_O_FDC(p_done_Z_p_O_FDCinv_sqrt_),.p_desc946_p_O_FDC(p_desc946_p_O_FDCinv_sqrt_),.p_desc947_p_O_FDC(p_desc947_p_O_FDCinv_sqrt_),.p_desc948_p_O_FDC(p_desc948_p_O_FDCinv_sqrt_),.p_desc949_p_O_FDC(p_desc949_p_O_FDCinv_sqrt_),.p_desc950_p_O_FDC(p_desc950_p_O_FDCinv_sqrt_));
  qr_decomp_ctl_mux_inj muxes(.single_in_R_sel(single_in_R_sel),.single_in_R_sel_0(single_in_R_sel_0),.w_col_sel_AQ_int(w_col_sel_AQ_int[1:0]),.col_sel_AQ(col_sel_AQ[1:0]),.wr_en_AQ_sel(wr_en_AQ_sel),.w_col_sel_AQ_mux_i_m3_lut6_2_O6(w_col_sel_AQ_mux_i_m3_lut6_2_O6),.w_col_sel_AQ_mux_i_m3_lut6_2_O5(w_col_sel_AQ_mux_i_m3_lut6_2_O5),.col_sel_AQ2_int(col_sel_AQ2_int[1:0]),.col_sel_AQ2_mux_i_m3_lut6_2_O6(col_sel_AQ2_mux_i_m3_lut6_2_O6),.col_sel_AQ2_mux_i_m3_lut6_2_O5(col_sel_AQ2_mux_i_m3_lut6_2_O5),.state_0(state[3:3]),.state_2(state[5:5]),.state_5(state[8:8]),.wr_en_AQ_sel_0(wr_en_AQ_sel_0),.col_sel_R(col_sel_R[1:0]),.col_sel_R_int(col_sel_R_int[1:0]),.col_sel_R_mux_i_m3_lut6_2_O6(col_sel_R_mux_i_m3_lut6_2_O6),.col_sel_R_mux_i_m3_lut6_2_O5(col_sel_R_mux_i_m3_lut6_2_O5),.in_a_r_reg_0_0(in_a_r_reg_0[0:0]),.in_a_r_reg_0_11(in_a_r_reg_0[11:11]),.out_r_vec_sub_0(out_r_vec_sub_0[11:11]),.in_a_i_reg_1(in_a_i_reg_1[11:11]),.vec_in_AQ_sel(vec_in_AQ_sel[1:0]),.in_a_r_reg_3(in_a_r_reg_3[11:11]),.in_a_i_reg_0(in_a_i_reg_0[11:11]),.in_a_i_reg_3(in_a_i_reg_3[11:11]),.in_a_r_reg_1(in_a_r_reg_1[11:11]),.pre_out_4(pre_out_0[11:11]),.pre_out_0({pre_out_2[11:11],pre_out_1[10:9],pre_out_0[8:8],pre_out_1[7:7],pre_out_0[6:6],pre_out_1[5:5],pre_out_0[4:4],pre_out_1[3:2],pre_out[1:1]}),.in_a_r_reg_2(in_a_r_reg_2[11:11]),.pre_out_5(pre_out_1[11:11]),.pre_out_1({pre_out_3[11:11],pre_out[10:9],pre_out_3[8:8],pre_out[7:2],pre_out_0[1:1]}),.in_a_i_reg_2(in_a_i_reg_2[11:11]),.pre_out_6(pre_out_4[11:11]),.pre_out_3_9(pre_out_5[11:11]),.pre_out_3_1(pre_out_3[3:3]),.pre_out_3_7(pre_out_3[9:9]),.pre_out_3_3(pre_out_3[5:5]),.pre_out_3_8(pre_out_3[10:10]),.pre_out_3_5(pre_out_3[7:7]),.pre_out_3_6(pre_out_2[8:8]),.pre_out_3_0(pre_out_3[2:2]),.pre_out_2({pre_out_6[11:11],pre_out_0[10:9],pre_out[8:8],pre_out_0[7:7],pre_out_2[6:6],pre_out_0[5:5],pre_out_2[4:4],pre_out_0[3:2],pre_out_2[1:1]}),.out_inner_prod_i(out_inner_prod_i[11:0]),.pre_out_10(pre_out[11:11]),.pre_out_9(pre_out_2[10:10]),.pre_out_0_d0(pre_out_1[1:1]),.pre_out_1_d0(pre_out_2[2:2]),.pre_out_3_d0(pre_out_1[4:4]),.pre_out_6_d0(pre_out_2[7:7]),.pre_out_7(pre_out_1[8:8]),.pre_out_8(pre_out_2[9:9]),.pre_out_5_d0(pre_out_1[6:6]),.pre_out_4_d0(pre_out_2[5:5]),.pre_out_2_d0(pre_out_2[3:3]),.pre_out_18(pre_out[19:19]),.pre_out_19(pre_out[20:20]),.pre_out_20(pre_out[21:21]),.pre_out_21(pre_out[22:22]),.pre_out_reg(pre_out_reg[23:23]),.out_r_vec_mult_2(out_r_vec_mult_2[11:0]),.vec_in_r_AQ_mux_2(vec_in_r_AQ_mux_2[11:0]),.out_r_vec_mult_1(out_r_vec_mult_1[11:0]),.vec_in_r_AQ_mux_1(vec_in_r_AQ_mux_1[11:0]),.pre_out_i_m({pre_out_i_m[10:2],pre_out_i_m_0[1:1],pre_out_i_m_3}),.out_i_vec_mult_3(out_i_vec_mult_3[11:0]),.pre_out_i_m_1(pre_out_i_m_4),.vec_in_i_AQ_mux_3(vec_in_i_AQ_mux_3[11:0]),.output_iv({output_iv[10:10],output_iv_0[9:9],output_iv[8:8],output_iv_0[7:7],output_iv[6:5],output_iv_0[4:3],output_iv[2:2],output_iv_0[1:1],output_iv[0:0]}),.out_i_vec_mult_0(out_i_vec_mult_0[11:0]),.vec_in_i_AQ_mux_0_11(vec_in_i_AQ_mux_0[11:11]),.vec_in_i_AQ_mux_0_1(vec_in_i_AQ_mux_0[1:1]),.vec_in_i_AQ_mux_0_5(vec_in_i_AQ_mux_0[5:5]),.vec_in_i_AQ_mux_0_0(vec_in_i_AQ_mux_0[0:0]),.vec_in_i_AQ_mux_0_8(vec_in_i_AQ_mux_0[8:8]),.vec_in_i_AQ_mux_0_10(vec_in_i_AQ_mux_0[10:10]),.vec_in_i_AQ_mux_0_7(vec_in_i_AQ_mux_0[7:7]),.vec_in_i_AQ_mux_0_6(vec_in_i_AQ_mux_0[6:6]),.vec_in_i_AQ_mux_0_9(vec_in_i_AQ_mux_0[9:9]),.vec_in_i_AQ_mux_0_4(vec_in_i_AQ_mux_0[4:4]),.out_r_vec_mult_0(out_r_vec_mult_0[11:0]),.output_iv_0_2(output_iv[3:3]),.output_iv_0_4(output_iv_0[5:5]),.output_iv_0_1(output_iv_0[2:2]),.output_iv_0_0(output_iv[1:1]),.output_iv_0_9(output_iv_0[10:10]),.output_iv_0_6(output_iv[7:7]),.output_iv_0_8(output_iv[9:9]),.output_iv_0_3(output_iv[4:4]),.output_iv_0_7(output_iv_0[8:8]),.vec_in_r_AQ_mux_0_10(vec_in_r_AQ_mux_0[11:11]),.vec_in_r_AQ_mux_0_2(vec_in_r_AQ_mux_0[3:3]),.vec_in_r_AQ_mux_0_4(vec_in_r_AQ_mux_0[5:5]),.vec_in_r_AQ_mux_0_3(vec_in_r_AQ_mux_0[4:4]),.vec_in_r_AQ_mux_0_6(vec_in_r_AQ_mux_0[7:7]),.vec_in_r_AQ_mux_0_1(vec_in_r_AQ_mux_0[2:2]),.vec_in_r_AQ_mux_0_9(vec_in_r_AQ_mux_0[10:10]),.vec_in_r_AQ_mux_0_8(vec_in_r_AQ_mux_0[9:9]),.vec_in_r_AQ_mux_0_0(vec_in_r_AQ_mux_0[1:1]),.vec_in_r_AQ_mux_0_7(vec_in_r_AQ_mux_0[8:8]),.pre_out_i_m_0_0(pre_out_i_m_2),.pre_out_i_m_0_6(pre_out_i_m_0[6:6]),.pre_out_i_m_0_4(pre_out_i_m_0[4:4]),.pre_out_i_m_0_1(pre_out_i_m[1:1]),.in_A_r(in_A_r[47:0]),.out_r_vec_mult_3(out_r_vec_mult_3[11:0]),.pre_out_i_m_2(pre_out_i_m[0:0]),.vec_in_r_AQ_mux_3(vec_in_r_AQ_mux_3[11:0]),.out_i_vec_mult_2(out_i_vec_mult_2[11:0]),.pre_out_i_m_3(pre_out_i_m_1),.vec_in_i_AQ_mux_2(vec_in_i_AQ_mux_2[11:0]),.in_A_i(in_A_i[47:0]),.out_i_vec_mult_1(out_i_vec_mult_1[11:0]),.pre_out_i_m_4(pre_out_i_m_0[0:0]),.vec_in_i_AQ_mux_1(vec_in_i_AQ_mux_1[11:0]),.un8_rnd_out_P(un8_rnd_out_P[19:19]),.single_in_r_R_mux(single_in_r_R_mux[11:11]),.out_inner_prod_r(out_inner_prod_r[11:0]),.un8_rnd_out(un8_rnd_out[10:0]),.N_390_i(N_390_i),.N_393_i(N_393_i),.done_inv_sqrt(done_inv_sqrt),.N_391_i(N_391_i),.N_394_i(N_394_i),.N_396_i(N_396_i),.N_395_i(N_395_i),.N_397_i(N_397_i),.N_398_i(N_398_i),.N_400_i(N_400_i),.N_399_i(N_399_i),.N_401_i(N_401_i),.wr_en_AQ_int(wr_en_AQ_int),.wr_A_QR(wr_A_QR),.start_QR(start_QR),.wr_en_AQ_mux_i_m3_lut6_2_O6(wr_en_AQ_mux_i_m3_lut6_2_O6),.N_501(N_501),.N_392_i(N_392_i),.PATTERNDETECT_32(PATTERNDETECT_32),.N_500(N_500),.N_508(N_508),.N_507(N_507),.N_506(N_506),.N_505(N_505),.un5_output(un5_output_0),.un5_output_0(un5_output),.un5_output_1(un5_output_4),.un5_output_2(un5_output_1),.un5_output_3(un5_output_3),.un5_output_4(un5_output_2),.N_389_i(N_389_i),.N_388_i(N_388_i),.N_387_i(N_387_i),.N_386_i(N_386_i),.N_385_i(N_385_i),.N_384_i(N_384_i),.N_383_i(N_383_i),.N_34_i(N_34_i),.N_32_i(N_32_i),.N_30_i(N_30_i),.N_28_i(N_28_i));
  qr_decomp_ctl_inj the_ctl(.col_sel_AQ_int(col_sel_AQ_int[1:0]),.col_sel_AQ2_int(col_sel_AQ2_int[1:0]),.row_sel_AQ(row_sel_AQ[1:0]),.state_5(state[5:5]),.state_8(state[8:8]),.state_3(state[3:3]),.in_b_inner_prod_sel(in_b_inner_prod_sel),.w_col_sel_AQ_int(w_col_sel_AQ_int[1:0]),.col_sel_R_int(col_sel_R_int[1:0]),.row_sel_R(row_sel_R[1:0]),.in_a_inner_prod_sel(in_a_inner_prod_sel),.vec_in_AQ_sel(vec_in_AQ_sel[1:0]),.single_in_R_sel(single_in_R_sel),.single_in_R_sel_0(single_in_R_sel_0),.wr_en_AQ_sel(wr_en_AQ_sel),.wr_en_AQ_sel_0(wr_en_AQ_sel_0),.in_b_vec_mult_sel(in_b_vec_mult_sel),.red_mat_reg(red_mat_reg),.rst(rst),.done_inv_sqrt(done_inv_sqrt),.N_512_i(N_512_i),.done_inner_prod(done_inner_prod),.start_inv_sqrt(start_inv_sqrt),.clk(clk),.start_inner_prod(start_inner_prod),.wr_en_AQ_int(wr_en_AQ_int),.wr_en_R(wr_en_R),.w_in_a_vec_sub(w_in_a_vec_sub),.done_QR(done_QR),.start_QR(start_QR),.red_mat_reg_0(red_mat_reg_0),.p_desc1255_p_O_FDC(p_desc1255_p_O_FDCqr_decomp_ctl_),.p_desc1256_p_O_FDC(p_desc1256_p_O_FDCqr_decomp_ctl_),.p_desc1257_p_O_FDC(p_desc1257_p_O_FDCqr_decomp_ctl_),.p_desc1258_p_O_FDC(p_desc1258_p_O_FDCqr_decomp_ctl_),.p_start_inner_prod_Z_p_O_FDC(p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_),.p_wr_en_AQ_int_Z_p_O_FDC(p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_),.p_wr_en_R_Z_p_O_FDC(p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_),.p_w_in_a_vec_sub_Z_p_O_FDC(p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_),.p_start_inv_sqrt_Z_p_O_FDC(p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_),.p_desc1274_p_O_FDC(p_desc1274_p_O_FDCqr_decomp_ctl_),.p_pre_red_mat_reg_Z_p_O_FDC(p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_),.p_done_Z_p_O_FDC(p_done_Z_p_O_FDCqr_decomp_ctl_),.p_desc1275_p_O_FDC(p_desc1275_p_O_FDCqr_decomp_ctl_),.p_desc1276_p_O_FDC(p_desc1276_p_O_FDCqr_decomp_ctl_),.p_desc1277_p_O_FDC(p_desc1277_p_O_FDCqr_decomp_ctl_),.p_desc1278_p_O_FDC(p_desc1278_p_O_FDCqr_decomp_ctl_),.p_desc1279_p_O_FDC(p_desc1279_p_O_FDCqr_decomp_ctl_),.p_desc1281_p_O_FDC(p_desc1281_p_O_FDCqr_decomp_ctl_),.p_desc1282_p_O_FDC(p_desc1282_p_O_FDCqr_decomp_ctl_),.p_desc1283_p_O_FDC(p_desc1283_p_O_FDCqr_decomp_ctl_),.p_desc1284_p_O_FDC(p_desc1284_p_O_FDCqr_decomp_ctl_),.p_desc1285_p_O_FDC(p_desc1285_p_O_FDCqr_decomp_ctl_),.p_desc1286_p_O_FDC(p_desc1286_p_O_FDCqr_decomp_ctl_),.p_desc1287_p_O_FDC(p_desc1287_p_O_FDCqr_decomp_ctl_),.p_desc1288_p_O_FDC(p_desc1288_p_O_FDCqr_decomp_ctl_),.p_desc1265_p_O_FDP(p_desc1265_p_O_FDPqr_decomp_ctl_),.p_desc1268_p_O_FDP(p_desc1268_p_O_FDPqr_decomp_ctl_),.p_desc1280_p_O_FDP(p_desc1280_p_O_FDPqr_decomp_ctl_),.p_desc1263_p_O_FDCE(p_desc1263_p_O_FDCEqr_decomp_ctl_),.p_desc1264_p_O_FDCE(p_desc1264_p_O_FDCEqr_decomp_ctl_),.p_desc1266_p_O_FDCE(p_desc1266_p_O_FDCEqr_decomp_ctl_),.p_desc1267_p_O_FDCE(p_desc1267_p_O_FDCEqr_decomp_ctl_),.p_desc1269_p_O_FDCE(p_desc1269_p_O_FDCEqr_decomp_ctl_),.p_desc1270_p_O_FDCE(p_desc1270_p_O_FDCEqr_decomp_ctl_),.p_desc1271_p_O_FDCE(p_desc1271_p_O_FDCEqr_decomp_ctl_),.p_desc1272_p_O_FDCE(p_desc1272_p_O_FDCEqr_decomp_ctl_),.p_desc1273_p_O_FDCE(p_desc1273_p_O_FDCEqr_decomp_ctl_));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module qr_decomp_ctl_inj (col_sel_AQ_int,col_sel_AQ2_int,row_sel_AQ,state_5,state_8,state_3,in_b_inner_prod_sel,w_col_sel_AQ_int,col_sel_R_int,row_sel_R,in_a_inner_prod_sel,vec_in_AQ_sel,single_in_R_sel,single_in_R_sel_0,wr_en_AQ_sel,wr_en_AQ_sel_0,in_b_vec_mult_sel,red_mat_reg,rst,done_inv_sqrt,N_512_i,done_inner_prod,start_inv_sqrt,clk,start_inner_prod,wr_en_AQ_int,wr_en_R,w_in_a_vec_sub,done_QR,start_QR,red_mat_reg_0,p_desc1255_p_O_FDC,p_desc1256_p_O_FDC,p_desc1257_p_O_FDC,p_desc1258_p_O_FDC,p_start_inner_prod_Z_p_O_FDC,p_wr_en_AQ_int_Z_p_O_FDC,p_wr_en_R_Z_p_O_FDC,p_w_in_a_vec_sub_Z_p_O_FDC,p_start_inv_sqrt_Z_p_O_FDC,p_desc1274_p_O_FDC,p_pre_red_mat_reg_Z_p_O_FDC,p_done_Z_p_O_FDC,p_desc1275_p_O_FDC,p_desc1276_p_O_FDC,p_desc1277_p_O_FDC,p_desc1278_p_O_FDC,p_desc1279_p_O_FDC,p_desc1281_p_O_FDC,p_desc1282_p_O_FDC,p_desc1283_p_O_FDC,p_desc1284_p_O_FDC,p_desc1285_p_O_FDC,p_desc1286_p_O_FDC,p_desc1287_p_O_FDC,p_desc1288_p_O_FDC,p_desc1265_p_O_FDP,p_desc1268_p_O_FDP,p_desc1280_p_O_FDP,p_desc1263_p_O_FDCE,p_desc1264_p_O_FDCE,p_desc1266_p_O_FDCE,p_desc1267_p_O_FDCE,p_desc1269_p_O_FDCE,p_desc1270_p_O_FDCE,p_desc1271_p_O_FDCE,p_desc1272_p_O_FDCE,p_desc1273_p_O_FDCE);
output [1:0] col_sel_AQ_int ;
output [1:0] col_sel_AQ2_int ;
output [1:0] row_sel_AQ ;
output state_5 ;
output state_8 ;
output state_3 ;
output in_b_inner_prod_sel ;
output [1:0] w_col_sel_AQ_int ;
output [1:0] col_sel_R_int ;
output [1:0] row_sel_R ;
output in_a_inner_prod_sel ;
output [1:0] vec_in_AQ_sel ;
output single_in_R_sel ;
input single_in_R_sel_0 ;
output wr_en_AQ_sel ;
input wr_en_AQ_sel_0 ;
output in_b_vec_mult_sel ;
output red_mat_reg ;
input rst ;
input done_inv_sqrt ;
output N_512_i ;
input done_inner_prod ;
output start_inv_sqrt ;
input clk ;
output start_inner_prod ;
output wr_en_AQ_int ;
output wr_en_R ;
output w_in_a_vec_sub ;
output done_QR ;
input start_QR ;
input red_mat_reg_0 ;
wire state_5 ;
wire state_8 ;
wire state_3 ;
wire red_mat_reg ;
wire rst ;
wire done_inv_sqrt ;
wire N_512_i ;
wire done_inner_prod ;
wire start_inv_sqrt ;
wire clk ;
wire start_inner_prod ;
wire wr_en_AQ_int ;
wire wr_en_R ;
wire w_in_a_vec_sub ;
wire done_QR ;
wire start_QR ;
wire red_mat_reg_0 ;
wire [7:0] state ;
wire [2:0] mult_counter ;
wire [5:5] state_ns_2_tz ;
wire [7:1] state_ns ;
wire in_b_inner_prod_sel_0 ;
wire [1:0] w_col_sel_AQ_int_4_i_m2_i_m3 ;
wire [1:0] col_sel_R_int_4_i_m2_i_m3 ;
wire in_a_inner_prod_sel_0 ;
wire [1:1] j_RNO ;
wire VCC ;
wire N_676 ;
wire N_210_i ;
wire N_526 ;
wire row_sel_R_0_sqmuxa ;
wire row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_O5 ;
wire N_662 ;
wire N_201_2 ;
wire N_706 ;
wire N_686 ;
wire N_495 ;
wire N_503 ;
wire N_652 ;
wire un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_O6 ;
wire un1_state_10_0_o6_0_o2_lut6_2_O6 ;
wire N_653 ;
wire start_inv_sqrt_0 ;
wire un1_state_23_0_0_o2_lut6_2_O6 ;
wire N_513_i ;
wire N_218_i ;
wire un1_state_33_0_0 ;
wire N_220_i ;
wire start_inner_prod_0 ;
wire wr_en_AQ_int_0 ;
wire un1_state_29_0_0 ;
wire N_514_i ;
wire wr_en_R_0 ;
wire w_in_a_vec_sub_0 ;
wire pre_red_mat_reg ;
wire done ;
wire N_214_i ;
wire N_216_i ;
wire N_231_i ;
wire N_201_i ;
wire N_196_3 ;
wire N_106_1 ;
wire N_527 ;
wire N_106_2 ;
wire N_123 ;
wire N_122 ;
wire N_121 ;
wire N_120 ;
wire N_119 ;
wire N_118 ;
wire N_117 ;
wire N_116 ;
wire N_115 ;
wire GND ;
input p_desc1255_p_O_FDC ;
input p_desc1256_p_O_FDC ;
input p_desc1257_p_O_FDC ;
input p_desc1258_p_O_FDC ;
input p_start_inner_prod_Z_p_O_FDC ;
input p_wr_en_AQ_int_Z_p_O_FDC ;
input p_wr_en_R_Z_p_O_FDC ;
input p_w_in_a_vec_sub_Z_p_O_FDC ;
input p_start_inv_sqrt_Z_p_O_FDC ;
input p_desc1274_p_O_FDC ;
input p_pre_red_mat_reg_Z_p_O_FDC ;
input p_done_Z_p_O_FDC ;
input p_desc1275_p_O_FDC ;
input p_desc1276_p_O_FDC ;
input p_desc1277_p_O_FDC ;
input p_desc1278_p_O_FDC ;
input p_desc1279_p_O_FDC ;
input p_desc1281_p_O_FDC ;
input p_desc1282_p_O_FDC ;
input p_desc1283_p_O_FDC ;
input p_desc1284_p_O_FDC ;
input p_desc1285_p_O_FDC ;
input p_desc1286_p_O_FDC ;
input p_desc1287_p_O_FDC ;
input p_desc1288_p_O_FDC ;
input p_desc1265_p_O_FDP ;
input p_desc1268_p_O_FDP ;
input p_desc1280_p_O_FDP ;
input p_desc1263_p_O_FDCE ;
input p_desc1264_p_O_FDCE ;
input p_desc1266_p_O_FDCE ;
input p_desc1267_p_O_FDCE ;
input p_desc1269_p_O_FDCE ;
input p_desc1270_p_O_FDCE ;
input p_desc1271_p_O_FDCE ;
input p_desc1272_p_O_FDCE ;
input p_desc1273_p_O_FDCE ;
// instances
  p_O_FDC desc1255(.Q(w_col_sel_AQ_int[1:1]),.D(w_col_sel_AQ_int_4_i_m2_i_m3[1:1]),.C(clk),.CLR(rst),.E(p_desc1255_p_O_FDC));
  p_O_FDC desc1256(.Q(w_col_sel_AQ_int[0:0]),.D(w_col_sel_AQ_int_4_i_m2_i_m3[0:0]),.C(clk),.CLR(rst),.E(p_desc1256_p_O_FDC));
  p_O_FDC desc1257(.Q(col_sel_R_int[1:1]),.D(col_sel_R_int_4_i_m2_i_m3[1:1]),.C(clk),.CLR(rst),.E(p_desc1257_p_O_FDC));
  p_O_FDC desc1258(.Q(col_sel_R_int[0:0]),.D(col_sel_R_int_4_i_m2_i_m3[0:0]),.C(clk),.CLR(rst),.E(p_desc1258_p_O_FDC));
  LUT5 desc1259(.I0(col_sel_AQ2_int[0:0]),.I1(state[7:7]),.I2(col_sel_AQ_int[0:0]),.I3(w_col_sel_AQ_int[0:0]),.I4(un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_O6),.O(w_col_sel_AQ_int_4_i_m2_i_m3[0:0]));
defparam desc1259.INIT=32'hE2E2FF00;
  LUT5 desc1260(.I0(col_sel_AQ2_int[1:1]),.I1(state[7:7]),.I2(col_sel_AQ_int[1:1]),.I3(w_col_sel_AQ_int[1:1]),.I4(un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_O6),.O(w_col_sel_AQ_int_4_i_m2_i_m3[1:1]));
defparam desc1260.INIT=32'hE2E2FF00;
  LUT5 desc1261(.I0(col_sel_AQ2_int[0:0]),.I1(state_5),.I2(col_sel_AQ_int[0:0]),.I3(col_sel_R_int[0:0]),.I4(un1_state_23_0_0_o2_lut6_2_O6),.O(col_sel_R_int_4_i_m2_i_m3[0:0]));
defparam desc1261.INIT=32'hE2E2FF00;
  LUT5 desc1262(.I0(col_sel_AQ2_int[1:1]),.I1(state_5),.I2(col_sel_AQ_int[1:1]),.I3(col_sel_R_int[1:1]),.I4(un1_state_23_0_0_o2_lut6_2_O6),.O(col_sel_R_int_4_i_m2_i_m3[1:1]));
defparam desc1262.INIT=32'hE2E2FF00;
  p_O_FDCE desc1263(.Q(row_sel_R[0:0]),.D(col_sel_AQ_int[0:0]),.C(clk),.CLR(rst),.CE(row_sel_R_0_sqmuxa),.E(p_desc1263_p_O_FDCE));
  p_O_FDCE desc1264(.Q(row_sel_R[1:1]),.D(col_sel_AQ_int[1:1]),.C(clk),.CLR(rst),.CE(row_sel_R_0_sqmuxa),.E(p_desc1264_p_O_FDCE));
  p_O_FDP desc1265(.Q(in_b_inner_prod_sel),.D(in_b_inner_prod_sel_0),.C(clk),.PRE(rst),.E(p_desc1265_p_O_FDP));
  p_O_FDCE desc1266(.Q(row_sel_AQ[0:0]),.D(N_218_i),.C(clk),.CLR(rst),.CE(un1_state_33_0_0),.E(p_desc1266_p_O_FDCE));
  p_O_FDCE desc1267(.Q(row_sel_AQ[1:1]),.D(N_220_i),.C(clk),.CLR(rst),.CE(un1_state_33_0_0),.E(p_desc1267_p_O_FDCE));
  p_O_FDC start_inner_prod_Z(.Q(start_inner_prod),.D(start_inner_prod_0),.C(clk),.CLR(rst),.E(p_start_inner_prod_Z_p_O_FDC));
  p_O_FDP desc1268(.Q(in_a_inner_prod_sel),.D(in_a_inner_prod_sel_0),.C(clk),.PRE(rst),.E(p_desc1268_p_O_FDP));
  p_O_FDC wr_en_AQ_int_Z(.Q(wr_en_AQ_int),.D(wr_en_AQ_int_0),.C(clk),.CLR(rst),.E(p_wr_en_AQ_int_Z_p_O_FDC));
  p_O_FDCE desc1269(.Q(mult_counter[0:0]),.D(un1_state_23_0_0_o2_lut6_2_O6),.C(clk),.CLR(rst),.CE(un1_state_29_0_0),.E(p_desc1269_p_O_FDCE));
  p_O_FDCE desc1270(.Q(mult_counter[1:1]),.D(N_513_i),.C(clk),.CLR(rst),.CE(un1_state_29_0_0),.E(p_desc1270_p_O_FDCE));
  p_O_FDCE desc1271(.Q(mult_counter[2:2]),.D(N_514_i),.C(clk),.CLR(rst),.CE(un1_state_29_0_0),.E(p_desc1271_p_O_FDCE));
  p_O_FDC wr_en_R_Z(.Q(wr_en_R),.D(wr_en_R_0),.C(clk),.CLR(rst),.E(p_wr_en_R_Z_p_O_FDC));
  p_O_FDCE desc1272(.Q(vec_in_AQ_sel[0:0]),.D(state_5),.C(clk),.CLR(rst),.CE(row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_O5),.E(p_desc1272_p_O_FDCE));
  p_O_FDCE desc1273(.Q(vec_in_AQ_sel[1:1]),.D(state[2:2]),.C(clk),.CLR(rst),.CE(row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_O5),.E(p_desc1273_p_O_FDCE));
  p_O_FDC w_in_a_vec_sub_Z(.Q(w_in_a_vec_sub),.D(w_in_a_vec_sub_0),.C(clk),.CLR(rst),.E(p_w_in_a_vec_sub_Z_p_O_FDC));
  p_O_FDC start_inv_sqrt_Z(.Q(start_inv_sqrt),.D(start_inv_sqrt_0),.C(clk),.CLR(rst),.E(p_start_inv_sqrt_Z_p_O_FDC));
  p_O_FDC desc1274(.Q(single_in_R_sel),.D(single_in_R_sel_0),.C(clk),.CLR(rst),.E(p_desc1274_p_O_FDC));
  p_O_FDC pre_red_mat_reg_Z(.Q(red_mat_reg),.D(pre_red_mat_reg),.C(clk),.CLR(rst),.E(p_pre_red_mat_reg_Z_p_O_FDC));
  p_O_FDC done_Z(.Q(done_QR),.D(done),.C(clk),.CLR(rst),.E(p_done_Z_p_O_FDC));
  p_O_FDC desc1275(.Q(wr_en_AQ_sel),.D(wr_en_AQ_sel_0),.C(clk),.CLR(rst),.E(p_desc1275_p_O_FDC));
  p_O_FDC desc1276(.Q(col_sel_AQ_int[0:0]),.D(N_214_i),.C(clk),.CLR(rst),.E(p_desc1276_p_O_FDC));
  p_O_FDC desc1277(.Q(col_sel_AQ_int[1:1]),.D(N_216_i),.C(clk),.CLR(rst),.E(p_desc1277_p_O_FDC));
  p_O_FDC desc1278(.Q(col_sel_AQ2_int[0:0]),.D(N_231_i),.C(clk),.CLR(rst),.E(p_desc1278_p_O_FDC));
  p_O_FDC desc1279(.Q(col_sel_AQ2_int[1:1]),.D(j_RNO[1:1]),.C(clk),.CLR(rst),.E(p_desc1279_p_O_FDC));
  p_O_FDP desc1280(.Q(state_8),.D(N_201_i),.C(clk),.PRE(rst),.E(p_desc1280_p_O_FDP));
  p_O_FDC desc1281(.Q(state[7:7]),.D(state_ns[1:1]),.C(clk),.CLR(rst),.E(p_desc1281_p_O_FDC));
  p_O_FDC desc1282(.Q(state[6:6]),.D(state_ns[2:2]),.C(clk),.CLR(rst),.E(p_desc1282_p_O_FDC));
  p_O_FDC desc1283(.Q(state_5),.D(state_ns[3:3]),.C(clk),.CLR(rst),.E(p_desc1283_p_O_FDC));
  p_O_FDC desc1284(.Q(state[4:4]),.D(state_ns[4:4]),.C(clk),.CLR(rst),.E(p_desc1284_p_O_FDC));
  p_O_FDC desc1285(.Q(state_3),.D(state_ns[5:5]),.C(clk),.CLR(rst),.E(p_desc1285_p_O_FDC));
  p_O_FDC desc1286(.Q(state[2:2]),.D(state_ns[6:6]),.C(clk),.CLR(rst),.E(p_desc1286_p_O_FDC));
  p_O_FDC desc1287(.Q(state[1:1]),.D(state_ns[7:7]),.C(clk),.CLR(rst),.E(p_desc1287_p_O_FDC));
  p_O_FDC desc1288(.Q(state[0:0]),.D(N_210_i),.C(clk),.CLR(rst),.E(p_desc1288_p_O_FDC));
  FDPE desc1289(.Q(in_b_vec_mult_sel),.D(row_sel_R_0_sqmuxa),.C(clk),.PRE(rst),.CE(un1_state_23_0_0_o2_lut6_2_O6));
  LUT6 un1_state_29_0_0_cZ(.I0(done_inner_prod),.I1(state[1:1]),.I2(state[2:2]),.I3(state[4:4]),.I4(state_5),.I5(done_inv_sqrt),.O(un1_state_29_0_0));
defparam un1_state_29_0_0_cZ.INIT=64'hFFFFFFECFFECFFEC;
  LUT5_L desc1290(.I0(mult_counter[1:1]),.I1(done_inner_prod),.I2(state[2:2]),.I3(state_5),.I4(done_inv_sqrt),.LO(N_514_i));
defparam desc1290.INIT=32'h002A2A2A;
  LUT6_L desc1291(.I0(state_3),.I1(state[1:1]),.I2(mult_counter[2:2]),.I3(state_ns_2_tz[5:5]),.I4(N_526),.I5(N_676),.LO(state_ns[5:5]));
defparam desc1291.INIT=64'hFFFFFFFFEAAAC000;
  LUT6_L desc1292(.I0(start_QR),.I1(state[1:1]),.I2(mult_counter[2:2]),.I3(state_8),.I4(row_sel_AQ[0:0]),.I5(N_676),.LO(N_218_i));
defparam desc1292.INIT=64'h000000000000153F;
  LUT6_L desc1293(.I0(state_3),.I1(state[7:7]),.I2(state_8),.I3(in_a_inner_prod_sel),.I4(N_676),.I5(N_652),.LO(in_a_inner_prod_sel_0));
defparam desc1293.INIT=64'hFEFEFEFEFEFEFFEE;
  LUT6 un1_state_33_0_0_cZ(.I0(state_3),.I1(start_QR),.I2(state[7:7]),.I3(state_8),.I4(N_706),.I5(N_676),.O(un1_state_33_0_0));
defparam un1_state_33_0_0_cZ.INIT=64'hFFFFFFFFFFFFFEFA;
  LUT6_L un1_state_28_i_0_3(.I0(state[7:7]),.I1(done_inner_prod),.I2(state[2:2]),.I3(state_5),.I4(state_8),.I5(N_662),.LO(N_196_3));
defparam un1_state_28_i_0_3.INIT=64'hFFFFFFFFFFFFFFBA;
  LUT6_L desc1294(.I0(state[6:6]),.I1(state[7:7]),.I2(done_inner_prod),.I3(red_mat_reg),.I4(row_sel_AQ[1:1]),.I5(row_sel_AQ[0:0]),.LO(state_ns[2:2]));
defparam desc1294.INIT=64'hCECECE0A0A0A0A0A;
  LUT6_L desc1295(.I0(state_3),.I1(done_inner_prod),.I2(state[2:2]),.I3(red_mat_reg),.I4(row_sel_AQ[1:1]),.I5(row_sel_AQ[0:0]),.LO(state_ns[6:6]));
defparam desc1295.INIT=64'hBABABA3030303030;
  LUT6 desc1296(.I0(col_sel_AQ2_int[0:0]),.I1(state[1:1]),.I2(state[4:4]),.I3(mult_counter[2:2]),.I4(col_sel_AQ_int[1:1]),.I5(col_sel_AQ_int[0:0]),.O(N_106_1));
defparam desc1296.INIT=64'h00008800F8000000;
  LUT4_L w_in_a_vec_sub_e(.I0(done_inner_prod),.I1(state[1:1]),.I2(state[2:2]),.I3(w_in_a_vec_sub),.LO(w_in_a_vec_sub_0));
defparam w_in_a_vec_sub_e.INIT=16'hB3A0;
  LUT6_L desc1297(.I0(col_sel_AQ2_int[1:1]),.I1(red_mat_reg),.I2(mult_counter[2:2]),.I3(state_8),.I4(col_sel_AQ_int[0:0]),.I5(N_495),.LO(N_214_i));
defparam desc1297.INIT=64'h00FF0000001F00E0;
  LUT4_L desc1298(.I0(state[6:6]),.I1(done_inner_prod),.I2(state_5),.I3(done_inv_sqrt),.LO(state_ns[3:3]));
defparam desc1298.INIT=16'h88F8;
  LUT4_L pre_red_mat_reg_e(.I0(red_mat_reg_0),.I1(start_QR),.I2(red_mat_reg),.I3(state_8),.LO(pre_red_mat_reg));
defparam pre_red_mat_reg_e.INIT=16'hB8F0;
  LUT3_L done_e(.I0(done_QR),.I1(state[0:0]),.I2(state_8),.LO(done));
defparam done_e.INIT=8'hCE;
  LUT6 un1_state_1_sqmuxa_3_0_o2_0(.I0(col_sel_AQ2_int[1:1]),.I1(red_mat_reg),.I2(mult_counter[2:2]),.I3(state_8),.I4(col_sel_AQ_int[1:1]),.I5(N_495),.O(N_652));
defparam un1_state_1_sqmuxa_3_0_o2_0.INIT=64'hFF00FF00FFE0FFC0;
  LUT6 desc1299(.I0(col_sel_AQ2_int[1:1]),.I1(state[4:4]),.I2(red_mat_reg),.I3(col_sel_AQ_int[1:1]),.I4(col_sel_AQ_int[0:0]),.I5(N_495),.O(N_527));
defparam desc1299.INIT=64'h000C0000050D0505;
  LUT5_L desc1300(.I0(start_QR),.I1(state[7:7]),.I2(state_8),.I3(N_526),.I4(N_503),.LO(state_ns[1:1]));
defparam desc1300.INIT=32'hECA0FFFF;
  LUT6_L desc1301(.I0(state[0:0]),.I1(state[6:6]),.I2(start_QR),.I3(state[2:2]),.I4(state_5),.I5(N_201_2),.LO(N_201_i));
defparam desc1301.INIT=64'h0000000000000023;
  LUT6_L wr_en_AQ_int_e(.I0(wr_en_AQ_int),.I1(state[6:6]),.I2(state[2:2]),.I3(mult_counter[2:2]),.I4(un1_state_10_0_o6_0_o2_lut6_2_O6),.I5(N_653),.LO(wr_en_AQ_int_0));
defparam wr_en_AQ_int_e.INIT=64'hAAAAAAAAABAAA8A8;
  LUT5_L wr_en_R_e(.I0(state[6:6]),.I1(wr_en_R),.I2(state[2:2]),.I3(state[4:4]),.I4(N_196_3),.LO(wr_en_R_0));
defparam wr_en_R_e.INIT=32'hCCCCDDD8;
  LUT6_L desc1302(.I0(col_sel_AQ2_int[1:1]),.I1(state[1:1]),.I2(mult_counter[2:2]),.I3(state_8),.I4(col_sel_AQ_int[0:0]),.I5(N_527),.LO(N_106_2));
defparam desc1302.INIT=64'hF0FAF0FA002A000A;
  LUT4_L desc1303(.I0(state_8),.I1(col_sel_AQ_int[1:1]),.I2(col_sel_AQ_int[0:0]),.I3(N_503),.LO(N_216_i));
defparam desc1303.INIT=16'h4414;
  LUT6_L desc1304(.I0(start_QR),.I1(state_8),.I2(row_sel_AQ[1:1]),.I3(row_sel_AQ[0:0]),.I4(N_706),.I5(N_676),.LO(N_220_i));
defparam desc1304.INIT=64'h0000000000000770;
  LUT6_L start_inner_prod_e(.I0(start_QR),.I1(state_8),.I2(start_inner_prod),.I3(un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_O6),.I4(N_706),.I5(N_676),.LO(start_inner_prod_0));
defparam start_inner_prod_e.INIT=64'hFFFFFFFFFFFF88B8;
  LUT6_L desc1305(.I0(col_sel_AQ2_int[1:1]),.I1(state[4:4]),.I2(state_8),.I3(N_495),.I4(N_106_1),.I5(N_106_2),.LO(j_RNO[1:1]));
defparam desc1305.INIT=64'hFFFFFFFFFFFF0200;
  LUT6_L desc1306(.I0(mult_counter[2:2]),.I1(state_8),.I2(col_sel_AQ_int[0:0]),.I3(N_495),.I4(N_686),.I5(N_527),.LO(N_231_i));
defparam desc1306.INIT=64'h0000111100003313;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 un1_state_23_0_0_o2_lut6_2_o6(.I0(done_inner_prod),.I1(state[2:2]),.I2(state_5),.I3(done_inv_sqrt),.O(un1_state_23_0_0_o2_lut6_2_O6));
defparam un1_state_23_0_0_o2_lut6_2_o6.INIT=16'hF888;
  LUT5 un1_state_23_0_0_o2_lut6_2_o5(.I0(mult_counter[0:0]),.I1(done_inner_prod),.I2(state[2:2]),.I3(state_5),.I4(done_inv_sqrt),.O(N_513_i));
defparam un1_state_23_0_0_o2_lut6_2_o5.INIT=32'h002A2A2A;
  LUT2 un1_state_25_0_0_o2_lut6_2_o6(.I0(state_5),.I1(state_8),.O(N_653));
defparam un1_state_25_0_0_o2_lut6_2_o6.INIT=4'hE;
  LUT5 un1_state_25_0_0_o2_lut6_2_o5(.I0(state[6:6]),.I1(done_inner_prod),.I2(state_5),.I3(start_inv_sqrt),.I4(state_8),.O(start_inv_sqrt_0));
defparam un1_state_25_0_0_o2_lut6_2_o5.INIT=32'hAAAAAFA8;
  LUT2 un1_state_10_0_o6_0_o2_lut6_2_o6(.I0(state[1:1]),.I1(state[4:4]),.O(un1_state_10_0_o6_0_o2_lut6_2_O6));
defparam un1_state_10_0_o6_0_o2_lut6_2_o6.INIT=4'hE;
  LUT4 un1_state_10_0_o6_0_o2_lut6_2_o5(.I0(state[1:1]),.I1(done_inner_prod),.I2(state[2:2]),.I3(mult_counter[2:2]),.O(state_ns[7:7]));
defparam un1_state_10_0_o6_0_o2_lut6_2_o5.INIT=16'hC0EA;
  LUT2 un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_o6(.I0(state_3),.I1(state[7:7]),.O(un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_O6));
defparam un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_o6.INIT=4'hE;
  LUT5 un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_o5(.I0(state_3),.I1(state[7:7]),.I2(state_8),.I3(in_b_inner_prod_sel),.I4(N_652),.O(in_b_inner_prod_sel_0));
defparam un1_state_1_sqmuxa_3_0_o6_0_o2_lut6_2_o5.INIT=32'hFEFEFFEE;
  LUT2 desc1307(.I0(col_sel_AQ2_int[0:0]),.I1(state[1:1]),.O(N_495));
defparam desc1307.INIT=4'h7;
  LUT5 desc1308(.I0(col_sel_AQ2_int[0:0]),.I1(col_sel_AQ2_int[1:1]),.I2(state[1:1]),.I3(red_mat_reg),.I4(mult_counter[2:2]),.O(N_503));
defparam desc1308.INIT=32'h5F7FFFFF;
  LUT2 un1_state_1_sqmuxa_4_0_0_a3_lut6_2_o6(.I0(state[1:1]),.I1(mult_counter[2:2]),.O(N_706));
defparam un1_state_1_sqmuxa_4_0_0_a3_lut6_2_o6.INIT=4'h8;
  LUT5 un1_state_1_sqmuxa_4_0_0_a3_lut6_2_o5(.I0(col_sel_AQ2_int[0:0]),.I1(state[1:1]),.I2(state[4:4]),.I3(mult_counter[2:2]),.I4(col_sel_AQ_int[0:0]),.O(N_686));
defparam un1_state_1_sqmuxa_4_0_0_a3_lut6_2_o5.INIT=32'h11550155;
  LUT2 desc1309(.I0(state[4:4]),.I1(mult_counter[2:2]),.O(N_662));
defparam desc1309.INIT=4'h2;
  LUT4 desc1310(.I0(state_3),.I1(state[7:7]),.I2(state[4:4]),.I3(state[1:1]),.O(N_201_2));
defparam desc1310.INIT=16'hFFFE;
  LUT2 row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_o6(.I0(state_5),.I1(done_inv_sqrt),.O(row_sel_R_0_sqmuxa));
defparam row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_o6.INIT=4'h8;
  LUT5 row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_o5(.I0(done_inner_prod),.I1(state[2:2]),.I2(state_5),.I3(state_8),.I4(done_inv_sqrt),.O(row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_O5));
defparam row_sel_R_0_sqmuxa_0_a6_0_a2_lut6_2_o5.INIT=32'hFFF8FF88;
  LUT2 desc1311(.I0(rst),.I1(state[4:4]),.O(N_512_i));
defparam desc1311.INIT=4'h4;
  LUT4 desc1312(.I0(state[4:4]),.I1(mult_counter[2:2]),.I2(state_5),.I3(done_inv_sqrt),.O(state_ns[4:4]));
defparam desc1312.INIT=16'hF222;
  LUT3 desc1313(.I0(red_mat_reg),.I1(row_sel_AQ[1:1]),.I2(row_sel_AQ[0:0]),.O(N_526));
defparam desc1313.INIT=8'h1F;
  LUT3 desc1314(.I0(col_sel_AQ2_int[0:0]),.I1(col_sel_AQ2_int[1:1]),.I2(red_mat_reg),.O(state_ns_2_tz[5:5]));
defparam desc1314.INIT=8'h57;
  LUT5 desc1315(.I0(state[4:4]),.I1(red_mat_reg),.I2(mult_counter[2:2]),.I3(col_sel_AQ_int[1:1]),.I4(col_sel_AQ_int[0:0]),.O(N_676));
defparam desc1315.INIT=32'h0020A0A0;
  LUT5 desc1316(.I0(state[4:4]),.I1(red_mat_reg),.I2(mult_counter[2:2]),.I3(col_sel_AQ_int[1:1]),.I4(col_sel_AQ_int[0:0]),.O(N_210_i));
defparam desc1316.INIT=32'hA0800000;
endmodule
module qr_decomp_ctl_mux_inj (single_in_R_sel,single_in_R_sel_0,w_col_sel_AQ_int,col_sel_AQ,wr_en_AQ_sel,w_col_sel_AQ_mux_i_m3_lut6_2_O6,w_col_sel_AQ_mux_i_m3_lut6_2_O5,col_sel_AQ2_int,col_sel_AQ2_mux_i_m3_lut6_2_O6,col_sel_AQ2_mux_i_m3_lut6_2_O5,state_0,state_2,state_5,wr_en_AQ_sel_0,col_sel_R,col_sel_R_int,col_sel_R_mux_i_m3_lut6_2_O6,col_sel_R_mux_i_m3_lut6_2_O5,in_a_r_reg_0_0,in_a_r_reg_0_11,out_r_vec_sub_0,in_a_i_reg_1,vec_in_AQ_sel,in_a_r_reg_3,in_a_i_reg_0,in_a_i_reg_3,in_a_r_reg_1,pre_out_4,pre_out_0,in_a_r_reg_2,pre_out_5,pre_out_1,in_a_i_reg_2,pre_out_6,pre_out_3_9,pre_out_3_1,pre_out_3_7,pre_out_3_3,pre_out_3_8,pre_out_3_5,pre_out_3_6,pre_out_3_0,pre_out_2,out_inner_prod_i,pre_out_10,pre_out_9,pre_out_0_d0,pre_out_1_d0,pre_out_3_d0,pre_out_6_d0,pre_out_7,pre_out_8,pre_out_5_d0,pre_out_4_d0,pre_out_2_d0,pre_out_18,pre_out_19,pre_out_20,pre_out_21,pre_out_reg,out_r_vec_mult_2,vec_in_r_AQ_mux_2,out_r_vec_mult_1,vec_in_r_AQ_mux_1,pre_out_i_m,out_i_vec_mult_3,pre_out_i_m_1,vec_in_i_AQ_mux_3,output_iv,out_i_vec_mult_0,vec_in_i_AQ_mux_0_11,vec_in_i_AQ_mux_0_1,vec_in_i_AQ_mux_0_5,vec_in_i_AQ_mux_0_0,vec_in_i_AQ_mux_0_8,vec_in_i_AQ_mux_0_10,vec_in_i_AQ_mux_0_7,vec_in_i_AQ_mux_0_6,vec_in_i_AQ_mux_0_9,vec_in_i_AQ_mux_0_4,out_r_vec_mult_0,output_iv_0_2,output_iv_0_4,output_iv_0_1,output_iv_0_0,output_iv_0_9,output_iv_0_6,output_iv_0_8,output_iv_0_3,output_iv_0_7,vec_in_r_AQ_mux_0_10,vec_in_r_AQ_mux_0_2,vec_in_r_AQ_mux_0_4,vec_in_r_AQ_mux_0_3,vec_in_r_AQ_mux_0_6,vec_in_r_AQ_mux_0_1,vec_in_r_AQ_mux_0_9,vec_in_r_AQ_mux_0_8,vec_in_r_AQ_mux_0_0,vec_in_r_AQ_mux_0_7,pre_out_i_m_0_0,pre_out_i_m_0_6,pre_out_i_m_0_4,pre_out_i_m_0_1,in_A_r,out_r_vec_mult_3,pre_out_i_m_2,vec_in_r_AQ_mux_3,out_i_vec_mult_2,pre_out_i_m_3,vec_in_i_AQ_mux_2,in_A_i,out_i_vec_mult_1,pre_out_i_m_4,vec_in_i_AQ_mux_1,un8_rnd_out_P,single_in_r_R_mux,out_inner_prod_r,un8_rnd_out,N_390_i,N_393_i,done_inv_sqrt,N_391_i,N_394_i,N_396_i,N_395_i,N_397_i,N_398_i,N_400_i,N_399_i,N_401_i,wr_en_AQ_int,wr_A_QR,start_QR,wr_en_AQ_mux_i_m3_lut6_2_O6,N_501,N_392_i,PATTERNDETECT_32,N_500,N_508,N_507,N_506,N_505,un5_output,un5_output_0,un5_output_1,un5_output_2,un5_output_3,un5_output_4,N_389_i,N_388_i,N_387_i,N_386_i,N_385_i,N_384_i,N_383_i,N_34_i,N_32_i,N_30_i,N_28_i);
input single_in_R_sel ;
output single_in_R_sel_0 ;
input [1:0] w_col_sel_AQ_int ;
input [1:0] col_sel_AQ ;
input wr_en_AQ_sel ;
output w_col_sel_AQ_mux_i_m3_lut6_2_O6 ;
output w_col_sel_AQ_mux_i_m3_lut6_2_O5 ;
input [1:0] col_sel_AQ2_int ;
output col_sel_AQ2_mux_i_m3_lut6_2_O6 ;
output col_sel_AQ2_mux_i_m3_lut6_2_O5 ;
input state_0 ;
input state_2 ;
input state_5 ;
output wr_en_AQ_sel_0 ;
input [1:0] col_sel_R ;
input [1:0] col_sel_R_int ;
output col_sel_R_mux_i_m3_lut6_2_O6 ;
output col_sel_R_mux_i_m3_lut6_2_O5 ;
input in_a_r_reg_0_0 ;
input in_a_r_reg_0_11 ;
output [11:11] out_r_vec_sub_0 ;
input [11:11] in_a_i_reg_1 ;
input [1:0] vec_in_AQ_sel ;
input [11:11] in_a_r_reg_3 ;
input [11:11] in_a_i_reg_0 ;
input [11:11] in_a_i_reg_3 ;
input [11:11] in_a_r_reg_1 ;
input [11:11] pre_out_4 ;
input [11:1] pre_out_0 ;
input [11:11] in_a_r_reg_2 ;
input [11:11] pre_out_5 ;
input [11:1] pre_out_1 ;
input [11:11] in_a_i_reg_2 ;
input [11:11] pre_out_6 ;
input pre_out_3_9 ;
input pre_out_3_1 ;
input pre_out_3_7 ;
input pre_out_3_3 ;
input pre_out_3_8 ;
input pre_out_3_5 ;
input pre_out_3_6 ;
input pre_out_3_0 ;
input [11:1] pre_out_2 ;
input [11:0] out_inner_prod_i ;
input pre_out_10 ;
input pre_out_9 ;
input pre_out_0_d0 ;
input pre_out_1_d0 ;
input pre_out_3_d0 ;
input pre_out_6_d0 ;
input pre_out_7 ;
input pre_out_8 ;
input pre_out_5_d0 ;
input pre_out_4_d0 ;
input pre_out_2_d0 ;
input pre_out_18 ;
input pre_out_19 ;
input pre_out_20 ;
input pre_out_21 ;
input [23:23] pre_out_reg ;
input [11:0] out_r_vec_mult_2 ;
output [11:0] vec_in_r_AQ_mux_2 ;
input [11:0] out_r_vec_mult_1 ;
output [11:0] vec_in_r_AQ_mux_1 ;
input [10:0] pre_out_i_m ;
input [11:0] out_i_vec_mult_3 ;
input pre_out_i_m_1 ;
output [11:0] vec_in_i_AQ_mux_3 ;
input [10:0] output_iv ;
input [11:0] out_i_vec_mult_0 ;
output vec_in_i_AQ_mux_0_11 ;
output vec_in_i_AQ_mux_0_1 ;
output vec_in_i_AQ_mux_0_5 ;
output vec_in_i_AQ_mux_0_0 ;
output vec_in_i_AQ_mux_0_8 ;
output vec_in_i_AQ_mux_0_10 ;
output vec_in_i_AQ_mux_0_7 ;
output vec_in_i_AQ_mux_0_6 ;
output vec_in_i_AQ_mux_0_9 ;
output vec_in_i_AQ_mux_0_4 ;
input [11:0] out_r_vec_mult_0 ;
input output_iv_0_2 ;
input output_iv_0_4 ;
input output_iv_0_1 ;
input output_iv_0_0 ;
input output_iv_0_9 ;
input output_iv_0_6 ;
input output_iv_0_8 ;
input output_iv_0_3 ;
input output_iv_0_7 ;
output vec_in_r_AQ_mux_0_10 ;
output vec_in_r_AQ_mux_0_2 ;
output vec_in_r_AQ_mux_0_4 ;
output vec_in_r_AQ_mux_0_3 ;
output vec_in_r_AQ_mux_0_6 ;
output vec_in_r_AQ_mux_0_1 ;
output vec_in_r_AQ_mux_0_9 ;
output vec_in_r_AQ_mux_0_8 ;
output vec_in_r_AQ_mux_0_0 ;
output vec_in_r_AQ_mux_0_7 ;
input pre_out_i_m_0_0 ;
input pre_out_i_m_0_6 ;
input pre_out_i_m_0_4 ;
input pre_out_i_m_0_1 ;
input [47:0] in_A_r ;
input [11:0] out_r_vec_mult_3 ;
input pre_out_i_m_2 ;
output [11:0] vec_in_r_AQ_mux_3 ;
input [11:0] out_i_vec_mult_2 ;
input pre_out_i_m_3 ;
output [11:0] vec_in_i_AQ_mux_2 ;
input [47:0] in_A_i ;
input [11:0] out_i_vec_mult_1 ;
input pre_out_i_m_4 ;
output [11:0] vec_in_i_AQ_mux_1 ;
input [19:19] un8_rnd_out_P ;
output [11:11] single_in_r_R_mux ;
input [11:0] out_inner_prod_r ;
input [10:0] un8_rnd_out ;
output N_390_i ;
output N_393_i ;
input done_inv_sqrt ;
output N_391_i ;
output N_394_i ;
output N_396_i ;
output N_395_i ;
output N_397_i ;
output N_398_i ;
output N_400_i ;
output N_399_i ;
output N_401_i ;
input wr_en_AQ_int ;
input wr_A_QR ;
input start_QR ;
output wr_en_AQ_mux_i_m3_lut6_2_O6 ;
output N_501 ;
output N_392_i ;
input PATTERNDETECT_32 ;
input N_500 ;
output N_508 ;
output N_507 ;
output N_506 ;
output N_505 ;
input un5_output ;
input un5_output_0 ;
input un5_output_1 ;
input un5_output_2 ;
input un5_output_3 ;
input un5_output_4 ;
output N_389_i ;
output N_388_i ;
output N_387_i ;
output N_386_i ;
output N_385_i ;
output N_384_i ;
output N_383_i ;
output N_34_i ;
output N_32_i ;
output N_30_i ;
output N_28_i ;
wire state_0 ;
wire state_2 ;
wire state_5 ;
wire in_a_r_reg_0_0 ;
wire in_a_r_reg_0_11 ;
wire pre_out_3_9 ;
wire pre_out_3_1 ;
wire pre_out_3_7 ;
wire pre_out_3_3 ;
wire pre_out_3_8 ;
wire pre_out_3_5 ;
wire pre_out_3_6 ;
wire pre_out_3_0 ;
wire pre_out_10 ;
wire pre_out_9 ;
wire pre_out_0_d0 ;
wire pre_out_1_d0 ;
wire pre_out_3_d0 ;
wire pre_out_6_d0 ;
wire pre_out_7 ;
wire pre_out_8 ;
wire pre_out_5_d0 ;
wire pre_out_4_d0 ;
wire pre_out_2_d0 ;
wire pre_out_18 ;
wire pre_out_19 ;
wire pre_out_20 ;
wire pre_out_21 ;
wire vec_in_i_AQ_mux_0_11 ;
wire vec_in_i_AQ_mux_0_1 ;
wire vec_in_i_AQ_mux_0_5 ;
wire vec_in_i_AQ_mux_0_0 ;
wire vec_in_i_AQ_mux_0_8 ;
wire vec_in_i_AQ_mux_0_10 ;
wire vec_in_i_AQ_mux_0_7 ;
wire vec_in_i_AQ_mux_0_6 ;
wire vec_in_i_AQ_mux_0_9 ;
wire vec_in_i_AQ_mux_0_4 ;
wire output_iv_0_2 ;
wire output_iv_0_4 ;
wire output_iv_0_1 ;
wire output_iv_0_0 ;
wire output_iv_0_9 ;
wire output_iv_0_6 ;
wire output_iv_0_8 ;
wire output_iv_0_3 ;
wire output_iv_0_7 ;
wire vec_in_r_AQ_mux_0_10 ;
wire vec_in_r_AQ_mux_0_2 ;
wire vec_in_r_AQ_mux_0_4 ;
wire vec_in_r_AQ_mux_0_3 ;
wire vec_in_r_AQ_mux_0_6 ;
wire vec_in_r_AQ_mux_0_1 ;
wire vec_in_r_AQ_mux_0_9 ;
wire vec_in_r_AQ_mux_0_8 ;
wire vec_in_r_AQ_mux_0_0 ;
wire vec_in_r_AQ_mux_0_7 ;
wire pre_out_i_m_0_0 ;
wire pre_out_i_m_0_6 ;
wire pre_out_i_m_0_4 ;
wire pre_out_i_m_0_1 ;
wire N_390_i ;
wire N_393_i ;
wire done_inv_sqrt ;
wire N_391_i ;
wire N_394_i ;
wire N_396_i ;
wire N_395_i ;
wire N_397_i ;
wire N_398_i ;
wire N_400_i ;
wire N_399_i ;
wire N_401_i ;
wire wr_en_AQ_int ;
wire wr_A_QR ;
wire start_QR ;
wire wr_en_AQ_mux_i_m3_lut6_2_O6 ;
wire N_501 ;
wire N_392_i ;
wire PATTERNDETECT_32 ;
wire N_500 ;
wire N_508 ;
wire N_507 ;
wire N_506 ;
wire N_505 ;
wire un5_output ;
wire un5_output_0 ;
wire un5_output_1 ;
wire un5_output_2 ;
wire un5_output_3 ;
wire un5_output_4 ;
wire N_389_i ;
wire N_388_i ;
wire N_387_i ;
wire N_386_i ;
wire N_385_i ;
wire N_384_i ;
wire N_383_i ;
wire N_34_i ;
wire N_32_i ;
wire N_30_i ;
wire N_28_i ;
wire GND ;
wire VCC ;
wire N_161 ;
wire N_162 ;
wire N_163 ;
wire N_164 ;
wire N_165 ;
wire N_148 ;
wire N_166 ;
wire N_167 ;
wire N_168 ;
wire N_169 ;
wire N_149 ;
wire N_150 ;
wire N_151 ;
wire N_152 ;
wire N_153 ;
wire N_154 ;
wire N_155 ;
wire N_143 ;
wire N_156 ;
wire N_157 ;
wire N_37 ;
wire N_38 ;
wire N_39 ;
wire N_40 ;
wire N_41 ;
wire N_50 ;
wire N_60 ;
wire N_66 ;
wire N_61 ;
wire N_62 ;
wire N_64 ;
wire N_65 ;
wire N_68 ;
wire N_69 ;
wire N_48 ;
wire N_49 ;
wire N_51 ;
wire N_52 ;
wire N_54 ;
wire N_55 ;
wire N_56 ;
wire N_57 ;
wire N_42 ;
wire N_43 ;
wire N_44 ;
wire N_45 ;
wire N_160 ;
wire N_95 ;
wire N_122 ;
// instances
  LUT6 desc1091(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_169),.I4(pre_out_9),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[10:10]));
defparam desc1091.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1092(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_160),.I4(pre_out_0_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[1:1]));
defparam desc1092.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1093(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_161),.I4(pre_out_1_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[2:2]));
defparam desc1093.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1094(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_163),.I4(pre_out_3_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[4:4]));
defparam desc1094.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1095(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_166),.I4(pre_out_6_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[7:7]));
defparam desc1095.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1096(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_167),.I4(pre_out_7),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[8:8]));
defparam desc1096.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1097(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_168),.I4(pre_out_8),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[9:9]));
defparam desc1097.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1098(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_165),.I4(pre_out_5_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[6:6]));
defparam desc1098.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1099(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_164),.I4(pre_out_4_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[5:5]));
defparam desc1099.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1100(.I0(out_i_vec_mult_1[11:11]),.I1(in_a_i_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_162),.I4(pre_out_2_d0),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[3:3]));
defparam desc1100.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1101(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_41),.I4(pre_out_0[6:6]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[6:6]));
defparam desc1101.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1102(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_44),.I4(pre_out_0[9:9]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[9:9]));
defparam desc1102.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1103(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_37),.I4(pre_out_0[2:2]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[2:2]));
defparam desc1103.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1104(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_39),.I4(pre_out_0[4:4]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[4:4]));
defparam desc1104.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1105(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_40),.I4(pre_out_0[5:5]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[5:5]));
defparam desc1105.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1106(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_45),.I4(pre_out_0[10:10]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[10:10]));
defparam desc1106.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1107(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_38),.I4(pre_out_0[3:3]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[3:3]));
defparam desc1107.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1108(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_42),.I4(pre_out_0[7:7]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[7:7]));
defparam desc1108.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1109(.I0(out_r_vec_mult_3[11:11]),.I1(in_a_r_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_43),.I4(pre_out_0[8:8]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[8:8]));
defparam desc1109.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1110(.I0(in_A_i[47:47]),.I1(out_i_vec_mult_0[11:11]),.I2(in_a_i_reg_0[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_2[11:11]),.O(vec_in_i_AQ_mux_0_11));
defparam desc1110.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1111(.I0(in_A_r[47:47]),.I1(out_r_vec_mult_0[11:11]),.I2(in_a_r_reg_0_11),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_10),.O(vec_in_r_AQ_mux_0_10));
defparam desc1111.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1112(.I0(out_i_vec_mult_3[11:11]),.I1(in_a_i_reg_3[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_143),.I4(pre_out_1[8:8]),.I5(pre_out_3_9),.O(vec_in_i_AQ_mux_3[8:8]));
defparam desc1112.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1113(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_62),.I4(pre_out_1[3:3]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[3:3]));
defparam desc1113.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1114(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_65),.I4(pre_out_1[6:6]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[6:6]));
defparam desc1114.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1115(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_64),.I4(pre_out_1[5:5]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[5:5]));
defparam desc1115.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1116(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_69),.I4(pre_out_1[10:10]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[10:10]));
defparam desc1116.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1117(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_60),.I4(pre_out_0[1:1]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[1:1]));
defparam desc1117.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1118(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_68),.I4(pre_out_1[9:9]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[9:9]));
defparam desc1118.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1119(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_61),.I4(pre_out_1[2:2]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[2:2]));
defparam desc1119.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1120(.I0(out_r_vec_mult_1[11:11]),.I1(in_a_r_reg_1[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_66),.I4(pre_out_1[7:7]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[7:7]));
defparam desc1120.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1121(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_51),.I4(pre_out_1[4:4]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[4:4]));
defparam desc1121.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1122(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_55),.I4(pre_out_2[8:8]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[8:8]));
defparam desc1122.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1123(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_54),.I4(pre_out_2[7:7]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[7:7]));
defparam desc1123.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1124(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_48),.I4(pre_out_1[1:1]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[1:1]));
defparam desc1124.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1125(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_50),.I4(pre_out_2[3:3]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[3:3]));
defparam desc1125.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1126(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_57),.I4(pre_out_2[10:10]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[10:10]));
defparam desc1126.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1127(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_52),.I4(pre_out_2[5:5]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[5:5]));
defparam desc1127.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1128(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_49),.I4(pre_out_2[2:2]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[2:2]));
defparam desc1128.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1129(.I0(out_r_vec_mult_2[11:11]),.I1(in_a_r_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_56),.I4(pre_out_2[9:9]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[9:9]));
defparam desc1129.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1130(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_150),.I4(pre_out_3_1),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[3:3]));
defparam desc1130.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1131(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_156),.I4(pre_out_3_7),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[9:9]));
defparam desc1131.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1132(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_152),.I4(pre_out_3_3),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[5:5]));
defparam desc1132.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1133(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_157),.I4(pre_out_3_8),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[10:10]));
defparam desc1133.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1134(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_151),.I4(pre_out_2[4:4]),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[4:4]));
defparam desc1134.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1135(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_154),.I4(pre_out_3_5),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[7:7]));
defparam desc1135.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1136(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_155),.I4(pre_out_3_6),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[8:8]));
defparam desc1136.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1137(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_149),.I4(pre_out_3_0),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[2:2]));
defparam desc1137.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1138(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_153),.I4(pre_out_2[6:6]),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[6:6]));
defparam desc1138.INIT=64'hFFF02F20BFB00F00;
  LUT6 desc1139(.I0(out_i_vec_mult_2[11:11]),.I1(in_a_i_reg_2[11:11]),.I2(vec_in_AQ_sel[1:1]),.I3(N_148),.I4(pre_out_2[1:1]),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[1:1]));
defparam desc1139.INIT=64'hFFF02F20BFB00F00;
  LUT3 desc1140(.I0(in_A_i[25:25]),.I1(out_i_vec_mult_1[1:1]),.I2(vec_in_AQ_sel[0:0]),.O(N_160));
defparam desc1140.INIT=8'hCA;
  LUT2 N_392_i_c(.I0(out_inner_prod_i[2:2]),.I1(single_in_R_sel),.O(N_392_i));
defparam N_392_i_c.INIT=4'h8;
  LUT6 single_in_r_R_mux_i_a3_a(.I0(single_in_R_sel),.I1(pre_out_18),.I2(pre_out_19),.I3(pre_out_20),.I4(pre_out_21),.I5(PATTERNDETECT_32),.O(N_95));
defparam single_in_r_R_mux_i_a3_a.INIT=64'h1555555500000000;
  LUT6 desc1141(.I0(single_in_R_sel),.I1(pre_out_reg[23:23]),.I2(pre_out_18),.I3(pre_out_19),.I4(pre_out_20),.I5(pre_out_21),.O(N_122));
defparam desc1141.INIT=64'h4444444444444445;
  LUT5 desc1142(.I0(in_A_r[42:42]),.I1(out_r_vec_mult_0[6:6]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(N_500),.O(N_508));
defparam desc1142.INIT=32'h00CAFFCA;
  LUT5 desc1143(.I0(in_A_r[36:36]),.I1(out_r_vec_mult_0[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(N_501),.O(N_507));
defparam desc1143.INIT=32'h00CAFFCA;
  LUT5 desc1144(.I0(in_A_i[39:39]),.I1(out_i_vec_mult_0[3:3]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[3:3]),.O(N_506));
defparam desc1144.INIT=32'h00CAFFCA;
  LUT5 desc1145(.I0(in_A_i[38:38]),.I1(out_i_vec_mult_0[2:2]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[2:2]),.O(N_505));
defparam desc1145.INIT=32'h00CAFFCA;
  LUT5 desc1146(.I0(in_A_r[39:39]),.I1(out_r_vec_mult_0[3:3]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_2),.O(vec_in_r_AQ_mux_0_2));
defparam desc1146.INIT=32'h00CAFFCA;
  LUT6 desc1147(.I0(in_A_r[11:11]),.I1(out_r_vec_mult_3[11:11]),.I2(in_a_r_reg_3[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_1[11:11]),.O(vec_in_r_AQ_mux_3[11:11]));
defparam desc1147.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1148(.I0(in_A_r[23:23]),.I1(out_r_vec_mult_2[11:11]),.I2(in_a_r_reg_2[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_5[11:11]),.O(vec_in_r_AQ_mux_2[11:11]));
defparam desc1148.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1149(.I0(in_A_r[18:18]),.I1(out_r_vec_mult_2[6:6]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[6:6]),.I5(un5_output),.O(vec_in_r_AQ_mux_2[6:6]));
defparam desc1149.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1150(.I0(in_A_r[12:12]),.I1(out_r_vec_mult_2[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[0:0]),.I5(un5_output),.O(vec_in_r_AQ_mux_2[0:0]));
defparam desc1150.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1151(.I0(in_A_r[35:35]),.I1(out_r_vec_mult_1[11:11]),.I2(in_a_r_reg_1[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_4[11:11]),.O(vec_in_r_AQ_mux_1[11:11]));
defparam desc1151.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1152(.I0(in_A_r[32:32]),.I1(out_r_vec_mult_1[8:8]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[8:8]),.I5(un5_output_0),.O(vec_in_r_AQ_mux_1[8:8]));
defparam desc1152.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1153(.I0(in_A_r[28:28]),.I1(out_r_vec_mult_1[4:4]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[4:4]),.I5(un5_output_0),.O(vec_in_r_AQ_mux_1[4:4]));
defparam desc1153.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1154(.I0(in_A_r[24:24]),.I1(out_r_vec_mult_1[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_0_0),.I5(un5_output_0),.O(vec_in_r_AQ_mux_1[0:0]));
defparam desc1154.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1155(.I0(in_A_i[11:11]),.I1(out_i_vec_mult_3[11:11]),.I2(in_a_i_reg_3[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_3_9),.O(vec_in_i_AQ_mux_3[11:11]));
defparam desc1155.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1156(.I0(in_A_i[10:10]),.I1(out_i_vec_mult_3[10:10]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[10:10]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[10:10]));
defparam desc1156.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1157(.I0(in_A_i[9:9]),.I1(out_i_vec_mult_3[9:9]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[9:9]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[9:9]));
defparam desc1157.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1158(.I0(in_A_i[7:7]),.I1(out_i_vec_mult_3[7:7]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[7:7]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[7:7]));
defparam desc1158.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1159(.I0(in_A_i[6:6]),.I1(out_i_vec_mult_3[6:6]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_0_6),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[6:6]));
defparam desc1159.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1160(.I0(in_A_i[5:5]),.I1(out_i_vec_mult_3[5:5]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[5:5]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[5:5]));
defparam desc1160.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1161(.I0(in_A_i[4:4]),.I1(out_i_vec_mult_3[4:4]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_0_4),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[4:4]));
defparam desc1161.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1162(.I0(in_A_i[3:3]),.I1(out_i_vec_mult_3[3:3]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[3:3]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[3:3]));
defparam desc1162.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1163(.I0(in_A_i[2:2]),.I1(out_i_vec_mult_3[2:2]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[2:2]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[2:2]));
defparam desc1163.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1164(.I0(in_A_i[1:1]),.I1(out_i_vec_mult_3[1:1]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m[1:1]),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[1:1]));
defparam desc1164.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1165(.I0(in_A_i[0:0]),.I1(out_i_vec_mult_3[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_1),.I5(un5_output_1),.O(vec_in_i_AQ_mux_3[0:0]));
defparam desc1165.INIT=64'h00CAFFCA00CA00CA;
  LUT5 desc1166(.I0(in_A_i[37:37]),.I1(out_i_vec_mult_0[1:1]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[1:1]),.O(vec_in_i_AQ_mux_0_1));
defparam desc1166.INIT=32'h00CAFFCA;
  LUT5 desc1167(.I0(in_A_r[41:41]),.I1(out_r_vec_mult_0[5:5]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[5:5]),.O(vec_in_r_AQ_mux_0_4));
defparam desc1167.INIT=32'h00CAFFCA;
  LUT5 desc1168(.I0(in_A_r[40:40]),.I1(out_r_vec_mult_0[4:4]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[4:4]),.O(vec_in_r_AQ_mux_0_3));
defparam desc1168.INIT=32'h00CAFFCA;
  LUT5 desc1169(.I0(in_A_i[41:41]),.I1(out_i_vec_mult_0[5:5]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_4),.O(vec_in_i_AQ_mux_0_5));
defparam desc1169.INIT=32'h00CAFFCA;
  LUT5 desc1170(.I0(in_A_i[36:36]),.I1(out_i_vec_mult_0[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[0:0]),.O(vec_in_i_AQ_mux_0_0));
defparam desc1170.INIT=32'h00CAFFCA;
  LUT5 desc1171(.I0(in_A_r[43:43]),.I1(out_r_vec_mult_0[7:7]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[7:7]),.O(vec_in_r_AQ_mux_0_6));
defparam desc1171.INIT=32'h00CAFFCA;
  LUT5 desc1172(.I0(in_A_r[38:38]),.I1(out_r_vec_mult_0[2:2]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_1),.O(vec_in_r_AQ_mux_0_1));
defparam desc1172.INIT=32'h00CAFFCA;
  LUT5 desc1173(.I0(in_A_i[44:44]),.I1(out_i_vec_mult_0[8:8]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[8:8]),.O(vec_in_i_AQ_mux_0_8));
defparam desc1173.INIT=32'h00CAFFCA;
  LUT5 desc1174(.I0(in_A_r[46:46]),.I1(out_r_vec_mult_0[10:10]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[10:10]),.O(vec_in_r_AQ_mux_0_9));
defparam desc1174.INIT=32'h00CAFFCA;
  LUT5 desc1175(.I0(in_A_r[45:45]),.I1(out_r_vec_mult_0[9:9]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[9:9]),.O(vec_in_r_AQ_mux_0_8));
defparam desc1175.INIT=32'h00CAFFCA;
  LUT5 desc1176(.I0(in_A_r[37:37]),.I1(out_r_vec_mult_0[1:1]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_0),.O(vec_in_r_AQ_mux_0_0));
defparam desc1176.INIT=32'h00CAFFCA;
  LUT5 desc1177(.I0(in_A_i[46:46]),.I1(out_i_vec_mult_0[10:10]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_9),.O(vec_in_i_AQ_mux_0_10));
defparam desc1177.INIT=32'h00CAFFCA;
  LUT5 desc1178(.I0(in_A_i[43:43]),.I1(out_i_vec_mult_0[7:7]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_6),.O(vec_in_i_AQ_mux_0_7));
defparam desc1178.INIT=32'h00CAFFCA;
  LUT5 desc1179(.I0(in_A_i[42:42]),.I1(out_i_vec_mult_0[6:6]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv[6:6]),.O(vec_in_i_AQ_mux_0_6));
defparam desc1179.INIT=32'h00CAFFCA;
  LUT5 desc1180(.I0(in_A_i[45:45]),.I1(out_i_vec_mult_0[9:9]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_8),.O(vec_in_i_AQ_mux_0_9));
defparam desc1180.INIT=32'h00CAFFCA;
  LUT5 desc1181(.I0(in_A_i[40:40]),.I1(out_i_vec_mult_0[4:4]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_3),.O(vec_in_i_AQ_mux_0_4));
defparam desc1181.INIT=32'h00CAFFCA;
  LUT5 desc1182(.I0(in_A_r[44:44]),.I1(out_r_vec_mult_0[8:8]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(output_iv_0_7),.O(vec_in_r_AQ_mux_0_7));
defparam desc1182.INIT=32'h00CAFFCA;
  LUT6 desc1183(.I0(in_A_r[1:1]),.I1(out_r_vec_mult_3[1:1]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_0_1),.I5(un5_output_2),.O(vec_in_r_AQ_mux_3[1:1]));
defparam desc1183.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1184(.I0(in_A_r[0:0]),.I1(out_r_vec_mult_3[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(pre_out_i_m_2),.I5(un5_output_2),.O(vec_in_r_AQ_mux_3[0:0]));
defparam desc1184.INIT=64'h00CAFFCA00CA00CA;
  LUT6 desc1185(.I0(in_A_i[23:23]),.I1(out_i_vec_mult_2[11:11]),.I2(in_a_i_reg_2[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_6[11:11]),.O(vec_in_i_AQ_mux_2[11:11]));
defparam desc1185.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1186(.I0(in_A_i[12:12]),.I1(out_i_vec_mult_2[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(un5_output_3),.I5(pre_out_i_m_3),.O(vec_in_i_AQ_mux_2[0:0]));
defparam desc1186.INIT=64'h00CA00CAFFCA00CA;
  LUT6 desc1187(.I0(in_A_i[35:35]),.I1(out_i_vec_mult_1[11:11]),.I2(in_a_i_reg_1[11:11]),.I3(vec_in_AQ_sel[0:0]),.I4(vec_in_AQ_sel[1:1]),.I5(pre_out_0[11:11]),.O(vec_in_i_AQ_mux_1[11:11]));
defparam desc1187.INIT=64'hF3F3CCAA3030CCAA;
  LUT6 desc1188(.I0(in_A_i[24:24]),.I1(out_i_vec_mult_1[0:0]),.I2(vec_in_AQ_sel[0:0]),.I3(vec_in_AQ_sel[1:1]),.I4(un5_output_4),.I5(pre_out_i_m_4),.O(vec_in_i_AQ_mux_1[0:0]));
defparam desc1188.INIT=64'h00CA00CAFFCA00CA;
  LUT5 desc1189(.I0(single_in_R_sel),.I1(out_inner_prod_r[11:11]),.I2(un8_rnd_out_P[19:19]),.I3(N_122),.I4(N_95),.O(single_in_r_R_mux[11:11]));
defparam desc1189.INIT=32'hFFFFF888;
  LUT5 desc1190(.I0(out_inner_prod_r[10:10]),.I1(single_in_R_sel),.I2(un8_rnd_out[10:10]),.I3(N_122),.I4(N_95),.O(N_389_i));
defparam desc1190.INIT=32'h0000B0BB;
  LUT5 desc1191(.I0(out_inner_prod_r[9:9]),.I1(single_in_R_sel),.I2(un8_rnd_out[9:9]),.I3(N_122),.I4(N_95),.O(N_388_i));
defparam desc1191.INIT=32'h0000B0BB;
  LUT5 desc1192(.I0(out_inner_prod_r[8:8]),.I1(single_in_R_sel),.I2(un8_rnd_out[8:8]),.I3(N_122),.I4(N_95),.O(N_387_i));
defparam desc1192.INIT=32'h0000B0BB;
  LUT5 desc1193(.I0(out_inner_prod_r[7:7]),.I1(single_in_R_sel),.I2(un8_rnd_out[7:7]),.I3(N_122),.I4(N_95),.O(N_386_i));
defparam desc1193.INIT=32'h0000B0BB;
  LUT5 desc1194(.I0(out_inner_prod_r[6:6]),.I1(single_in_R_sel),.I2(un8_rnd_out[6:6]),.I3(N_122),.I4(N_95),.O(N_385_i));
defparam desc1194.INIT=32'h0000B0BB;
  LUT5 desc1195(.I0(out_inner_prod_r[5:5]),.I1(single_in_R_sel),.I2(un8_rnd_out[5:5]),.I3(N_122),.I4(N_95),.O(N_384_i));
defparam desc1195.INIT=32'h0000B0BB;
  LUT5 desc1196(.I0(out_inner_prod_r[4:4]),.I1(single_in_R_sel),.I2(un8_rnd_out[4:4]),.I3(N_122),.I4(N_95),.O(N_383_i));
defparam desc1196.INIT=32'h0000B0BB;
  LUT5 desc1197(.I0(out_inner_prod_r[3:3]),.I1(single_in_R_sel),.I2(un8_rnd_out[3:3]),.I3(N_122),.I4(N_95),.O(N_34_i));
defparam desc1197.INIT=32'h0000B0BB;
  LUT5 desc1198(.I0(out_inner_prod_r[2:2]),.I1(single_in_R_sel),.I2(un8_rnd_out[2:2]),.I3(N_122),.I4(N_95),.O(N_32_i));
defparam desc1198.INIT=32'h0000B0BB;
  LUT5 desc1199(.I0(out_inner_prod_r[1:1]),.I1(single_in_R_sel),.I2(un8_rnd_out[1:1]),.I3(N_122),.I4(N_95),.O(N_30_i));
defparam desc1199.INIT=32'h0000B0BB;
  LUT5 desc1200(.I0(out_inner_prod_r[0:0]),.I1(single_in_R_sel),.I2(un8_rnd_out[0:0]),.I3(N_122),.I4(N_95),.O(N_28_i));
defparam desc1200.INIT=32'h0000B0BB;
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT5 desc1201(.I0(out_r_vec_mult_0[0:0]),.I1(in_a_r_reg_0_0),.I2(out_r_vec_mult_0[11:11]),.I3(in_a_r_reg_0_11),.I4(pre_out_10),.O(N_501));
defparam desc1201.INIT=32'h99099F99;
  LUT3 desc1202(.I0(out_r_vec_mult_0[11:11]),.I1(in_a_r_reg_0_11),.I2(pre_out_10),.O(out_r_vec_sub_0[11:11]));
defparam desc1202.INIT=8'hD4;
  LUT3 desc1203(.I0(col_sel_R_int[0:0]),.I1(col_sel_R[0:0]),.I2(wr_en_AQ_sel),.O(col_sel_R_mux_i_m3_lut6_2_O6));
defparam desc1203.INIT=8'hAC;
  LUT3 desc1204(.I0(col_sel_R[1:1]),.I1(col_sel_R_int[1:1]),.I2(wr_en_AQ_sel),.O(col_sel_R_mux_i_m3_lut6_2_O5));
defparam desc1204.INIT=8'hCA;
  LUT3 wr_en_AQ_mux_i_m3_lut6_2_o6(.I0(wr_en_AQ_int),.I1(wr_A_QR),.I2(wr_en_AQ_sel),.O(wr_en_AQ_mux_i_m3_lut6_2_O6));
defparam wr_en_AQ_mux_i_m3_lut6_2_o6.INIT=8'hAC;
  LUT3 wr_en_AQ_mux_i_m3_lut6_2_o5(.I0(start_QR),.I1(state_5),.I2(wr_en_AQ_sel),.O(wr_en_AQ_sel_0));
defparam wr_en_AQ_mux_i_m3_lut6_2_o5.INIT=8'hB8;
  LUT3 desc1205(.I0(col_sel_AQ[0:0]),.I1(col_sel_AQ2_int[0:0]),.I2(wr_en_AQ_sel),.O(col_sel_AQ2_mux_i_m3_lut6_2_O6));
defparam desc1205.INIT=8'hCA;
  LUT3 desc1206(.I0(col_sel_AQ[1:1]),.I1(col_sel_AQ2_int[1:1]),.I2(wr_en_AQ_sel),.O(col_sel_AQ2_mux_i_m3_lut6_2_O5));
defparam desc1206.INIT=8'hCA;
  LUT3 desc1207(.I0(w_col_sel_AQ_int[0:0]),.I1(col_sel_AQ[0:0]),.I2(wr_en_AQ_sel),.O(w_col_sel_AQ_mux_i_m3_lut6_2_O6));
defparam desc1207.INIT=8'hAC;
  LUT3 desc1208(.I0(w_col_sel_AQ_int[1:1]),.I1(col_sel_AQ[1:1]),.I2(wr_en_AQ_sel),.O(w_col_sel_AQ_mux_i_m3_lut6_2_O5));
defparam desc1208.INIT=8'hAC;
  LUT3 desc1209(.I0(in_A_r[9:9]),.I1(out_r_vec_mult_3[9:9]),.I2(vec_in_AQ_sel[0:0]),.O(N_44));
defparam desc1209.INIT=8'hCA;
  LUT3 desc1210(.I0(in_A_r[10:10]),.I1(out_r_vec_mult_3[10:10]),.I2(vec_in_AQ_sel[0:0]),.O(N_45));
defparam desc1210.INIT=8'hCA;
  LUT3 desc1211(.I0(in_A_r[7:7]),.I1(out_r_vec_mult_3[7:7]),.I2(vec_in_AQ_sel[0:0]),.O(N_42));
defparam desc1211.INIT=8'hCA;
  LUT3 desc1212(.I0(in_A_r[8:8]),.I1(out_r_vec_mult_3[8:8]),.I2(vec_in_AQ_sel[0:0]),.O(N_43));
defparam desc1212.INIT=8'hCA;
  LUT3 desc1213(.I0(in_A_r[21:21]),.I1(out_r_vec_mult_2[9:9]),.I2(vec_in_AQ_sel[0:0]),.O(N_56));
defparam desc1213.INIT=8'hCA;
  LUT3 desc1214(.I0(in_A_r[22:22]),.I1(out_r_vec_mult_2[10:10]),.I2(vec_in_AQ_sel[0:0]),.O(N_57));
defparam desc1214.INIT=8'hCA;
  LUT3 desc1215(.I0(in_A_r[19:19]),.I1(out_r_vec_mult_2[7:7]),.I2(vec_in_AQ_sel[0:0]),.O(N_54));
defparam desc1215.INIT=8'hCA;
  LUT3 desc1216(.I0(in_A_r[20:20]),.I1(out_r_vec_mult_2[8:8]),.I2(vec_in_AQ_sel[0:0]),.O(N_55));
defparam desc1216.INIT=8'hCA;
  LUT3 desc1217(.I0(in_A_r[16:16]),.I1(out_r_vec_mult_2[4:4]),.I2(vec_in_AQ_sel[0:0]),.O(N_51));
defparam desc1217.INIT=8'hCA;
  LUT3 desc1218(.I0(in_A_r[17:17]),.I1(out_r_vec_mult_2[5:5]),.I2(vec_in_AQ_sel[0:0]),.O(N_52));
defparam desc1218.INIT=8'hCA;
  LUT3 desc1219(.I0(in_A_r[13:13]),.I1(out_r_vec_mult_2[1:1]),.I2(vec_in_AQ_sel[0:0]),.O(N_48));
defparam desc1219.INIT=8'hCA;
  LUT3 desc1220(.I0(in_A_r[14:14]),.I1(out_r_vec_mult_2[2:2]),.I2(vec_in_AQ_sel[0:0]),.O(N_49));
defparam desc1220.INIT=8'hCA;
  LUT3 desc1221(.I0(in_A_r[33:33]),.I1(out_r_vec_mult_1[9:9]),.I2(vec_in_AQ_sel[0:0]),.O(N_68));
defparam desc1221.INIT=8'hCA;
  LUT3 desc1222(.I0(in_A_r[34:34]),.I1(out_r_vec_mult_1[10:10]),.I2(vec_in_AQ_sel[0:0]),.O(N_69));
defparam desc1222.INIT=8'hCA;
  LUT3 desc1223(.I0(in_A_r[29:29]),.I1(out_r_vec_mult_1[5:5]),.I2(vec_in_AQ_sel[0:0]),.O(N_64));
defparam desc1223.INIT=8'hCA;
  LUT3 desc1224(.I0(in_A_r[30:30]),.I1(out_r_vec_mult_1[6:6]),.I2(vec_in_AQ_sel[0:0]),.O(N_65));
defparam desc1224.INIT=8'hCA;
  LUT3 desc1225(.I0(in_A_r[26:26]),.I1(out_r_vec_mult_1[2:2]),.I2(vec_in_AQ_sel[0:0]),.O(N_61));
defparam desc1225.INIT=8'hCA;
  LUT3 desc1226(.I0(in_A_r[27:27]),.I1(out_r_vec_mult_1[3:3]),.I2(vec_in_AQ_sel[0:0]),.O(N_62));
defparam desc1226.INIT=8'hCA;
  LUT3 desc1227(.I0(in_A_r[25:25]),.I1(out_r_vec_mult_1[1:1]),.I2(vec_in_AQ_sel[0:0]),.O(N_60));
defparam desc1227.INIT=8'hCA;
  LUT3 desc1228(.I0(in_A_r[31:31]),.I1(out_r_vec_mult_1[7:7]),.I2(vec_in_AQ_sel[0:0]),.O(N_66));
defparam desc1228.INIT=8'hCA;
  LUT3 desc1229(.I0(in_A_r[6:6]),.I1(out_r_vec_mult_3[6:6]),.I2(vec_in_AQ_sel[0:0]),.O(N_41));
defparam desc1229.INIT=8'hCA;
  LUT3 desc1230(.I0(in_A_r[15:15]),.I1(out_r_vec_mult_2[3:3]),.I2(vec_in_AQ_sel[0:0]),.O(N_50));
defparam desc1230.INIT=8'hCA;
  LUT3 desc1231(.I0(in_A_r[4:4]),.I1(out_r_vec_mult_3[4:4]),.I2(vec_in_AQ_sel[0:0]),.O(N_39));
defparam desc1231.INIT=8'hCA;
  LUT3 desc1232(.I0(in_A_r[5:5]),.I1(out_r_vec_mult_3[5:5]),.I2(vec_in_AQ_sel[0:0]),.O(N_40));
defparam desc1232.INIT=8'hCA;
  LUT3 desc1233(.I0(in_A_r[2:2]),.I1(out_r_vec_mult_3[2:2]),.I2(vec_in_AQ_sel[0:0]),.O(N_37));
defparam desc1233.INIT=8'hCA;
  LUT3 desc1234(.I0(in_A_r[3:3]),.I1(out_r_vec_mult_3[3:3]),.I2(vec_in_AQ_sel[0:0]),.O(N_38));
defparam desc1234.INIT=8'hCA;
  LUT3 desc1235(.I0(in_A_i[21:21]),.I1(out_i_vec_mult_2[9:9]),.I2(vec_in_AQ_sel[0:0]),.O(N_156));
defparam desc1235.INIT=8'hCA;
  LUT3 desc1236(.I0(in_A_i[22:22]),.I1(out_i_vec_mult_2[10:10]),.I2(vec_in_AQ_sel[0:0]),.O(N_157));
defparam desc1236.INIT=8'hCA;
  LUT3 desc1237(.I0(in_A_i[20:20]),.I1(out_i_vec_mult_2[8:8]),.I2(vec_in_AQ_sel[0:0]),.O(N_155));
defparam desc1237.INIT=8'hCA;
  LUT3 desc1238(.I0(in_A_i[8:8]),.I1(out_i_vec_mult_3[8:8]),.I2(vec_in_AQ_sel[0:0]),.O(N_143));
defparam desc1238.INIT=8'hCA;
  LUT3 desc1239(.I0(in_A_i[18:18]),.I1(out_i_vec_mult_2[6:6]),.I2(vec_in_AQ_sel[0:0]),.O(N_153));
defparam desc1239.INIT=8'hCA;
  LUT3 desc1240(.I0(in_A_i[19:19]),.I1(out_i_vec_mult_2[7:7]),.I2(vec_in_AQ_sel[0:0]),.O(N_154));
defparam desc1240.INIT=8'hCA;
  LUT3 desc1241(.I0(in_A_i[16:16]),.I1(out_i_vec_mult_2[4:4]),.I2(vec_in_AQ_sel[0:0]),.O(N_151));
defparam desc1241.INIT=8'hCA;
  LUT3 desc1242(.I0(in_A_i[17:17]),.I1(out_i_vec_mult_2[5:5]),.I2(vec_in_AQ_sel[0:0]),.O(N_152));
defparam desc1242.INIT=8'hCA;
  LUT3 desc1243(.I0(in_A_i[14:14]),.I1(out_i_vec_mult_2[2:2]),.I2(vec_in_AQ_sel[0:0]),.O(N_149));
defparam desc1243.INIT=8'hCA;
  LUT3 desc1244(.I0(in_A_i[15:15]),.I1(out_i_vec_mult_2[3:3]),.I2(vec_in_AQ_sel[0:0]),.O(N_150));
defparam desc1244.INIT=8'hCA;
  LUT3 desc1245(.I0(in_A_i[33:33]),.I1(out_i_vec_mult_1[9:9]),.I2(vec_in_AQ_sel[0:0]),.O(N_168));
defparam desc1245.INIT=8'hCA;
  LUT3 desc1246(.I0(in_A_i[34:34]),.I1(out_i_vec_mult_1[10:10]),.I2(vec_in_AQ_sel[0:0]),.O(N_169));
defparam desc1246.INIT=8'hCA;
  LUT3 desc1247(.I0(in_A_i[31:31]),.I1(out_i_vec_mult_1[7:7]),.I2(vec_in_AQ_sel[0:0]),.O(N_166));
defparam desc1247.INIT=8'hCA;
  LUT3 desc1248(.I0(in_A_i[32:32]),.I1(out_i_vec_mult_1[8:8]),.I2(vec_in_AQ_sel[0:0]),.O(N_167));
defparam desc1248.INIT=8'hCA;
  LUT3 desc1249(.I0(in_A_i[30:30]),.I1(out_i_vec_mult_1[6:6]),.I2(vec_in_AQ_sel[0:0]),.O(N_165));
defparam desc1249.INIT=8'hCA;
  LUT3 desc1250(.I0(in_A_i[13:13]),.I1(out_i_vec_mult_2[1:1]),.I2(vec_in_AQ_sel[0:0]),.O(N_148));
defparam desc1250.INIT=8'hCA;
  LUT3 desc1251(.I0(in_A_i[28:28]),.I1(out_i_vec_mult_1[4:4]),.I2(vec_in_AQ_sel[0:0]),.O(N_163));
defparam desc1251.INIT=8'hCA;
  LUT3 desc1252(.I0(in_A_i[29:29]),.I1(out_i_vec_mult_1[5:5]),.I2(vec_in_AQ_sel[0:0]),.O(N_164));
defparam desc1252.INIT=8'hCA;
  LUT3 desc1253(.I0(in_A_i[26:26]),.I1(out_i_vec_mult_1[2:2]),.I2(vec_in_AQ_sel[0:0]),.O(N_161));
defparam desc1253.INIT=8'hCA;
  LUT3 desc1254(.I0(in_A_i[27:27]),.I1(out_i_vec_mult_1[3:3]),.I2(vec_in_AQ_sel[0:0]),.O(N_162));
defparam desc1254.INIT=8'hCA;
  LUT2 N_399_i_lut6_2_o6(.I0(out_inner_prod_i[9:9]),.I1(single_in_R_sel),.O(N_399_i));
defparam N_399_i_lut6_2_o6.INIT=4'h8;
  LUT2 N_399_i_lut6_2_o5(.I0(single_in_R_sel),.I1(out_inner_prod_i[11:11]),.O(N_401_i));
defparam N_399_i_lut6_2_o5.INIT=4'h8;
  LUT2 N_398_i_lut6_2_o6(.I0(out_inner_prod_i[8:8]),.I1(single_in_R_sel),.O(N_398_i));
defparam N_398_i_lut6_2_o6.INIT=4'h8;
  LUT2 N_398_i_lut6_2_o5(.I0(out_inner_prod_i[10:10]),.I1(single_in_R_sel),.O(N_400_i));
defparam N_398_i_lut6_2_o5.INIT=4'h8;
  LUT2 N_395_i_lut6_2_o6(.I0(out_inner_prod_i[5:5]),.I1(single_in_R_sel),.O(N_395_i));
defparam N_395_i_lut6_2_o6.INIT=4'h8;
  LUT2 N_395_i_lut6_2_o5(.I0(out_inner_prod_i[7:7]),.I1(single_in_R_sel),.O(N_397_i));
defparam N_395_i_lut6_2_o5.INIT=4'h8;
  LUT2 N_394_i_lut6_2_o6(.I0(out_inner_prod_i[4:4]),.I1(single_in_R_sel),.O(N_394_i));
defparam N_394_i_lut6_2_o6.INIT=4'h8;
  LUT2 N_394_i_lut6_2_o5(.I0(out_inner_prod_i[6:6]),.I1(single_in_R_sel),.O(N_396_i));
defparam N_394_i_lut6_2_o5.INIT=4'h8;
  LUT2 N_391_i_lut6_2_o6(.I0(out_inner_prod_i[1:1]),.I1(single_in_R_sel),.O(N_391_i));
defparam N_391_i_lut6_2_o6.INIT=4'h8;
  LUT4 N_391_i_lut6_2_o5(.I0(state_0),.I1(state_2),.I2(single_in_R_sel),.I3(done_inv_sqrt),.O(single_in_R_sel_0));
defparam N_391_i_lut6_2_o5.INIT=16'hBAFA;
  LUT2 N_390_i_lut6_2_o6(.I0(out_inner_prod_i[0:0]),.I1(single_in_R_sel),.O(N_390_i));
defparam N_390_i_lut6_2_o6.INIT=4'h8;
  LUT2 N_390_i_lut6_2_o5(.I0(out_inner_prod_i[3:3]),.I1(single_in_R_sel),.O(N_393_i));
defparam N_390_i_lut6_2_o5.INIT=4'h8;
endmodule
module qr_wrapper_inj (out_Q_r,out_Q_i,out_R_i,out_R_r,in_A_r,in_A_i,clk,rst,valid_out,ready,request_out,start,reduced_matrix,p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_,p_desc951_p_O_FDEinv_sqrt_qr_decomp_,p_desc952_p_O_FDEinv_sqrt_qr_decomp_,p_desc953_p_O_FDEinv_sqrt_qr_decomp_,p_desc954_p_O_FDEinv_sqrt_qr_decomp_,p_desc955_p_O_FDEinv_sqrt_qr_decomp_,p_desc956_p_O_FDEinv_sqrt_qr_decomp_,p_desc957_p_O_FDEinv_sqrt_qr_decomp_,p_desc958_p_O_FDEinv_sqrt_qr_decomp_,p_desc959_p_O_FDEinv_sqrt_qr_decomp_,p_desc960_p_O_FDEinv_sqrt_qr_decomp_,p_desc961_p_O_FDEinv_sqrt_qr_decomp_,p_desc962_p_O_FDEinv_sqrt_qr_decomp_,p_desc48_p_O_FDEr_mat_regs_qr_decomp_,p_desc49_p_O_FDEr_mat_regs_qr_decomp_,p_desc50_p_O_FDEr_mat_regs_qr_decomp_,p_desc51_p_O_FDEr_mat_regs_qr_decomp_,p_desc52_p_O_FDEr_mat_regs_qr_decomp_,p_desc53_p_O_FDEr_mat_regs_qr_decomp_,p_desc54_p_O_FDEr_mat_regs_qr_decomp_,p_desc55_p_O_FDEr_mat_regs_qr_decomp_,p_desc56_p_O_FDEr_mat_regs_qr_decomp_,p_desc57_p_O_FDEr_mat_regs_qr_decomp_,p_desc58_p_O_FDEr_mat_regs_qr_decomp_,p_desc59_p_O_FDEr_mat_regs_qr_decomp_,p_desc60_p_O_FDEr_mat_regs_qr_decomp_,p_desc61_p_O_FDEr_mat_regs_qr_decomp_,p_desc62_p_O_FDEr_mat_regs_qr_decomp_,p_desc63_p_O_FDEr_mat_regs_qr_decomp_,p_desc64_p_O_FDEr_mat_regs_qr_decomp_,p_desc65_p_O_FDEr_mat_regs_qr_decomp_,p_desc66_p_O_FDEr_mat_regs_qr_decomp_,p_desc67_p_O_FDEr_mat_regs_qr_decomp_,p_desc68_p_O_FDEr_mat_regs_qr_decomp_,p_desc69_p_O_FDEr_mat_regs_qr_decomp_,p_desc70_p_O_FDEr_mat_regs_qr_decomp_,p_desc71_p_O_FDEr_mat_regs_qr_decomp_,p_desc72_p_O_FDEr_mat_regs_qr_decomp_,p_desc73_p_O_FDEr_mat_regs_qr_decomp_,p_desc74_p_O_FDEr_mat_regs_qr_decomp_,p_desc75_p_O_FDEr_mat_regs_qr_decomp_,p_desc76_p_O_FDEr_mat_regs_qr_decomp_,p_desc77_p_O_FDEr_mat_regs_qr_decomp_,p_desc78_p_O_FDEr_mat_regs_qr_decomp_,p_desc79_p_O_FDEr_mat_regs_qr_decomp_,p_desc80_p_O_FDEr_mat_regs_qr_decomp_,p_desc81_p_O_FDEr_mat_regs_qr_decomp_,p_desc82_p_O_FDEr_mat_regs_qr_decomp_,p_desc83_p_O_FDEr_mat_regs_qr_decomp_,p_desc84_p_O_FDEr_mat_regs_qr_decomp_,p_desc85_p_O_FDEr_mat_regs_qr_decomp_,p_desc86_p_O_FDEr_mat_regs_qr_decomp_,p_desc87_p_O_FDEr_mat_regs_qr_decomp_,p_desc88_p_O_FDEr_mat_regs_qr_decomp_,p_desc89_p_O_FDEr_mat_regs_qr_decomp_,p_desc90_p_O_FDEr_mat_regs_qr_decomp_,p_desc91_p_O_FDEr_mat_regs_qr_decomp_,p_desc92_p_O_FDEr_mat_regs_qr_decomp_,p_desc93_p_O_FDEr_mat_regs_qr_decomp_,p_desc94_p_O_FDEr_mat_regs_qr_decomp_,p_desc95_p_O_FDEr_mat_regs_qr_decomp_,p_desc96_p_O_FDEr_mat_regs_qr_decomp_,p_desc97_p_O_FDEr_mat_regs_qr_decomp_,p_desc98_p_O_FDEr_mat_regs_qr_decomp_,p_desc99_p_O_FDEr_mat_regs_qr_decomp_,p_desc100_p_O_FDEr_mat_regs_qr_decomp_,p_desc101_p_O_FDEr_mat_regs_qr_decomp_,p_desc102_p_O_FDEr_mat_regs_qr_decomp_,p_desc103_p_O_FDEr_mat_regs_qr_decomp_,p_desc104_p_O_FDEr_mat_regs_qr_decomp_,p_desc105_p_O_FDEr_mat_regs_qr_decomp_,p_desc106_p_O_FDEr_mat_regs_qr_decomp_,p_desc107_p_O_FDEr_mat_regs_qr_decomp_,p_desc108_p_O_FDEr_mat_regs_qr_decomp_,p_desc109_p_O_FDEr_mat_regs_qr_decomp_,p_desc110_p_O_FDEr_mat_regs_qr_decomp_,p_desc111_p_O_FDEr_mat_regs_qr_decomp_,p_desc112_p_O_FDEr_mat_regs_qr_decomp_,p_desc113_p_O_FDEr_mat_regs_qr_decomp_,p_desc114_p_O_FDEr_mat_regs_qr_decomp_,p_desc115_p_O_FDEr_mat_regs_qr_decomp_,p_desc116_p_O_FDEr_mat_regs_qr_decomp_,p_desc117_p_O_FDEr_mat_regs_qr_decomp_,p_desc118_p_O_FDEr_mat_regs_qr_decomp_,p_desc119_p_O_FDEr_mat_regs_qr_decomp_,p_desc120_p_O_FDEr_mat_regs_qr_decomp_,p_desc121_p_O_FDEr_mat_regs_qr_decomp_,p_desc122_p_O_FDEr_mat_regs_qr_decomp_,p_desc123_p_O_FDEr_mat_regs_qr_decomp_,p_desc124_p_O_FDEr_mat_regs_qr_decomp_,p_desc125_p_O_FDEr_mat_regs_qr_decomp_,p_desc126_p_O_FDEr_mat_regs_qr_decomp_,p_desc127_p_O_FDEr_mat_regs_qr_decomp_,p_desc128_p_O_FDEr_mat_regs_qr_decomp_,p_desc129_p_O_FDEr_mat_regs_qr_decomp_,p_desc130_p_O_FDEr_mat_regs_qr_decomp_,p_desc131_p_O_FDEr_mat_regs_qr_decomp_,p_desc132_p_O_FDEr_mat_regs_qr_decomp_,p_desc133_p_O_FDEr_mat_regs_qr_decomp_,p_desc134_p_O_FDEr_mat_regs_qr_decomp_,p_desc135_p_O_FDEr_mat_regs_qr_decomp_,p_desc136_p_O_FDEr_mat_regs_qr_decomp_,p_desc137_p_O_FDEr_mat_regs_qr_decomp_,p_desc138_p_O_FDEr_mat_regs_qr_decomp_,p_desc139_p_O_FDEr_mat_regs_qr_decomp_,p_desc140_p_O_FDEr_mat_regs_qr_decomp_,p_desc141_p_O_FDEr_mat_regs_qr_decomp_,p_desc142_p_O_FDEr_mat_regs_qr_decomp_,p_desc143_p_O_FDEr_mat_regs_qr_decomp_,p_desc144_p_O_FDEr_mat_regs_qr_decomp_,p_desc145_p_O_FDEr_mat_regs_qr_decomp_,p_desc146_p_O_FDEr_mat_regs_qr_decomp_,p_desc147_p_O_FDEr_mat_regs_qr_decomp_,p_desc148_p_O_FDEr_mat_regs_qr_decomp_,p_desc149_p_O_FDEr_mat_regs_qr_decomp_,p_desc150_p_O_FDEr_mat_regs_qr_decomp_,p_desc151_p_O_FDEr_mat_regs_qr_decomp_,p_desc152_p_O_FDEr_mat_regs_qr_decomp_,p_desc153_p_O_FDEr_mat_regs_qr_decomp_,p_desc154_p_O_FDEr_mat_regs_qr_decomp_,p_desc155_p_O_FDEr_mat_regs_qr_decomp_,p_desc156_p_O_FDEr_mat_regs_qr_decomp_,p_desc157_p_O_FDEr_mat_regs_qr_decomp_,p_desc158_p_O_FDEr_mat_regs_qr_decomp_,p_desc159_p_O_FDEr_mat_regs_qr_decomp_,p_desc160_p_O_FDEr_mat_regs_qr_decomp_,p_desc161_p_O_FDEr_mat_regs_qr_decomp_,p_desc162_p_O_FDEr_mat_regs_qr_decomp_,p_desc163_p_O_FDEr_mat_regs_qr_decomp_,p_desc164_p_O_FDEr_mat_regs_qr_decomp_,p_desc165_p_O_FDEr_mat_regs_qr_decomp_,p_desc166_p_O_FDEr_mat_regs_qr_decomp_,p_desc167_p_O_FDEr_mat_regs_qr_decomp_,p_desc168_p_O_FDEr_mat_regs_qr_decomp_,p_desc169_p_O_FDEr_mat_regs_qr_decomp_,p_desc170_p_O_FDEr_mat_regs_qr_decomp_,p_desc171_p_O_FDEr_mat_regs_qr_decomp_,p_desc172_p_O_FDEr_mat_regs_qr_decomp_,p_desc173_p_O_FDEr_mat_regs_qr_decomp_,p_desc174_p_O_FDEr_mat_regs_qr_decomp_,p_desc175_p_O_FDEr_mat_regs_qr_decomp_,p_desc176_p_O_FDEr_mat_regs_qr_decomp_,p_desc177_p_O_FDEr_mat_regs_qr_decomp_,p_desc178_p_O_FDEr_mat_regs_qr_decomp_,p_desc179_p_O_FDEr_mat_regs_qr_decomp_,p_desc180_p_O_FDEr_mat_regs_qr_decomp_,p_desc181_p_O_FDEr_mat_regs_qr_decomp_,p_desc182_p_O_FDEr_mat_regs_qr_decomp_,p_desc183_p_O_FDEr_mat_regs_qr_decomp_,p_desc184_p_O_FDEr_mat_regs_qr_decomp_,p_desc185_p_O_FDEr_mat_regs_qr_decomp_,p_desc186_p_O_FDEr_mat_regs_qr_decomp_,p_desc187_p_O_FDEr_mat_regs_qr_decomp_,p_desc188_p_O_FDEr_mat_regs_qr_decomp_,p_desc189_p_O_FDEr_mat_regs_qr_decomp_,p_desc190_p_O_FDEr_mat_regs_qr_decomp_,p_desc191_p_O_FDEr_mat_regs_qr_decomp_,p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_,p_desc739_p_O_FDEvec_sub_qr_decomp_,p_desc740_p_O_FDEvec_sub_qr_decomp_,p_desc741_p_O_FDEvec_sub_qr_decomp_,p_desc742_p_O_FDEvec_sub_qr_decomp_,p_desc743_p_O_FDEvec_sub_qr_decomp_,p_desc744_p_O_FDEvec_sub_qr_decomp_,p_desc745_p_O_FDEvec_sub_qr_decomp_,p_desc746_p_O_FDEvec_sub_qr_decomp_,p_desc747_p_O_FDEvec_sub_qr_decomp_,p_desc748_p_O_FDEvec_sub_qr_decomp_,p_desc749_p_O_FDEvec_sub_qr_decomp_,p_desc750_p_O_FDEvec_sub_qr_decomp_,p_desc751_p_O_FDEvec_sub_qr_decomp_,p_desc752_p_O_FDEvec_sub_qr_decomp_,p_desc753_p_O_FDEvec_sub_qr_decomp_,p_desc754_p_O_FDEvec_sub_qr_decomp_,p_desc755_p_O_FDEvec_sub_qr_decomp_,p_desc756_p_O_FDEvec_sub_qr_decomp_,p_desc757_p_O_FDEvec_sub_qr_decomp_,p_desc758_p_O_FDEvec_sub_qr_decomp_,p_desc759_p_O_FDEvec_sub_qr_decomp_,p_desc760_p_O_FDEvec_sub_qr_decomp_,p_desc761_p_O_FDEvec_sub_qr_decomp_,p_desc762_p_O_FDEvec_sub_qr_decomp_,p_desc763_p_O_FDEvec_sub_qr_decomp_,p_desc764_p_O_FDEvec_sub_qr_decomp_,p_desc765_p_O_FDEvec_sub_qr_decomp_,p_desc766_p_O_FDEvec_sub_qr_decomp_,p_desc767_p_O_FDEvec_sub_qr_decomp_,p_desc768_p_O_FDEvec_sub_qr_decomp_,p_desc769_p_O_FDEvec_sub_qr_decomp_,p_desc770_p_O_FDEvec_sub_qr_decomp_,p_desc771_p_O_FDEvec_sub_qr_decomp_,p_desc772_p_O_FDEvec_sub_qr_decomp_,p_desc773_p_O_FDEvec_sub_qr_decomp_,p_desc774_p_O_FDEvec_sub_qr_decomp_,p_desc775_p_O_FDEvec_sub_qr_decomp_,p_desc776_p_O_FDEvec_sub_qr_decomp_,p_desc777_p_O_FDEvec_sub_qr_decomp_,p_desc778_p_O_FDEvec_sub_qr_decomp_,p_desc779_p_O_FDEvec_sub_qr_decomp_,p_desc780_p_O_FDEvec_sub_qr_decomp_,p_desc781_p_O_FDEvec_sub_qr_decomp_,p_desc782_p_O_FDEvec_sub_qr_decomp_,p_desc783_p_O_FDEvec_sub_qr_decomp_,p_desc784_p_O_FDEvec_sub_qr_decomp_,p_desc785_p_O_FDEvec_sub_qr_decomp_,p_desc786_p_O_FDEvec_sub_qr_decomp_,p_desc787_p_O_FDEvec_sub_qr_decomp_,p_desc788_p_O_FDEvec_sub_qr_decomp_,p_desc789_p_O_FDEvec_sub_qr_decomp_,p_desc790_p_O_FDEvec_sub_qr_decomp_,p_desc791_p_O_FDEvec_sub_qr_decomp_,p_desc792_p_O_FDEvec_sub_qr_decomp_,p_desc793_p_O_FDEvec_sub_qr_decomp_,p_desc794_p_O_FDEvec_sub_qr_decomp_,p_desc795_p_O_FDEvec_sub_qr_decomp_,p_desc796_p_O_FDEvec_sub_qr_decomp_,p_desc797_p_O_FDEvec_sub_qr_decomp_,p_desc798_p_O_FDEvec_sub_qr_decomp_,p_desc799_p_O_FDEvec_sub_qr_decomp_,p_desc800_p_O_FDEvec_sub_qr_decomp_,p_desc801_p_O_FDEvec_sub_qr_decomp_,p_desc802_p_O_FDEvec_sub_qr_decomp_,p_desc803_p_O_FDEvec_sub_qr_decomp_,p_desc804_p_O_FDEvec_sub_qr_decomp_,p_desc805_p_O_FDEvec_sub_qr_decomp_,p_desc806_p_O_FDEvec_sub_qr_decomp_,p_desc807_p_O_FDEvec_sub_qr_decomp_,p_desc808_p_O_FDEvec_sub_qr_decomp_,p_desc809_p_O_FDEvec_sub_qr_decomp_,p_desc810_p_O_FDEvec_sub_qr_decomp_,p_desc811_p_O_FDEvec_sub_qr_decomp_,p_desc812_p_O_FDEvec_sub_qr_decomp_,p_desc813_p_O_FDEvec_sub_qr_decomp_,p_desc814_p_O_FDEvec_sub_qr_decomp_,p_desc815_p_O_FDEvec_sub_qr_decomp_,p_desc816_p_O_FDEvec_sub_qr_decomp_,p_desc817_p_O_FDEvec_sub_qr_decomp_,p_desc818_p_O_FDEvec_sub_qr_decomp_,p_desc819_p_O_FDEvec_sub_qr_decomp_,p_desc820_p_O_FDEvec_sub_qr_decomp_,p_desc821_p_O_FDEvec_sub_qr_decomp_,p_desc822_p_O_FDEvec_sub_qr_decomp_,p_desc823_p_O_FDEvec_sub_qr_decomp_,p_desc824_p_O_FDEvec_sub_qr_decomp_,p_desc825_p_O_FDEvec_sub_qr_decomp_,p_desc826_p_O_FDEvec_sub_qr_decomp_,p_desc827_p_O_FDEvec_sub_qr_decomp_,p_desc828_p_O_FDEvec_sub_qr_decomp_,p_desc829_p_O_FDEvec_sub_qr_decomp_,p_desc830_p_O_FDEvec_sub_qr_decomp_,p_desc831_p_O_FDEvec_sub_qr_decomp_,p_desc832_p_O_FDEvec_sub_qr_decomp_,p_desc833_p_O_FDEvec_sub_qr_decomp_,p_desc834_p_O_FDEvec_sub_qr_decomp_,p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_,p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_,p_desc318_p_O_FDCinner_prod_qr_decomp_,p_desc319_p_O_FDCinner_prod_qr_decomp_,p_desc320_p_O_FDCinner_prod_qr_decomp_,p_desc321_p_O_FDCinner_prod_qr_decomp_,p_desc322_p_O_FDCinner_prod_qr_decomp_,p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_,p_done_Z_p_O_FDCinner_prod_qr_decomp_,p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_,p_desc325_p_O_FDCinner_prod_qr_decomp_,p_desc326_p_O_FDCinner_prod_qr_decomp_,p_desc327_p_O_FDCinner_prod_qr_decomp_,p_desc328_p_O_FDCinner_prod_qr_decomp_,p_desc329_p_O_FDCinner_prod_qr_decomp_,p_desc330_p_O_FDCinner_prod_qr_decomp_,p_desc331_p_O_FDCinner_prod_qr_decomp_,p_desc332_p_O_FDCinner_prod_qr_decomp_,p_desc333_p_O_FDCinner_prod_qr_decomp_,p_desc334_p_O_FDCinner_prod_qr_decomp_,p_desc335_p_O_FDCinner_prod_qr_decomp_,p_desc336_p_O_FDCinner_prod_qr_decomp_,p_desc337_p_O_FDCinner_prod_qr_decomp_,p_desc338_p_O_FDCinner_prod_qr_decomp_,p_desc339_p_O_FDCinner_prod_qr_decomp_,p_desc340_p_O_FDCinner_prod_qr_decomp_,p_desc341_p_O_FDCinner_prod_qr_decomp_,p_desc342_p_O_FDCinner_prod_qr_decomp_,p_desc343_p_O_FDCinner_prod_qr_decomp_,p_desc344_p_O_FDCinner_prod_qr_decomp_,p_desc345_p_O_FDCinner_prod_qr_decomp_,p_desc346_p_O_FDCinner_prod_qr_decomp_,p_desc347_p_O_FDCinner_prod_qr_decomp_,p_desc348_p_O_FDCinner_prod_qr_decomp_,p_desc349_p_O_FDCinner_prod_qr_decomp_,p_desc350_p_O_FDCinner_prod_qr_decomp_,p_desc375_p_O_FDCinner_prod_qr_decomp_,p_desc376_p_O_FDCinner_prod_qr_decomp_,p_desc377_p_O_FDCinner_prod_qr_decomp_,p_desc378_p_O_FDCinner_prod_qr_decomp_,p_desc379_p_O_FDCinner_prod_qr_decomp_,p_desc380_p_O_FDCinner_prod_qr_decomp_,p_desc381_p_O_FDCinner_prod_qr_decomp_,p_desc382_p_O_FDCinner_prod_qr_decomp_,p_desc383_p_O_FDCinner_prod_qr_decomp_,p_desc384_p_O_FDCinner_prod_qr_decomp_,p_desc385_p_O_FDCinner_prod_qr_decomp_,p_desc386_p_O_FDCinner_prod_qr_decomp_,p_desc387_p_O_FDCinner_prod_qr_decomp_,p_desc388_p_O_FDCinner_prod_qr_decomp_,p_desc389_p_O_FDCinner_prod_qr_decomp_,p_desc390_p_O_FDCinner_prod_qr_decomp_,p_desc391_p_O_FDCinner_prod_qr_decomp_,p_desc392_p_O_FDCinner_prod_qr_decomp_,p_desc393_p_O_FDCinner_prod_qr_decomp_,p_desc394_p_O_FDCinner_prod_qr_decomp_,p_desc395_p_O_FDCinner_prod_qr_decomp_,p_desc396_p_O_FDCinner_prod_qr_decomp_,p_desc397_p_O_FDCinner_prod_qr_decomp_,p_desc398_p_O_FDCinner_prod_qr_decomp_,p_done_Z_p_O_FDCinv_sqrt_qr_decomp_,p_desc946_p_O_FDCinv_sqrt_qr_decomp_,p_desc947_p_O_FDCinv_sqrt_qr_decomp_,p_desc948_p_O_FDCinv_sqrt_qr_decomp_,p_desc949_p_O_FDCinv_sqrt_qr_decomp_,p_desc950_p_O_FDCinv_sqrt_qr_decomp_,p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_,p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_,p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_,p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_,p_start_QR_Z_p_O_FDC,p_wr_A_QR_Z_p_O_FDC,p_valid_out_Z_p_O_FDC,p_ready_Z_p_O_FDC,p_red_mat_reg_Z_p_O_FDC,p_desc1317_p_O_FDC,p_desc1318_p_O_FDC,p_desc1319_p_O_FDC,p_desc1320_p_O_FDC,p_desc1321_p_O_FDC,p_desc1322_p_O_FDC,p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_,p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_,p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_,p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_,p_desc324_p_O_FDCEinner_prod_qr_decomp_,p_desc351_p_O_FDCEinner_prod_qr_decomp_,p_desc352_p_O_FDCEinner_prod_qr_decomp_,p_desc353_p_O_FDCEinner_prod_qr_decomp_,p_desc354_p_O_FDCEinner_prod_qr_decomp_,p_desc355_p_O_FDCEinner_prod_qr_decomp_,p_desc356_p_O_FDCEinner_prod_qr_decomp_,p_desc357_p_O_FDCEinner_prod_qr_decomp_,p_desc358_p_O_FDCEinner_prod_qr_decomp_,p_desc359_p_O_FDCEinner_prod_qr_decomp_,p_desc360_p_O_FDCEinner_prod_qr_decomp_,p_desc361_p_O_FDCEinner_prod_qr_decomp_,p_desc362_p_O_FDCEinner_prod_qr_decomp_,p_desc363_p_O_FDCEinner_prod_qr_decomp_,p_desc364_p_O_FDCEinner_prod_qr_decomp_,p_desc365_p_O_FDCEinner_prod_qr_decomp_,p_desc366_p_O_FDCEinner_prod_qr_decomp_,p_desc367_p_O_FDCEinner_prod_qr_decomp_,p_desc368_p_O_FDCEinner_prod_qr_decomp_,p_desc369_p_O_FDCEinner_prod_qr_decomp_,p_desc370_p_O_FDCEinner_prod_qr_decomp_,p_desc371_p_O_FDCEinner_prod_qr_decomp_,p_desc372_p_O_FDCEinner_prod_qr_decomp_,p_desc373_p_O_FDCEinner_prod_qr_decomp_,p_desc374_p_O_FDCEinner_prod_qr_decomp_,p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_,p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_);
output [47:0] out_Q_r ;
output [47:0] out_Q_i ;
output [47:12] out_R_i ;
output [47:0] out_R_r ;
input [47:0] in_A_r ;
input [47:0] in_A_i ;
input clk ;
input rst ;
output valid_out ;
output ready ;
input request_out ;
input start ;
input reduced_matrix ;
wire clk ;
wire rst ;
wire valid_out ;
wire ready ;
wire request_out ;
wire start ;
wire reduced_matrix ;
wire [1:0] col_sel_AQ ;
wire [1:0] col_sel_AQ_4 ;
wire [1:0] col_sel_R ;
wire [1:0] state ;
wire [1:0] state_ns ;
wire start_QR ;
wire start_QR_0 ;
wire wr_A_QR ;
wire wr_A_QR_0 ;
wire valid_out_0 ;
wire ready_0 ;
wire red_mat_reg ;
wire red_mat_reg_0 ;
wire N_14_i ;
wire N_16_i ;
wire N_26 ;
wire done_QR ;
wire N_50 ;
wire N_49 ;
wire N_48 ;
wire N_47 ;
wire GND ;
wire VCC ;
input p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_ ;
input p_desc951_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc952_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc953_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc954_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc955_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc956_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc957_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc958_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc959_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc960_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc961_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc962_p_O_FDEinv_sqrt_qr_decomp_ ;
input p_desc48_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc49_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc50_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc51_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc52_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc53_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc54_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc55_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc56_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc57_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc58_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc59_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc60_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc61_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc62_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc63_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc64_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc65_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc66_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc67_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc68_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc69_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc70_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc71_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc72_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc73_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc74_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc75_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc76_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc77_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc78_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc79_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc80_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc81_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc82_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc83_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc84_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc85_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc86_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc87_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc88_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc89_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc90_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc91_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc92_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc93_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc94_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc95_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc96_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc97_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc98_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc99_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc100_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc101_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc102_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc103_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc104_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc105_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc106_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc107_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc108_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc109_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc110_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc111_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc112_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc113_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc114_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc115_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc116_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc117_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc118_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc119_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc120_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc121_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc122_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc123_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc124_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc125_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc126_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc127_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc128_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc129_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc130_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc131_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc132_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc133_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc134_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc135_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc136_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc137_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc138_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc139_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc140_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc141_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc142_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc143_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc144_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc145_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc146_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc147_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc148_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc149_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc150_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc151_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc152_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc153_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc154_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc155_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc156_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc157_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc158_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc159_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc160_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc161_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc162_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc163_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc164_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc165_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc166_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc167_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc168_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc169_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc170_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc171_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc172_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc173_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc174_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc175_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc176_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc177_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc178_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc179_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc180_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc181_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc182_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc183_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc184_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc185_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc186_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc187_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc188_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc189_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc190_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_desc191_p_O_FDEr_mat_regs_qr_decomp_ ;
input p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_ ;
input p_desc739_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc740_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc741_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc742_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc743_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc744_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc745_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc746_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc747_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc748_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc749_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc750_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc751_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc752_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc753_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc754_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc755_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc756_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc757_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc758_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc759_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc760_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc761_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc762_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc763_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc764_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc765_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc766_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc767_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc768_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc769_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc770_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc771_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc772_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc773_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc774_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc775_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc776_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc777_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc778_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc779_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc780_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc781_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc782_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc783_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc784_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc785_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc786_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc787_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc788_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc789_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc790_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc791_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc792_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc793_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc794_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc795_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc796_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc797_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc798_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc799_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc800_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc801_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc802_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc803_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc804_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc805_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc806_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc807_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc808_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc809_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc810_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc811_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc812_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc813_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc814_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc815_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc816_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc817_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc818_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc819_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc820_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc821_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc822_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc823_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc824_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc825_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc826_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc827_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc828_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc829_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc830_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc831_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc832_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc833_p_O_FDEvec_sub_qr_decomp_ ;
input p_desc834_p_O_FDEvec_sub_qr_decomp_ ;
input p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_ ;
input p_desc318_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc319_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc320_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc321_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc322_p_O_FDCinner_prod_qr_decomp_ ;
input p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_ ;
input p_done_Z_p_O_FDCinner_prod_qr_decomp_ ;
input p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc325_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc326_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc327_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc328_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc329_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc330_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc331_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc332_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc333_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc334_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc335_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc336_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc337_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc338_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc339_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc340_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc341_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc342_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc343_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc344_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc345_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc346_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc347_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc348_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc349_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc350_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc375_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc376_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc377_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc378_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc379_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc380_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc381_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc382_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc383_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc384_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc385_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc386_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc387_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc388_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc389_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc390_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc391_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc392_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc393_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc394_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc395_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc396_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc397_p_O_FDCinner_prod_qr_decomp_ ;
input p_desc398_p_O_FDCinner_prod_qr_decomp_ ;
input p_done_Z_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc946_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc947_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc948_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc949_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc950_p_O_FDCinv_sqrt_qr_decomp_ ;
input p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_ ;
input p_start_QR_Z_p_O_FDC ;
input p_wr_A_QR_Z_p_O_FDC ;
input p_valid_out_Z_p_O_FDC ;
input p_ready_Z_p_O_FDC ;
input p_red_mat_reg_Z_p_O_FDC ;
input p_desc1317_p_O_FDC ;
input p_desc1318_p_O_FDC ;
input p_desc1319_p_O_FDC ;
input p_desc1320_p_O_FDC ;
input p_desc1321_p_O_FDC ;
input p_desc1322_p_O_FDC ;
input p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_ ;
input p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_ ;
input p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_ ;
input p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_ ;
input p_desc324_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc351_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc352_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc353_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc354_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc355_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc356_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc357_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc358_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc359_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc360_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc361_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc362_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc363_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc364_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc365_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc366_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc367_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc368_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc369_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc370_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc371_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc372_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc373_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc374_p_O_FDCEinner_prod_qr_decomp_ ;
input p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
input p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_ ;
// instances
  p_O_FDC start_QR_Z(.Q(start_QR),.D(start_QR_0),.C(clk),.CLR(rst),.E(p_start_QR_Z_p_O_FDC));
  p_O_FDC wr_A_QR_Z(.Q(wr_A_QR),.D(wr_A_QR_0),.C(clk),.CLR(rst),.E(p_wr_A_QR_Z_p_O_FDC));
  p_O_FDC valid_out_Z(.Q(valid_out),.D(valid_out_0),.C(clk),.CLR(rst),.E(p_valid_out_Z_p_O_FDC));
  p_O_FDC ready_Z(.Q(ready),.D(ready_0),.C(clk),.CLR(rst),.E(p_ready_Z_p_O_FDC));
  p_O_FDC red_mat_reg_Z(.Q(red_mat_reg),.D(red_mat_reg_0),.C(clk),.CLR(rst),.E(p_red_mat_reg_Z_p_O_FDC));
  p_O_FDC desc1317(.Q(col_sel_AQ[1:1]),.D(col_sel_AQ_4[1:1]),.C(clk),.CLR(rst),.E(p_desc1317_p_O_FDC));
  p_O_FDC desc1318(.Q(col_sel_R[0:0]),.D(N_14_i),.C(clk),.CLR(rst),.E(p_desc1318_p_O_FDC));
  p_O_FDC desc1319(.Q(col_sel_R[1:1]),.D(N_16_i),.C(clk),.CLR(rst),.E(p_desc1319_p_O_FDC));
  p_O_FDC desc1320(.Q(col_sel_AQ[0:0]),.D(col_sel_AQ_4[0:0]),.C(clk),.CLR(rst),.E(p_desc1320_p_O_FDC));
  p_O_FDC desc1321(.Q(state[0:0]),.D(state_ns[0:0]),.C(clk),.CLR(rst),.E(p_desc1321_p_O_FDC));
  p_O_FDC desc1322(.Q(state[1:1]),.D(state_ns[1:1]),.C(clk),.CLR(rst),.E(p_desc1322_p_O_FDC));
  LUT6_L desc1323(.I0(request_out),.I1(start),.I2(col_sel_AQ[1:1]),.I3(col_sel_AQ[0:0]),.I4(state[0:0]),.I5(state[1:1]),.LO(col_sel_AQ_4[1:1]));
defparam desc1323.INIT=64'h0FF0F0F00FF01010;
  LUT6_L start_QR_e(.I0(red_mat_reg),.I1(col_sel_AQ[1:1]),.I2(col_sel_AQ[0:0]),.I3(start_QR),.I4(state[0:0]),.I5(state[1:1]),.LO(start_QR_0));
defparam start_QR_e.INIT=64'hFF000000FFE0FF00;
  LUT3 desc1324(.I0(red_mat_reg),.I1(col_sel_AQ[1:1]),.I2(col_sel_AQ[0:0]),.O(N_26));
defparam desc1324.INIT=8'h1F;
  LUT5_L ready_e(.I0(request_out),.I1(start),.I2(ready),.I3(state[0:0]),.I4(state[1:1]),.LO(ready_0));
defparam ready_e.INIT=32'hF0F0F011;
  LUT5_L red_mat_reg_e(.I0(reduced_matrix),.I1(start),.I2(red_mat_reg),.I3(state[0:0]),.I4(state[1:1]),.LO(red_mat_reg_0));
defparam red_mat_reg_e.INIT=32'hF0F0F0B8;
  LUT5_L desc1325(.I0(request_out),.I1(start),.I2(state[0:0]),.I3(state[1:1]),.I4(N_26),.LO(state_ns[0:0]));
defparam desc1325.INIT=32'hF0FE000E;
  LUT5_L desc1326(.I0(request_out),.I1(start),.I2(col_sel_AQ[0:0]),.I3(state[0:0]),.I4(state[1:1]),.LO(col_sel_AQ_4[0:0]));
defparam desc1326.INIT=32'h0FF00F10;
  LUT6_L desc1327(.I0(request_out),.I1(start),.I2(state[0:0]),.I3(state[1:1]),.I4(col_sel_R[0:0]),.I5(col_sel_R[1:1]),.LO(N_16_i));
defparam desc1327.INIT=64'h0FFDFFFDF0000000;
  LUT5_L desc1328(.I0(request_out),.I1(start),.I2(state[0:0]),.I3(state[1:1]),.I4(col_sel_R[0:0]),.LO(N_14_i));
defparam desc1328.INIT=32'h0FFDF000;
  LUT6_L valid_out_e(.I0(request_out),.I1(start),.I2(valid_out),.I3(state[0:0]),.I4(state[1:1]),.I5(N_26),.LO(valid_out_0));
defparam valid_out_e.INIT=64'hF0F0F0F200F0F0F2;
  LUT6_L desc1329(.I0(request_out),.I1(start),.I2(done_QR),.I3(state[0:0]),.I4(state[1:1]),.I5(N_26),.LO(state_ns[1:1]));
defparam desc1329.INIT=64'hFF0F0022000FFF22;
  LUT5_L wr_A_QR_e(.I0(start),.I1(wr_A_QR),.I2(state[0:0]),.I3(state[1:1]),.I4(N_26),.LO(wr_A_QR_0));
defparam wr_A_QR_e.INIT=32'hCCCECC0E;
  qr_decomp_inj qr_decomp_inst(.out_Q_r(out_Q_r[47:0]),.out_Q_i(out_Q_i[47:0]),.col_sel_R(col_sel_R[1:0]),.out_R_i(out_R_i[47:12]),.out_R_r(out_R_r[47:0]),.col_sel_AQ(col_sel_AQ[1:0]),.in_A_r(in_A_r[47:0]),.in_A_i(in_A_i[47:0]),.clk(clk),.rst(rst),.wr_A_QR(wr_A_QR),.start_QR(start_QR),.done_QR(done_QR),.red_mat_reg_0(red_mat_reg),.p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_(p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_(p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_(p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_),.p_desc951_p_O_FDEinv_sqrt_(p_desc951_p_O_FDEinv_sqrt_qr_decomp_),.p_desc952_p_O_FDEinv_sqrt_(p_desc952_p_O_FDEinv_sqrt_qr_decomp_),.p_desc953_p_O_FDEinv_sqrt_(p_desc953_p_O_FDEinv_sqrt_qr_decomp_),.p_desc954_p_O_FDEinv_sqrt_(p_desc954_p_O_FDEinv_sqrt_qr_decomp_),.p_desc955_p_O_FDEinv_sqrt_(p_desc955_p_O_FDEinv_sqrt_qr_decomp_),.p_desc956_p_O_FDEinv_sqrt_(p_desc956_p_O_FDEinv_sqrt_qr_decomp_),.p_desc957_p_O_FDEinv_sqrt_(p_desc957_p_O_FDEinv_sqrt_qr_decomp_),.p_desc958_p_O_FDEinv_sqrt_(p_desc958_p_O_FDEinv_sqrt_qr_decomp_),.p_desc959_p_O_FDEinv_sqrt_(p_desc959_p_O_FDEinv_sqrt_qr_decomp_),.p_desc960_p_O_FDEinv_sqrt_(p_desc960_p_O_FDEinv_sqrt_qr_decomp_),.p_desc961_p_O_FDEinv_sqrt_(p_desc961_p_O_FDEinv_sqrt_qr_decomp_),.p_desc962_p_O_FDEinv_sqrt_(p_desc962_p_O_FDEinv_sqrt_qr_decomp_),.p_desc48_p_O_FDEr_mat_regs_(p_desc48_p_O_FDEr_mat_regs_qr_decomp_),.p_desc49_p_O_FDEr_mat_regs_(p_desc49_p_O_FDEr_mat_regs_qr_decomp_),.p_desc50_p_O_FDEr_mat_regs_(p_desc50_p_O_FDEr_mat_regs_qr_decomp_),.p_desc51_p_O_FDEr_mat_regs_(p_desc51_p_O_FDEr_mat_regs_qr_decomp_),.p_desc52_p_O_FDEr_mat_regs_(p_desc52_p_O_FDEr_mat_regs_qr_decomp_),.p_desc53_p_O_FDEr_mat_regs_(p_desc53_p_O_FDEr_mat_regs_qr_decomp_),.p_desc54_p_O_FDEr_mat_regs_(p_desc54_p_O_FDEr_mat_regs_qr_decomp_),.p_desc55_p_O_FDEr_mat_regs_(p_desc55_p_O_FDEr_mat_regs_qr_decomp_),.p_desc56_p_O_FDEr_mat_regs_(p_desc56_p_O_FDEr_mat_regs_qr_decomp_),.p_desc57_p_O_FDEr_mat_regs_(p_desc57_p_O_FDEr_mat_regs_qr_decomp_),.p_desc58_p_O_FDEr_mat_regs_(p_desc58_p_O_FDEr_mat_regs_qr_decomp_),.p_desc59_p_O_FDEr_mat_regs_(p_desc59_p_O_FDEr_mat_regs_qr_decomp_),.p_desc60_p_O_FDEr_mat_regs_(p_desc60_p_O_FDEr_mat_regs_qr_decomp_),.p_desc61_p_O_FDEr_mat_regs_(p_desc61_p_O_FDEr_mat_regs_qr_decomp_),.p_desc62_p_O_FDEr_mat_regs_(p_desc62_p_O_FDEr_mat_regs_qr_decomp_),.p_desc63_p_O_FDEr_mat_regs_(p_desc63_p_O_FDEr_mat_regs_qr_decomp_),.p_desc64_p_O_FDEr_mat_regs_(p_desc64_p_O_FDEr_mat_regs_qr_decomp_),.p_desc65_p_O_FDEr_mat_regs_(p_desc65_p_O_FDEr_mat_regs_qr_decomp_),.p_desc66_p_O_FDEr_mat_regs_(p_desc66_p_O_FDEr_mat_regs_qr_decomp_),.p_desc67_p_O_FDEr_mat_regs_(p_desc67_p_O_FDEr_mat_regs_qr_decomp_),.p_desc68_p_O_FDEr_mat_regs_(p_desc68_p_O_FDEr_mat_regs_qr_decomp_),.p_desc69_p_O_FDEr_mat_regs_(p_desc69_p_O_FDEr_mat_regs_qr_decomp_),.p_desc70_p_O_FDEr_mat_regs_(p_desc70_p_O_FDEr_mat_regs_qr_decomp_),.p_desc71_p_O_FDEr_mat_regs_(p_desc71_p_O_FDEr_mat_regs_qr_decomp_),.p_desc72_p_O_FDEr_mat_regs_(p_desc72_p_O_FDEr_mat_regs_qr_decomp_),.p_desc73_p_O_FDEr_mat_regs_(p_desc73_p_O_FDEr_mat_regs_qr_decomp_),.p_desc74_p_O_FDEr_mat_regs_(p_desc74_p_O_FDEr_mat_regs_qr_decomp_),.p_desc75_p_O_FDEr_mat_regs_(p_desc75_p_O_FDEr_mat_regs_qr_decomp_),.p_desc76_p_O_FDEr_mat_regs_(p_desc76_p_O_FDEr_mat_regs_qr_decomp_),.p_desc77_p_O_FDEr_mat_regs_(p_desc77_p_O_FDEr_mat_regs_qr_decomp_),.p_desc78_p_O_FDEr_mat_regs_(p_desc78_p_O_FDEr_mat_regs_qr_decomp_),.p_desc79_p_O_FDEr_mat_regs_(p_desc79_p_O_FDEr_mat_regs_qr_decomp_),.p_desc80_p_O_FDEr_mat_regs_(p_desc80_p_O_FDEr_mat_regs_qr_decomp_),.p_desc81_p_O_FDEr_mat_regs_(p_desc81_p_O_FDEr_mat_regs_qr_decomp_),.p_desc82_p_O_FDEr_mat_regs_(p_desc82_p_O_FDEr_mat_regs_qr_decomp_),.p_desc83_p_O_FDEr_mat_regs_(p_desc83_p_O_FDEr_mat_regs_qr_decomp_),.p_desc84_p_O_FDEr_mat_regs_(p_desc84_p_O_FDEr_mat_regs_qr_decomp_),.p_desc85_p_O_FDEr_mat_regs_(p_desc85_p_O_FDEr_mat_regs_qr_decomp_),.p_desc86_p_O_FDEr_mat_regs_(p_desc86_p_O_FDEr_mat_regs_qr_decomp_),.p_desc87_p_O_FDEr_mat_regs_(p_desc87_p_O_FDEr_mat_regs_qr_decomp_),.p_desc88_p_O_FDEr_mat_regs_(p_desc88_p_O_FDEr_mat_regs_qr_decomp_),.p_desc89_p_O_FDEr_mat_regs_(p_desc89_p_O_FDEr_mat_regs_qr_decomp_),.p_desc90_p_O_FDEr_mat_regs_(p_desc90_p_O_FDEr_mat_regs_qr_decomp_),.p_desc91_p_O_FDEr_mat_regs_(p_desc91_p_O_FDEr_mat_regs_qr_decomp_),.p_desc92_p_O_FDEr_mat_regs_(p_desc92_p_O_FDEr_mat_regs_qr_decomp_),.p_desc93_p_O_FDEr_mat_regs_(p_desc93_p_O_FDEr_mat_regs_qr_decomp_),.p_desc94_p_O_FDEr_mat_regs_(p_desc94_p_O_FDEr_mat_regs_qr_decomp_),.p_desc95_p_O_FDEr_mat_regs_(p_desc95_p_O_FDEr_mat_regs_qr_decomp_),.p_desc96_p_O_FDEr_mat_regs_(p_desc96_p_O_FDEr_mat_regs_qr_decomp_),.p_desc97_p_O_FDEr_mat_regs_(p_desc97_p_O_FDEr_mat_regs_qr_decomp_),.p_desc98_p_O_FDEr_mat_regs_(p_desc98_p_O_FDEr_mat_regs_qr_decomp_),.p_desc99_p_O_FDEr_mat_regs_(p_desc99_p_O_FDEr_mat_regs_qr_decomp_),.p_desc100_p_O_FDEr_mat_regs_(p_desc100_p_O_FDEr_mat_regs_qr_decomp_),.p_desc101_p_O_FDEr_mat_regs_(p_desc101_p_O_FDEr_mat_regs_qr_decomp_),.p_desc102_p_O_FDEr_mat_regs_(p_desc102_p_O_FDEr_mat_regs_qr_decomp_),.p_desc103_p_O_FDEr_mat_regs_(p_desc103_p_O_FDEr_mat_regs_qr_decomp_),.p_desc104_p_O_FDEr_mat_regs_(p_desc104_p_O_FDEr_mat_regs_qr_decomp_),.p_desc105_p_O_FDEr_mat_regs_(p_desc105_p_O_FDEr_mat_regs_qr_decomp_),.p_desc106_p_O_FDEr_mat_regs_(p_desc106_p_O_FDEr_mat_regs_qr_decomp_),.p_desc107_p_O_FDEr_mat_regs_(p_desc107_p_O_FDEr_mat_regs_qr_decomp_),.p_desc108_p_O_FDEr_mat_regs_(p_desc108_p_O_FDEr_mat_regs_qr_decomp_),.p_desc109_p_O_FDEr_mat_regs_(p_desc109_p_O_FDEr_mat_regs_qr_decomp_),.p_desc110_p_O_FDEr_mat_regs_(p_desc110_p_O_FDEr_mat_regs_qr_decomp_),.p_desc111_p_O_FDEr_mat_regs_(p_desc111_p_O_FDEr_mat_regs_qr_decomp_),.p_desc112_p_O_FDEr_mat_regs_(p_desc112_p_O_FDEr_mat_regs_qr_decomp_),.p_desc113_p_O_FDEr_mat_regs_(p_desc113_p_O_FDEr_mat_regs_qr_decomp_),.p_desc114_p_O_FDEr_mat_regs_(p_desc114_p_O_FDEr_mat_regs_qr_decomp_),.p_desc115_p_O_FDEr_mat_regs_(p_desc115_p_O_FDEr_mat_regs_qr_decomp_),.p_desc116_p_O_FDEr_mat_regs_(p_desc116_p_O_FDEr_mat_regs_qr_decomp_),.p_desc117_p_O_FDEr_mat_regs_(p_desc117_p_O_FDEr_mat_regs_qr_decomp_),.p_desc118_p_O_FDEr_mat_regs_(p_desc118_p_O_FDEr_mat_regs_qr_decomp_),.p_desc119_p_O_FDEr_mat_regs_(p_desc119_p_O_FDEr_mat_regs_qr_decomp_),.p_desc120_p_O_FDEr_mat_regs_(p_desc120_p_O_FDEr_mat_regs_qr_decomp_),.p_desc121_p_O_FDEr_mat_regs_(p_desc121_p_O_FDEr_mat_regs_qr_decomp_),.p_desc122_p_O_FDEr_mat_regs_(p_desc122_p_O_FDEr_mat_regs_qr_decomp_),.p_desc123_p_O_FDEr_mat_regs_(p_desc123_p_O_FDEr_mat_regs_qr_decomp_),.p_desc124_p_O_FDEr_mat_regs_(p_desc124_p_O_FDEr_mat_regs_qr_decomp_),.p_desc125_p_O_FDEr_mat_regs_(p_desc125_p_O_FDEr_mat_regs_qr_decomp_),.p_desc126_p_O_FDEr_mat_regs_(p_desc126_p_O_FDEr_mat_regs_qr_decomp_),.p_desc127_p_O_FDEr_mat_regs_(p_desc127_p_O_FDEr_mat_regs_qr_decomp_),.p_desc128_p_O_FDEr_mat_regs_(p_desc128_p_O_FDEr_mat_regs_qr_decomp_),.p_desc129_p_O_FDEr_mat_regs_(p_desc129_p_O_FDEr_mat_regs_qr_decomp_),.p_desc130_p_O_FDEr_mat_regs_(p_desc130_p_O_FDEr_mat_regs_qr_decomp_),.p_desc131_p_O_FDEr_mat_regs_(p_desc131_p_O_FDEr_mat_regs_qr_decomp_),.p_desc132_p_O_FDEr_mat_regs_(p_desc132_p_O_FDEr_mat_regs_qr_decomp_),.p_desc133_p_O_FDEr_mat_regs_(p_desc133_p_O_FDEr_mat_regs_qr_decomp_),.p_desc134_p_O_FDEr_mat_regs_(p_desc134_p_O_FDEr_mat_regs_qr_decomp_),.p_desc135_p_O_FDEr_mat_regs_(p_desc135_p_O_FDEr_mat_regs_qr_decomp_),.p_desc136_p_O_FDEr_mat_regs_(p_desc136_p_O_FDEr_mat_regs_qr_decomp_),.p_desc137_p_O_FDEr_mat_regs_(p_desc137_p_O_FDEr_mat_regs_qr_decomp_),.p_desc138_p_O_FDEr_mat_regs_(p_desc138_p_O_FDEr_mat_regs_qr_decomp_),.p_desc139_p_O_FDEr_mat_regs_(p_desc139_p_O_FDEr_mat_regs_qr_decomp_),.p_desc140_p_O_FDEr_mat_regs_(p_desc140_p_O_FDEr_mat_regs_qr_decomp_),.p_desc141_p_O_FDEr_mat_regs_(p_desc141_p_O_FDEr_mat_regs_qr_decomp_),.p_desc142_p_O_FDEr_mat_regs_(p_desc142_p_O_FDEr_mat_regs_qr_decomp_),.p_desc143_p_O_FDEr_mat_regs_(p_desc143_p_O_FDEr_mat_regs_qr_decomp_),.p_desc144_p_O_FDEr_mat_regs_(p_desc144_p_O_FDEr_mat_regs_qr_decomp_),.p_desc145_p_O_FDEr_mat_regs_(p_desc145_p_O_FDEr_mat_regs_qr_decomp_),.p_desc146_p_O_FDEr_mat_regs_(p_desc146_p_O_FDEr_mat_regs_qr_decomp_),.p_desc147_p_O_FDEr_mat_regs_(p_desc147_p_O_FDEr_mat_regs_qr_decomp_),.p_desc148_p_O_FDEr_mat_regs_(p_desc148_p_O_FDEr_mat_regs_qr_decomp_),.p_desc149_p_O_FDEr_mat_regs_(p_desc149_p_O_FDEr_mat_regs_qr_decomp_),.p_desc150_p_O_FDEr_mat_regs_(p_desc150_p_O_FDEr_mat_regs_qr_decomp_),.p_desc151_p_O_FDEr_mat_regs_(p_desc151_p_O_FDEr_mat_regs_qr_decomp_),.p_desc152_p_O_FDEr_mat_regs_(p_desc152_p_O_FDEr_mat_regs_qr_decomp_),.p_desc153_p_O_FDEr_mat_regs_(p_desc153_p_O_FDEr_mat_regs_qr_decomp_),.p_desc154_p_O_FDEr_mat_regs_(p_desc154_p_O_FDEr_mat_regs_qr_decomp_),.p_desc155_p_O_FDEr_mat_regs_(p_desc155_p_O_FDEr_mat_regs_qr_decomp_),.p_desc156_p_O_FDEr_mat_regs_(p_desc156_p_O_FDEr_mat_regs_qr_decomp_),.p_desc157_p_O_FDEr_mat_regs_(p_desc157_p_O_FDEr_mat_regs_qr_decomp_),.p_desc158_p_O_FDEr_mat_regs_(p_desc158_p_O_FDEr_mat_regs_qr_decomp_),.p_desc159_p_O_FDEr_mat_regs_(p_desc159_p_O_FDEr_mat_regs_qr_decomp_),.p_desc160_p_O_FDEr_mat_regs_(p_desc160_p_O_FDEr_mat_regs_qr_decomp_),.p_desc161_p_O_FDEr_mat_regs_(p_desc161_p_O_FDEr_mat_regs_qr_decomp_),.p_desc162_p_O_FDEr_mat_regs_(p_desc162_p_O_FDEr_mat_regs_qr_decomp_),.p_desc163_p_O_FDEr_mat_regs_(p_desc163_p_O_FDEr_mat_regs_qr_decomp_),.p_desc164_p_O_FDEr_mat_regs_(p_desc164_p_O_FDEr_mat_regs_qr_decomp_),.p_desc165_p_O_FDEr_mat_regs_(p_desc165_p_O_FDEr_mat_regs_qr_decomp_),.p_desc166_p_O_FDEr_mat_regs_(p_desc166_p_O_FDEr_mat_regs_qr_decomp_),.p_desc167_p_O_FDEr_mat_regs_(p_desc167_p_O_FDEr_mat_regs_qr_decomp_),.p_desc168_p_O_FDEr_mat_regs_(p_desc168_p_O_FDEr_mat_regs_qr_decomp_),.p_desc169_p_O_FDEr_mat_regs_(p_desc169_p_O_FDEr_mat_regs_qr_decomp_),.p_desc170_p_O_FDEr_mat_regs_(p_desc170_p_O_FDEr_mat_regs_qr_decomp_),.p_desc171_p_O_FDEr_mat_regs_(p_desc171_p_O_FDEr_mat_regs_qr_decomp_),.p_desc172_p_O_FDEr_mat_regs_(p_desc172_p_O_FDEr_mat_regs_qr_decomp_),.p_desc173_p_O_FDEr_mat_regs_(p_desc173_p_O_FDEr_mat_regs_qr_decomp_),.p_desc174_p_O_FDEr_mat_regs_(p_desc174_p_O_FDEr_mat_regs_qr_decomp_),.p_desc175_p_O_FDEr_mat_regs_(p_desc175_p_O_FDEr_mat_regs_qr_decomp_),.p_desc176_p_O_FDEr_mat_regs_(p_desc176_p_O_FDEr_mat_regs_qr_decomp_),.p_desc177_p_O_FDEr_mat_regs_(p_desc177_p_O_FDEr_mat_regs_qr_decomp_),.p_desc178_p_O_FDEr_mat_regs_(p_desc178_p_O_FDEr_mat_regs_qr_decomp_),.p_desc179_p_O_FDEr_mat_regs_(p_desc179_p_O_FDEr_mat_regs_qr_decomp_),.p_desc180_p_O_FDEr_mat_regs_(p_desc180_p_O_FDEr_mat_regs_qr_decomp_),.p_desc181_p_O_FDEr_mat_regs_(p_desc181_p_O_FDEr_mat_regs_qr_decomp_),.p_desc182_p_O_FDEr_mat_regs_(p_desc182_p_O_FDEr_mat_regs_qr_decomp_),.p_desc183_p_O_FDEr_mat_regs_(p_desc183_p_O_FDEr_mat_regs_qr_decomp_),.p_desc184_p_O_FDEr_mat_regs_(p_desc184_p_O_FDEr_mat_regs_qr_decomp_),.p_desc185_p_O_FDEr_mat_regs_(p_desc185_p_O_FDEr_mat_regs_qr_decomp_),.p_desc186_p_O_FDEr_mat_regs_(p_desc186_p_O_FDEr_mat_regs_qr_decomp_),.p_desc187_p_O_FDEr_mat_regs_(p_desc187_p_O_FDEr_mat_regs_qr_decomp_),.p_desc188_p_O_FDEr_mat_regs_(p_desc188_p_O_FDEr_mat_regs_qr_decomp_),.p_desc189_p_O_FDEr_mat_regs_(p_desc189_p_O_FDEr_mat_regs_qr_decomp_),.p_desc190_p_O_FDEr_mat_regs_(p_desc190_p_O_FDEr_mat_regs_qr_decomp_),.p_desc191_p_O_FDEr_mat_regs_(p_desc191_p_O_FDEr_mat_regs_qr_decomp_),.p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_(p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_),.p_desc739_p_O_FDEvec_sub_(p_desc739_p_O_FDEvec_sub_qr_decomp_),.p_desc740_p_O_FDEvec_sub_(p_desc740_p_O_FDEvec_sub_qr_decomp_),.p_desc741_p_O_FDEvec_sub_(p_desc741_p_O_FDEvec_sub_qr_decomp_),.p_desc742_p_O_FDEvec_sub_(p_desc742_p_O_FDEvec_sub_qr_decomp_),.p_desc743_p_O_FDEvec_sub_(p_desc743_p_O_FDEvec_sub_qr_decomp_),.p_desc744_p_O_FDEvec_sub_(p_desc744_p_O_FDEvec_sub_qr_decomp_),.p_desc745_p_O_FDEvec_sub_(p_desc745_p_O_FDEvec_sub_qr_decomp_),.p_desc746_p_O_FDEvec_sub_(p_desc746_p_O_FDEvec_sub_qr_decomp_),.p_desc747_p_O_FDEvec_sub_(p_desc747_p_O_FDEvec_sub_qr_decomp_),.p_desc748_p_O_FDEvec_sub_(p_desc748_p_O_FDEvec_sub_qr_decomp_),.p_desc749_p_O_FDEvec_sub_(p_desc749_p_O_FDEvec_sub_qr_decomp_),.p_desc750_p_O_FDEvec_sub_(p_desc750_p_O_FDEvec_sub_qr_decomp_),.p_desc751_p_O_FDEvec_sub_(p_desc751_p_O_FDEvec_sub_qr_decomp_),.p_desc752_p_O_FDEvec_sub_(p_desc752_p_O_FDEvec_sub_qr_decomp_),.p_desc753_p_O_FDEvec_sub_(p_desc753_p_O_FDEvec_sub_qr_decomp_),.p_desc754_p_O_FDEvec_sub_(p_desc754_p_O_FDEvec_sub_qr_decomp_),.p_desc755_p_O_FDEvec_sub_(p_desc755_p_O_FDEvec_sub_qr_decomp_),.p_desc756_p_O_FDEvec_sub_(p_desc756_p_O_FDEvec_sub_qr_decomp_),.p_desc757_p_O_FDEvec_sub_(p_desc757_p_O_FDEvec_sub_qr_decomp_),.p_desc758_p_O_FDEvec_sub_(p_desc758_p_O_FDEvec_sub_qr_decomp_),.p_desc759_p_O_FDEvec_sub_(p_desc759_p_O_FDEvec_sub_qr_decomp_),.p_desc760_p_O_FDEvec_sub_(p_desc760_p_O_FDEvec_sub_qr_decomp_),.p_desc761_p_O_FDEvec_sub_(p_desc761_p_O_FDEvec_sub_qr_decomp_),.p_desc762_p_O_FDEvec_sub_(p_desc762_p_O_FDEvec_sub_qr_decomp_),.p_desc763_p_O_FDEvec_sub_(p_desc763_p_O_FDEvec_sub_qr_decomp_),.p_desc764_p_O_FDEvec_sub_(p_desc764_p_O_FDEvec_sub_qr_decomp_),.p_desc765_p_O_FDEvec_sub_(p_desc765_p_O_FDEvec_sub_qr_decomp_),.p_desc766_p_O_FDEvec_sub_(p_desc766_p_O_FDEvec_sub_qr_decomp_),.p_desc767_p_O_FDEvec_sub_(p_desc767_p_O_FDEvec_sub_qr_decomp_),.p_desc768_p_O_FDEvec_sub_(p_desc768_p_O_FDEvec_sub_qr_decomp_),.p_desc769_p_O_FDEvec_sub_(p_desc769_p_O_FDEvec_sub_qr_decomp_),.p_desc770_p_O_FDEvec_sub_(p_desc770_p_O_FDEvec_sub_qr_decomp_),.p_desc771_p_O_FDEvec_sub_(p_desc771_p_O_FDEvec_sub_qr_decomp_),.p_desc772_p_O_FDEvec_sub_(p_desc772_p_O_FDEvec_sub_qr_decomp_),.p_desc773_p_O_FDEvec_sub_(p_desc773_p_O_FDEvec_sub_qr_decomp_),.p_desc774_p_O_FDEvec_sub_(p_desc774_p_O_FDEvec_sub_qr_decomp_),.p_desc775_p_O_FDEvec_sub_(p_desc775_p_O_FDEvec_sub_qr_decomp_),.p_desc776_p_O_FDEvec_sub_(p_desc776_p_O_FDEvec_sub_qr_decomp_),.p_desc777_p_O_FDEvec_sub_(p_desc777_p_O_FDEvec_sub_qr_decomp_),.p_desc778_p_O_FDEvec_sub_(p_desc778_p_O_FDEvec_sub_qr_decomp_),.p_desc779_p_O_FDEvec_sub_(p_desc779_p_O_FDEvec_sub_qr_decomp_),.p_desc780_p_O_FDEvec_sub_(p_desc780_p_O_FDEvec_sub_qr_decomp_),.p_desc781_p_O_FDEvec_sub_(p_desc781_p_O_FDEvec_sub_qr_decomp_),.p_desc782_p_O_FDEvec_sub_(p_desc782_p_O_FDEvec_sub_qr_decomp_),.p_desc783_p_O_FDEvec_sub_(p_desc783_p_O_FDEvec_sub_qr_decomp_),.p_desc784_p_O_FDEvec_sub_(p_desc784_p_O_FDEvec_sub_qr_decomp_),.p_desc785_p_O_FDEvec_sub_(p_desc785_p_O_FDEvec_sub_qr_decomp_),.p_desc786_p_O_FDEvec_sub_(p_desc786_p_O_FDEvec_sub_qr_decomp_),.p_desc787_p_O_FDEvec_sub_(p_desc787_p_O_FDEvec_sub_qr_decomp_),.p_desc788_p_O_FDEvec_sub_(p_desc788_p_O_FDEvec_sub_qr_decomp_),.p_desc789_p_O_FDEvec_sub_(p_desc789_p_O_FDEvec_sub_qr_decomp_),.p_desc790_p_O_FDEvec_sub_(p_desc790_p_O_FDEvec_sub_qr_decomp_),.p_desc791_p_O_FDEvec_sub_(p_desc791_p_O_FDEvec_sub_qr_decomp_),.p_desc792_p_O_FDEvec_sub_(p_desc792_p_O_FDEvec_sub_qr_decomp_),.p_desc793_p_O_FDEvec_sub_(p_desc793_p_O_FDEvec_sub_qr_decomp_),.p_desc794_p_O_FDEvec_sub_(p_desc794_p_O_FDEvec_sub_qr_decomp_),.p_desc795_p_O_FDEvec_sub_(p_desc795_p_O_FDEvec_sub_qr_decomp_),.p_desc796_p_O_FDEvec_sub_(p_desc796_p_O_FDEvec_sub_qr_decomp_),.p_desc797_p_O_FDEvec_sub_(p_desc797_p_O_FDEvec_sub_qr_decomp_),.p_desc798_p_O_FDEvec_sub_(p_desc798_p_O_FDEvec_sub_qr_decomp_),.p_desc799_p_O_FDEvec_sub_(p_desc799_p_O_FDEvec_sub_qr_decomp_),.p_desc800_p_O_FDEvec_sub_(p_desc800_p_O_FDEvec_sub_qr_decomp_),.p_desc801_p_O_FDEvec_sub_(p_desc801_p_O_FDEvec_sub_qr_decomp_),.p_desc802_p_O_FDEvec_sub_(p_desc802_p_O_FDEvec_sub_qr_decomp_),.p_desc803_p_O_FDEvec_sub_(p_desc803_p_O_FDEvec_sub_qr_decomp_),.p_desc804_p_O_FDEvec_sub_(p_desc804_p_O_FDEvec_sub_qr_decomp_),.p_desc805_p_O_FDEvec_sub_(p_desc805_p_O_FDEvec_sub_qr_decomp_),.p_desc806_p_O_FDEvec_sub_(p_desc806_p_O_FDEvec_sub_qr_decomp_),.p_desc807_p_O_FDEvec_sub_(p_desc807_p_O_FDEvec_sub_qr_decomp_),.p_desc808_p_O_FDEvec_sub_(p_desc808_p_O_FDEvec_sub_qr_decomp_),.p_desc809_p_O_FDEvec_sub_(p_desc809_p_O_FDEvec_sub_qr_decomp_),.p_desc810_p_O_FDEvec_sub_(p_desc810_p_O_FDEvec_sub_qr_decomp_),.p_desc811_p_O_FDEvec_sub_(p_desc811_p_O_FDEvec_sub_qr_decomp_),.p_desc812_p_O_FDEvec_sub_(p_desc812_p_O_FDEvec_sub_qr_decomp_),.p_desc813_p_O_FDEvec_sub_(p_desc813_p_O_FDEvec_sub_qr_decomp_),.p_desc814_p_O_FDEvec_sub_(p_desc814_p_O_FDEvec_sub_qr_decomp_),.p_desc815_p_O_FDEvec_sub_(p_desc815_p_O_FDEvec_sub_qr_decomp_),.p_desc816_p_O_FDEvec_sub_(p_desc816_p_O_FDEvec_sub_qr_decomp_),.p_desc817_p_O_FDEvec_sub_(p_desc817_p_O_FDEvec_sub_qr_decomp_),.p_desc818_p_O_FDEvec_sub_(p_desc818_p_O_FDEvec_sub_qr_decomp_),.p_desc819_p_O_FDEvec_sub_(p_desc819_p_O_FDEvec_sub_qr_decomp_),.p_desc820_p_O_FDEvec_sub_(p_desc820_p_O_FDEvec_sub_qr_decomp_),.p_desc821_p_O_FDEvec_sub_(p_desc821_p_O_FDEvec_sub_qr_decomp_),.p_desc822_p_O_FDEvec_sub_(p_desc822_p_O_FDEvec_sub_qr_decomp_),.p_desc823_p_O_FDEvec_sub_(p_desc823_p_O_FDEvec_sub_qr_decomp_),.p_desc824_p_O_FDEvec_sub_(p_desc824_p_O_FDEvec_sub_qr_decomp_),.p_desc825_p_O_FDEvec_sub_(p_desc825_p_O_FDEvec_sub_qr_decomp_),.p_desc826_p_O_FDEvec_sub_(p_desc826_p_O_FDEvec_sub_qr_decomp_),.p_desc827_p_O_FDEvec_sub_(p_desc827_p_O_FDEvec_sub_qr_decomp_),.p_desc828_p_O_FDEvec_sub_(p_desc828_p_O_FDEvec_sub_qr_decomp_),.p_desc829_p_O_FDEvec_sub_(p_desc829_p_O_FDEvec_sub_qr_decomp_),.p_desc830_p_O_FDEvec_sub_(p_desc830_p_O_FDEvec_sub_qr_decomp_),.p_desc831_p_O_FDEvec_sub_(p_desc831_p_O_FDEvec_sub_qr_decomp_),.p_desc832_p_O_FDEvec_sub_(p_desc832_p_O_FDEvec_sub_qr_decomp_),.p_desc833_p_O_FDEvec_sub_(p_desc833_p_O_FDEvec_sub_qr_decomp_),.p_desc834_p_O_FDEvec_sub_(p_desc834_p_O_FDEvec_sub_qr_decomp_),.p_output_reg_pipe_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_(p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_),.p_desc318_p_O_FDCinner_prod_(p_desc318_p_O_FDCinner_prod_qr_decomp_),.p_desc319_p_O_FDCinner_prod_(p_desc319_p_O_FDCinner_prod_qr_decomp_),.p_desc320_p_O_FDCinner_prod_(p_desc320_p_O_FDCinner_prod_qr_decomp_),.p_desc321_p_O_FDCinner_prod_(p_desc321_p_O_FDCinner_prod_qr_decomp_),.p_desc322_p_O_FDCinner_prod_(p_desc322_p_O_FDCinner_prod_qr_decomp_),.p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_(p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_),.p_done_Z_p_O_FDCinner_prod_(p_done_Z_p_O_FDCinner_prod_qr_decomp_),.p_acc_enable_Z_p_O_FDCinner_prod_(p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_),.p_desc325_p_O_FDCinner_prod_(p_desc325_p_O_FDCinner_prod_qr_decomp_),.p_desc326_p_O_FDCinner_prod_(p_desc326_p_O_FDCinner_prod_qr_decomp_),.p_desc327_p_O_FDCinner_prod_(p_desc327_p_O_FDCinner_prod_qr_decomp_),.p_desc328_p_O_FDCinner_prod_(p_desc328_p_O_FDCinner_prod_qr_decomp_),.p_desc329_p_O_FDCinner_prod_(p_desc329_p_O_FDCinner_prod_qr_decomp_),.p_desc330_p_O_FDCinner_prod_(p_desc330_p_O_FDCinner_prod_qr_decomp_),.p_desc331_p_O_FDCinner_prod_(p_desc331_p_O_FDCinner_prod_qr_decomp_),.p_desc332_p_O_FDCinner_prod_(p_desc332_p_O_FDCinner_prod_qr_decomp_),.p_desc333_p_O_FDCinner_prod_(p_desc333_p_O_FDCinner_prod_qr_decomp_),.p_desc334_p_O_FDCinner_prod_(p_desc334_p_O_FDCinner_prod_qr_decomp_),.p_desc335_p_O_FDCinner_prod_(p_desc335_p_O_FDCinner_prod_qr_decomp_),.p_desc336_p_O_FDCinner_prod_(p_desc336_p_O_FDCinner_prod_qr_decomp_),.p_desc337_p_O_FDCinner_prod_(p_desc337_p_O_FDCinner_prod_qr_decomp_),.p_desc338_p_O_FDCinner_prod_(p_desc338_p_O_FDCinner_prod_qr_decomp_),.p_desc339_p_O_FDCinner_prod_(p_desc339_p_O_FDCinner_prod_qr_decomp_),.p_desc340_p_O_FDCinner_prod_(p_desc340_p_O_FDCinner_prod_qr_decomp_),.p_desc341_p_O_FDCinner_prod_(p_desc341_p_O_FDCinner_prod_qr_decomp_),.p_desc342_p_O_FDCinner_prod_(p_desc342_p_O_FDCinner_prod_qr_decomp_),.p_desc343_p_O_FDCinner_prod_(p_desc343_p_O_FDCinner_prod_qr_decomp_),.p_desc344_p_O_FDCinner_prod_(p_desc344_p_O_FDCinner_prod_qr_decomp_),.p_desc345_p_O_FDCinner_prod_(p_desc345_p_O_FDCinner_prod_qr_decomp_),.p_desc346_p_O_FDCinner_prod_(p_desc346_p_O_FDCinner_prod_qr_decomp_),.p_desc347_p_O_FDCinner_prod_(p_desc347_p_O_FDCinner_prod_qr_decomp_),.p_desc348_p_O_FDCinner_prod_(p_desc348_p_O_FDCinner_prod_qr_decomp_),.p_desc349_p_O_FDCinner_prod_(p_desc349_p_O_FDCinner_prod_qr_decomp_),.p_desc350_p_O_FDCinner_prod_(p_desc350_p_O_FDCinner_prod_qr_decomp_),.p_desc375_p_O_FDCinner_prod_(p_desc375_p_O_FDCinner_prod_qr_decomp_),.p_desc376_p_O_FDCinner_prod_(p_desc376_p_O_FDCinner_prod_qr_decomp_),.p_desc377_p_O_FDCinner_prod_(p_desc377_p_O_FDCinner_prod_qr_decomp_),.p_desc378_p_O_FDCinner_prod_(p_desc378_p_O_FDCinner_prod_qr_decomp_),.p_desc379_p_O_FDCinner_prod_(p_desc379_p_O_FDCinner_prod_qr_decomp_),.p_desc380_p_O_FDCinner_prod_(p_desc380_p_O_FDCinner_prod_qr_decomp_),.p_desc381_p_O_FDCinner_prod_(p_desc381_p_O_FDCinner_prod_qr_decomp_),.p_desc382_p_O_FDCinner_prod_(p_desc382_p_O_FDCinner_prod_qr_decomp_),.p_desc383_p_O_FDCinner_prod_(p_desc383_p_O_FDCinner_prod_qr_decomp_),.p_desc384_p_O_FDCinner_prod_(p_desc384_p_O_FDCinner_prod_qr_decomp_),.p_desc385_p_O_FDCinner_prod_(p_desc385_p_O_FDCinner_prod_qr_decomp_),.p_desc386_p_O_FDCinner_prod_(p_desc386_p_O_FDCinner_prod_qr_decomp_),.p_desc387_p_O_FDCinner_prod_(p_desc387_p_O_FDCinner_prod_qr_decomp_),.p_desc388_p_O_FDCinner_prod_(p_desc388_p_O_FDCinner_prod_qr_decomp_),.p_desc389_p_O_FDCinner_prod_(p_desc389_p_O_FDCinner_prod_qr_decomp_),.p_desc390_p_O_FDCinner_prod_(p_desc390_p_O_FDCinner_prod_qr_decomp_),.p_desc391_p_O_FDCinner_prod_(p_desc391_p_O_FDCinner_prod_qr_decomp_),.p_desc392_p_O_FDCinner_prod_(p_desc392_p_O_FDCinner_prod_qr_decomp_),.p_desc393_p_O_FDCinner_prod_(p_desc393_p_O_FDCinner_prod_qr_decomp_),.p_desc394_p_O_FDCinner_prod_(p_desc394_p_O_FDCinner_prod_qr_decomp_),.p_desc395_p_O_FDCinner_prod_(p_desc395_p_O_FDCinner_prod_qr_decomp_),.p_desc396_p_O_FDCinner_prod_(p_desc396_p_O_FDCinner_prod_qr_decomp_),.p_desc397_p_O_FDCinner_prod_(p_desc397_p_O_FDCinner_prod_qr_decomp_),.p_desc398_p_O_FDCinner_prod_(p_desc398_p_O_FDCinner_prod_qr_decomp_),.p_done_Z_p_O_FDCinv_sqrt_(p_done_Z_p_O_FDCinv_sqrt_qr_decomp_),.p_desc946_p_O_FDCinv_sqrt_(p_desc946_p_O_FDCinv_sqrt_qr_decomp_),.p_desc947_p_O_FDCinv_sqrt_(p_desc947_p_O_FDCinv_sqrt_qr_decomp_),.p_desc948_p_O_FDCinv_sqrt_(p_desc948_p_O_FDCinv_sqrt_qr_decomp_),.p_desc949_p_O_FDCinv_sqrt_(p_desc949_p_O_FDCinv_sqrt_qr_decomp_),.p_desc950_p_O_FDCinv_sqrt_(p_desc950_p_O_FDCinv_sqrt_qr_decomp_),.p_desc1255_p_O_FDCqr_decomp_ctl_(p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1256_p_O_FDCqr_decomp_ctl_(p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1257_p_O_FDCqr_decomp_ctl_(p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1258_p_O_FDCqr_decomp_ctl_(p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_(p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_(p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_(p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_(p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_(p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1274_p_O_FDCqr_decomp_ctl_(p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_(p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_done_Z_p_O_FDCqr_decomp_ctl_(p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1275_p_O_FDCqr_decomp_ctl_(p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1276_p_O_FDCqr_decomp_ctl_(p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1277_p_O_FDCqr_decomp_ctl_(p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1278_p_O_FDCqr_decomp_ctl_(p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1279_p_O_FDCqr_decomp_ctl_(p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1281_p_O_FDCqr_decomp_ctl_(p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1282_p_O_FDCqr_decomp_ctl_(p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1283_p_O_FDCqr_decomp_ctl_(p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1284_p_O_FDCqr_decomp_ctl_(p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1285_p_O_FDCqr_decomp_ctl_(p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1286_p_O_FDCqr_decomp_ctl_(p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1287_p_O_FDCqr_decomp_ctl_(p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_desc1288_p_O_FDCqr_decomp_ctl_(p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_),.p_acc_clear_Z_p_O_FDPinner_prod_(p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_),.p_desc1265_p_O_FDPqr_decomp_ctl_(p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_),.p_desc1268_p_O_FDPqr_decomp_ctl_(p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_),.p_desc1280_p_O_FDPqr_decomp_ctl_(p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_),.p_desc324_p_O_FDCEinner_prod_(p_desc324_p_O_FDCEinner_prod_qr_decomp_),.p_desc351_p_O_FDCEinner_prod_(p_desc351_p_O_FDCEinner_prod_qr_decomp_),.p_desc352_p_O_FDCEinner_prod_(p_desc352_p_O_FDCEinner_prod_qr_decomp_),.p_desc353_p_O_FDCEinner_prod_(p_desc353_p_O_FDCEinner_prod_qr_decomp_),.p_desc354_p_O_FDCEinner_prod_(p_desc354_p_O_FDCEinner_prod_qr_decomp_),.p_desc355_p_O_FDCEinner_prod_(p_desc355_p_O_FDCEinner_prod_qr_decomp_),.p_desc356_p_O_FDCEinner_prod_(p_desc356_p_O_FDCEinner_prod_qr_decomp_),.p_desc357_p_O_FDCEinner_prod_(p_desc357_p_O_FDCEinner_prod_qr_decomp_),.p_desc358_p_O_FDCEinner_prod_(p_desc358_p_O_FDCEinner_prod_qr_decomp_),.p_desc359_p_O_FDCEinner_prod_(p_desc359_p_O_FDCEinner_prod_qr_decomp_),.p_desc360_p_O_FDCEinner_prod_(p_desc360_p_O_FDCEinner_prod_qr_decomp_),.p_desc361_p_O_FDCEinner_prod_(p_desc361_p_O_FDCEinner_prod_qr_decomp_),.p_desc362_p_O_FDCEinner_prod_(p_desc362_p_O_FDCEinner_prod_qr_decomp_),.p_desc363_p_O_FDCEinner_prod_(p_desc363_p_O_FDCEinner_prod_qr_decomp_),.p_desc364_p_O_FDCEinner_prod_(p_desc364_p_O_FDCEinner_prod_qr_decomp_),.p_desc365_p_O_FDCEinner_prod_(p_desc365_p_O_FDCEinner_prod_qr_decomp_),.p_desc366_p_O_FDCEinner_prod_(p_desc366_p_O_FDCEinner_prod_qr_decomp_),.p_desc367_p_O_FDCEinner_prod_(p_desc367_p_O_FDCEinner_prod_qr_decomp_),.p_desc368_p_O_FDCEinner_prod_(p_desc368_p_O_FDCEinner_prod_qr_decomp_),.p_desc369_p_O_FDCEinner_prod_(p_desc369_p_O_FDCEinner_prod_qr_decomp_),.p_desc370_p_O_FDCEinner_prod_(p_desc370_p_O_FDCEinner_prod_qr_decomp_),.p_desc371_p_O_FDCEinner_prod_(p_desc371_p_O_FDCEinner_prod_qr_decomp_),.p_desc372_p_O_FDCEinner_prod_(p_desc372_p_O_FDCEinner_prod_qr_decomp_),.p_desc373_p_O_FDCEinner_prod_(p_desc373_p_O_FDCEinner_prod_qr_decomp_),.p_desc374_p_O_FDCEinner_prod_(p_desc374_p_O_FDCEinner_prod_qr_decomp_),.p_desc1263_p_O_FDCEqr_decomp_ctl_(p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1264_p_O_FDCEqr_decomp_ctl_(p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1266_p_O_FDCEqr_decomp_ctl_(p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1267_p_O_FDCEqr_decomp_ctl_(p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1269_p_O_FDCEqr_decomp_ctl_(p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1270_p_O_FDCEqr_decomp_ctl_(p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1271_p_O_FDCEqr_decomp_ctl_(p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1272_p_O_FDCEqr_decomp_ctl_(p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_),.p_desc1273_p_O_FDCEqr_decomp_ctl_(p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module qr_wrapper_wrapper_inj (clk,rst,reduced_matrix,start,request_out,valid_out,ready,in_A_r,in_A_i,sigma_in,out_Q_r,out_Q_i,out_R_r,out_R_i,permut,p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_desc951_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc952_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc953_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc954_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc955_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc956_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc957_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc958_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc959_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc960_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc961_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc962_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_,p_desc48_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc49_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc50_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc51_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc52_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc53_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc54_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc55_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc56_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc57_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc58_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc59_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc60_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc61_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc62_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc63_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc64_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc65_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc66_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc67_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc68_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc69_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc70_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc71_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc72_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc73_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc74_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc75_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc76_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc77_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc78_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc79_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc80_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc81_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc82_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc83_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc84_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc85_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc86_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc87_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc88_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc89_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc90_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc91_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc92_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc93_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc94_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc95_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc96_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc97_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc98_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc99_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc100_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc101_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc102_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc103_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc104_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc105_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc106_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc107_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc108_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc109_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc110_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc111_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc112_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc113_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc114_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc115_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc116_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc117_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc118_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc119_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc120_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc121_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc122_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc123_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc124_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc125_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc126_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc127_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc128_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc129_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc130_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc131_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc132_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc133_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc134_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc135_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc136_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc137_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc138_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc139_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc140_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc141_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc142_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc143_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc144_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc145_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc146_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc147_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc148_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc149_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc150_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc151_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc152_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc153_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc154_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc155_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc156_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc157_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc158_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc159_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc160_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc161_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc162_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc163_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc164_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc165_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc166_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc167_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc168_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc169_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc170_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc171_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc172_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc173_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc174_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc175_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc176_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc177_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc178_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc179_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc180_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc181_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc182_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc183_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc184_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc185_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc186_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc187_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc188_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc189_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc190_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_desc191_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_,p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_,p_desc739_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc740_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc741_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc742_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc743_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc744_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc745_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc746_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc747_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc748_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc749_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc750_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc751_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc752_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc753_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc754_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc755_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc756_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc757_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc758_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc759_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc760_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc761_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc762_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc763_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc764_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc765_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc766_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc767_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc768_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc769_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc770_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc771_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc772_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc773_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc774_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc775_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc776_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc777_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc778_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc779_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc780_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc781_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc782_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc783_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc784_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc785_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc786_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc787_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc788_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc789_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc790_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc791_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc792_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc793_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc794_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc795_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc796_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc797_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc798_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc799_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc800_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc801_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc802_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc803_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc804_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc805_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc806_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc807_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc808_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc809_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc810_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc811_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc812_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc813_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc814_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc815_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc816_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc817_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc818_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc819_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc820_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc821_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc822_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc823_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc824_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc825_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc826_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc827_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc828_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc829_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc830_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc831_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc832_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc833_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_desc834_p_O_FDEvec_sub_qr_decomp_qr_wrapper_,p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_,p_desc318_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc319_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc320_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc321_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc322_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_done_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc325_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc326_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc327_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc328_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc329_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc330_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc331_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc332_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc333_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc334_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc335_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc336_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc337_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc338_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc339_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc340_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc341_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc342_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc343_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc344_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc345_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc346_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc347_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc348_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc349_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc350_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc375_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc376_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc377_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc378_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc379_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc380_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc381_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc382_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc383_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc384_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc385_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc386_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc387_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc388_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc389_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc390_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc391_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc392_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc393_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc394_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc395_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc396_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc397_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_desc398_p_O_FDCinner_prod_qr_decomp_qr_wrapper_,p_done_Z_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc946_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc947_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc948_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc949_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc950_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_,p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_,p_start_QR_Z_p_O_FDCqr_wrapper_,p_wr_A_QR_Z_p_O_FDCqr_wrapper_,p_valid_out_Z_p_O_FDCqr_wrapper_,p_ready_Z_p_O_FDCqr_wrapper_,p_red_mat_reg_Z_p_O_FDCqr_wrapper_,p_desc1317_p_O_FDCqr_wrapper_,p_desc1318_p_O_FDCqr_wrapper_,p_desc1319_p_O_FDCqr_wrapper_,p_desc1320_p_O_FDCqr_wrapper_,p_desc1321_p_O_FDCqr_wrapper_,p_desc1322_p_O_FDCqr_wrapper_,p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_qr_wrapper_,p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc324_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc351_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc352_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc353_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc354_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc355_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc356_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc357_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc358_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc359_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc360_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc361_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc362_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc363_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc364_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc365_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc366_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc367_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc368_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc369_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc370_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc371_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc372_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc373_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc374_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_,p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_,p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_);
input clk ;
input rst ;
input reduced_matrix ;
input start ;
input request_out ;
output valid_out ;
output ready ;
input [47:0] in_A_r ;
input [47:0] in_A_i ;
input [11:0] sigma_in ;
output [47:0] out_Q_r ;
output [47:0] out_Q_i ;
output [47:0] out_R_r ;
output [47:0] out_R_i ;
output [7:0] permut ;
wire clk ;
wire rst ;
wire reduced_matrix ;
wire start ;
wire request_out ;
wire valid_out ;
wire ready ;
wire VCC ;
wire GND ;
input p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc951_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc952_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc953_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc954_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc955_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc956_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc957_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc958_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc959_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc960_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc961_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc962_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc48_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc49_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc50_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc51_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc52_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc53_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc54_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc55_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc56_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc57_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc58_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc59_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc60_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc61_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc62_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc63_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc64_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc65_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc66_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc67_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc68_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc69_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc70_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc71_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc72_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc73_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc74_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc75_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc76_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc77_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc78_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc79_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc80_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc81_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc82_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc83_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc84_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc85_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc86_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc87_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc88_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc89_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc90_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc91_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc92_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc93_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc94_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc95_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc96_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc97_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc98_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc99_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc100_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc101_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc102_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc103_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc104_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc105_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc106_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc107_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc108_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc109_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc110_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc111_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc112_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc113_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc114_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc115_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc116_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc117_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc118_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc119_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc120_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc121_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc122_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc123_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc124_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc125_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc126_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc127_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc128_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc129_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc130_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc131_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc132_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc133_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc134_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc135_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc136_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc137_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc138_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc139_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc140_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc141_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc142_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc143_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc144_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc145_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc146_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc147_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc148_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc149_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc150_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc151_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc152_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc153_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc154_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc155_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc156_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc157_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc158_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc159_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc160_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc161_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc162_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc163_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc164_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc165_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc166_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc167_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc168_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc169_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc170_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc171_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc172_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc173_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc174_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc175_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc176_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc177_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc178_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc179_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc180_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc181_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc182_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc183_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc184_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc185_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc186_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc187_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc188_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc189_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc190_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_desc191_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc739_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc740_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc741_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc742_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc743_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc744_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc745_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc746_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc747_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc748_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc749_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc750_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc751_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc752_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc753_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc754_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc755_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc756_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc757_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc758_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc759_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc760_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc761_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc762_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc763_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc764_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc765_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc766_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc767_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc768_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc769_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc770_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc771_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc772_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc773_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc774_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc775_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc776_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc777_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc778_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc779_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc780_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc781_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc782_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc783_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc784_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc785_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc786_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc787_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc788_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc789_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc790_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc791_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc792_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc793_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc794_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc795_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc796_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc797_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc798_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc799_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc800_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc801_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc802_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc803_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc804_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc805_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc806_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc807_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc808_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc809_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc810_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc811_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc812_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc813_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc814_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc815_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc816_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc817_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc818_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc819_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc820_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc821_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc822_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc823_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc824_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc825_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc826_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc827_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc828_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc829_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc830_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc831_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc832_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc833_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_desc834_p_O_FDEvec_sub_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc318_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc319_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc320_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc321_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc322_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_done_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc325_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc326_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc327_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc328_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc329_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc330_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc331_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc332_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc333_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc334_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc335_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc336_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc337_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc338_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc339_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc340_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc341_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc342_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc343_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc344_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc345_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc346_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc347_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc348_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc349_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc350_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc375_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc376_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc377_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc378_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc379_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc380_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc381_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc382_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc383_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc384_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc385_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc386_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc387_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc388_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc389_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc390_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc391_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc392_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc393_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc394_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc395_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc396_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc397_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc398_p_O_FDCinner_prod_qr_decomp_qr_wrapper_ ;
input p_done_Z_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc946_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc947_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc948_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc949_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc950_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_ ;
input p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_start_QR_Z_p_O_FDCqr_wrapper_ ;
input p_wr_A_QR_Z_p_O_FDCqr_wrapper_ ;
input p_valid_out_Z_p_O_FDCqr_wrapper_ ;
input p_ready_Z_p_O_FDCqr_wrapper_ ;
input p_red_mat_reg_Z_p_O_FDCqr_wrapper_ ;
input p_desc1317_p_O_FDCqr_wrapper_ ;
input p_desc1318_p_O_FDCqr_wrapper_ ;
input p_desc1319_p_O_FDCqr_wrapper_ ;
input p_desc1320_p_O_FDCqr_wrapper_ ;
input p_desc1321_p_O_FDCqr_wrapper_ ;
input p_desc1322_p_O_FDCqr_wrapper_ ;
input p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc324_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc351_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc352_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc353_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc354_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc355_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc356_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc357_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc358_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc359_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc360_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc361_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc362_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc363_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc364_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc365_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc366_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc367_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc368_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc369_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc370_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc371_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc372_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc373_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc374_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_ ;
input p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
input p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_ ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  qr_wrapper_inj qr_wrapper_inst(.out_Q_r(out_Q_r[47:0]),.out_Q_i(out_Q_i[47:0]),.out_R_i(out_R_i[47:12]),.out_R_r(out_R_r[47:0]),.in_A_r(in_A_r[47:0]),.in_A_i(in_A_i[47:0]),.clk(clk),.rst(rst),.valid_out(valid_out),.ready(ready),.request_out(request_out),.start(start),.reduced_matrix(reduced_matrix),.p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_desc951_p_O_FDEinv_sqrt_qr_decomp_(p_desc951_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc952_p_O_FDEinv_sqrt_qr_decomp_(p_desc952_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc953_p_O_FDEinv_sqrt_qr_decomp_(p_desc953_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc954_p_O_FDEinv_sqrt_qr_decomp_(p_desc954_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc955_p_O_FDEinv_sqrt_qr_decomp_(p_desc955_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc956_p_O_FDEinv_sqrt_qr_decomp_(p_desc956_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc957_p_O_FDEinv_sqrt_qr_decomp_(p_desc957_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc958_p_O_FDEinv_sqrt_qr_decomp_(p_desc958_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc959_p_O_FDEinv_sqrt_qr_decomp_(p_desc959_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc960_p_O_FDEinv_sqrt_qr_decomp_(p_desc960_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc961_p_O_FDEinv_sqrt_qr_decomp_(p_desc961_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc962_p_O_FDEinv_sqrt_qr_decomp_(p_desc962_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_),.p_desc48_p_O_FDEr_mat_regs_qr_decomp_(p_desc48_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc49_p_O_FDEr_mat_regs_qr_decomp_(p_desc49_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc50_p_O_FDEr_mat_regs_qr_decomp_(p_desc50_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc51_p_O_FDEr_mat_regs_qr_decomp_(p_desc51_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc52_p_O_FDEr_mat_regs_qr_decomp_(p_desc52_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc53_p_O_FDEr_mat_regs_qr_decomp_(p_desc53_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc54_p_O_FDEr_mat_regs_qr_decomp_(p_desc54_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc55_p_O_FDEr_mat_regs_qr_decomp_(p_desc55_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc56_p_O_FDEr_mat_regs_qr_decomp_(p_desc56_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc57_p_O_FDEr_mat_regs_qr_decomp_(p_desc57_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc58_p_O_FDEr_mat_regs_qr_decomp_(p_desc58_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc59_p_O_FDEr_mat_regs_qr_decomp_(p_desc59_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc60_p_O_FDEr_mat_regs_qr_decomp_(p_desc60_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc61_p_O_FDEr_mat_regs_qr_decomp_(p_desc61_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc62_p_O_FDEr_mat_regs_qr_decomp_(p_desc62_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc63_p_O_FDEr_mat_regs_qr_decomp_(p_desc63_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc64_p_O_FDEr_mat_regs_qr_decomp_(p_desc64_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc65_p_O_FDEr_mat_regs_qr_decomp_(p_desc65_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc66_p_O_FDEr_mat_regs_qr_decomp_(p_desc66_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc67_p_O_FDEr_mat_regs_qr_decomp_(p_desc67_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc68_p_O_FDEr_mat_regs_qr_decomp_(p_desc68_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc69_p_O_FDEr_mat_regs_qr_decomp_(p_desc69_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc70_p_O_FDEr_mat_regs_qr_decomp_(p_desc70_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc71_p_O_FDEr_mat_regs_qr_decomp_(p_desc71_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc72_p_O_FDEr_mat_regs_qr_decomp_(p_desc72_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc73_p_O_FDEr_mat_regs_qr_decomp_(p_desc73_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc74_p_O_FDEr_mat_regs_qr_decomp_(p_desc74_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc75_p_O_FDEr_mat_regs_qr_decomp_(p_desc75_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc76_p_O_FDEr_mat_regs_qr_decomp_(p_desc76_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc77_p_O_FDEr_mat_regs_qr_decomp_(p_desc77_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc78_p_O_FDEr_mat_regs_qr_decomp_(p_desc78_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc79_p_O_FDEr_mat_regs_qr_decomp_(p_desc79_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc80_p_O_FDEr_mat_regs_qr_decomp_(p_desc80_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc81_p_O_FDEr_mat_regs_qr_decomp_(p_desc81_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc82_p_O_FDEr_mat_regs_qr_decomp_(p_desc82_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc83_p_O_FDEr_mat_regs_qr_decomp_(p_desc83_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc84_p_O_FDEr_mat_regs_qr_decomp_(p_desc84_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc85_p_O_FDEr_mat_regs_qr_decomp_(p_desc85_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc86_p_O_FDEr_mat_regs_qr_decomp_(p_desc86_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc87_p_O_FDEr_mat_regs_qr_decomp_(p_desc87_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc88_p_O_FDEr_mat_regs_qr_decomp_(p_desc88_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc89_p_O_FDEr_mat_regs_qr_decomp_(p_desc89_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc90_p_O_FDEr_mat_regs_qr_decomp_(p_desc90_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc91_p_O_FDEr_mat_regs_qr_decomp_(p_desc91_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc92_p_O_FDEr_mat_regs_qr_decomp_(p_desc92_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc93_p_O_FDEr_mat_regs_qr_decomp_(p_desc93_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc94_p_O_FDEr_mat_regs_qr_decomp_(p_desc94_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc95_p_O_FDEr_mat_regs_qr_decomp_(p_desc95_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc96_p_O_FDEr_mat_regs_qr_decomp_(p_desc96_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc97_p_O_FDEr_mat_regs_qr_decomp_(p_desc97_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc98_p_O_FDEr_mat_regs_qr_decomp_(p_desc98_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc99_p_O_FDEr_mat_regs_qr_decomp_(p_desc99_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc100_p_O_FDEr_mat_regs_qr_decomp_(p_desc100_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc101_p_O_FDEr_mat_regs_qr_decomp_(p_desc101_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc102_p_O_FDEr_mat_regs_qr_decomp_(p_desc102_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc103_p_O_FDEr_mat_regs_qr_decomp_(p_desc103_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc104_p_O_FDEr_mat_regs_qr_decomp_(p_desc104_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc105_p_O_FDEr_mat_regs_qr_decomp_(p_desc105_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc106_p_O_FDEr_mat_regs_qr_decomp_(p_desc106_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc107_p_O_FDEr_mat_regs_qr_decomp_(p_desc107_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc108_p_O_FDEr_mat_regs_qr_decomp_(p_desc108_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc109_p_O_FDEr_mat_regs_qr_decomp_(p_desc109_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc110_p_O_FDEr_mat_regs_qr_decomp_(p_desc110_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc111_p_O_FDEr_mat_regs_qr_decomp_(p_desc111_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc112_p_O_FDEr_mat_regs_qr_decomp_(p_desc112_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc113_p_O_FDEr_mat_regs_qr_decomp_(p_desc113_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc114_p_O_FDEr_mat_regs_qr_decomp_(p_desc114_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc115_p_O_FDEr_mat_regs_qr_decomp_(p_desc115_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc116_p_O_FDEr_mat_regs_qr_decomp_(p_desc116_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc117_p_O_FDEr_mat_regs_qr_decomp_(p_desc117_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc118_p_O_FDEr_mat_regs_qr_decomp_(p_desc118_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc119_p_O_FDEr_mat_regs_qr_decomp_(p_desc119_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc120_p_O_FDEr_mat_regs_qr_decomp_(p_desc120_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc121_p_O_FDEr_mat_regs_qr_decomp_(p_desc121_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc122_p_O_FDEr_mat_regs_qr_decomp_(p_desc122_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc123_p_O_FDEr_mat_regs_qr_decomp_(p_desc123_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc124_p_O_FDEr_mat_regs_qr_decomp_(p_desc124_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc125_p_O_FDEr_mat_regs_qr_decomp_(p_desc125_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc126_p_O_FDEr_mat_regs_qr_decomp_(p_desc126_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc127_p_O_FDEr_mat_regs_qr_decomp_(p_desc127_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc128_p_O_FDEr_mat_regs_qr_decomp_(p_desc128_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc129_p_O_FDEr_mat_regs_qr_decomp_(p_desc129_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc130_p_O_FDEr_mat_regs_qr_decomp_(p_desc130_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc131_p_O_FDEr_mat_regs_qr_decomp_(p_desc131_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc132_p_O_FDEr_mat_regs_qr_decomp_(p_desc132_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc133_p_O_FDEr_mat_regs_qr_decomp_(p_desc133_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc134_p_O_FDEr_mat_regs_qr_decomp_(p_desc134_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc135_p_O_FDEr_mat_regs_qr_decomp_(p_desc135_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc136_p_O_FDEr_mat_regs_qr_decomp_(p_desc136_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc137_p_O_FDEr_mat_regs_qr_decomp_(p_desc137_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc138_p_O_FDEr_mat_regs_qr_decomp_(p_desc138_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc139_p_O_FDEr_mat_regs_qr_decomp_(p_desc139_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc140_p_O_FDEr_mat_regs_qr_decomp_(p_desc140_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc141_p_O_FDEr_mat_regs_qr_decomp_(p_desc141_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc142_p_O_FDEr_mat_regs_qr_decomp_(p_desc142_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc143_p_O_FDEr_mat_regs_qr_decomp_(p_desc143_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc144_p_O_FDEr_mat_regs_qr_decomp_(p_desc144_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc145_p_O_FDEr_mat_regs_qr_decomp_(p_desc145_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc146_p_O_FDEr_mat_regs_qr_decomp_(p_desc146_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc147_p_O_FDEr_mat_regs_qr_decomp_(p_desc147_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc148_p_O_FDEr_mat_regs_qr_decomp_(p_desc148_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc149_p_O_FDEr_mat_regs_qr_decomp_(p_desc149_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc150_p_O_FDEr_mat_regs_qr_decomp_(p_desc150_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc151_p_O_FDEr_mat_regs_qr_decomp_(p_desc151_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc152_p_O_FDEr_mat_regs_qr_decomp_(p_desc152_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc153_p_O_FDEr_mat_regs_qr_decomp_(p_desc153_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc154_p_O_FDEr_mat_regs_qr_decomp_(p_desc154_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc155_p_O_FDEr_mat_regs_qr_decomp_(p_desc155_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc156_p_O_FDEr_mat_regs_qr_decomp_(p_desc156_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc157_p_O_FDEr_mat_regs_qr_decomp_(p_desc157_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc158_p_O_FDEr_mat_regs_qr_decomp_(p_desc158_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc159_p_O_FDEr_mat_regs_qr_decomp_(p_desc159_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc160_p_O_FDEr_mat_regs_qr_decomp_(p_desc160_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc161_p_O_FDEr_mat_regs_qr_decomp_(p_desc161_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc162_p_O_FDEr_mat_regs_qr_decomp_(p_desc162_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc163_p_O_FDEr_mat_regs_qr_decomp_(p_desc163_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc164_p_O_FDEr_mat_regs_qr_decomp_(p_desc164_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc165_p_O_FDEr_mat_regs_qr_decomp_(p_desc165_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc166_p_O_FDEr_mat_regs_qr_decomp_(p_desc166_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc167_p_O_FDEr_mat_regs_qr_decomp_(p_desc167_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc168_p_O_FDEr_mat_regs_qr_decomp_(p_desc168_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc169_p_O_FDEr_mat_regs_qr_decomp_(p_desc169_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc170_p_O_FDEr_mat_regs_qr_decomp_(p_desc170_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc171_p_O_FDEr_mat_regs_qr_decomp_(p_desc171_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc172_p_O_FDEr_mat_regs_qr_decomp_(p_desc172_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc173_p_O_FDEr_mat_regs_qr_decomp_(p_desc173_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc174_p_O_FDEr_mat_regs_qr_decomp_(p_desc174_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc175_p_O_FDEr_mat_regs_qr_decomp_(p_desc175_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc176_p_O_FDEr_mat_regs_qr_decomp_(p_desc176_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc177_p_O_FDEr_mat_regs_qr_decomp_(p_desc177_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc178_p_O_FDEr_mat_regs_qr_decomp_(p_desc178_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc179_p_O_FDEr_mat_regs_qr_decomp_(p_desc179_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc180_p_O_FDEr_mat_regs_qr_decomp_(p_desc180_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc181_p_O_FDEr_mat_regs_qr_decomp_(p_desc181_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc182_p_O_FDEr_mat_regs_qr_decomp_(p_desc182_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc183_p_O_FDEr_mat_regs_qr_decomp_(p_desc183_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc184_p_O_FDEr_mat_regs_qr_decomp_(p_desc184_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc185_p_O_FDEr_mat_regs_qr_decomp_(p_desc185_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc186_p_O_FDEr_mat_regs_qr_decomp_(p_desc186_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc187_p_O_FDEr_mat_regs_qr_decomp_(p_desc187_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc188_p_O_FDEr_mat_regs_qr_decomp_(p_desc188_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc189_p_O_FDEr_mat_regs_qr_decomp_(p_desc189_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc190_p_O_FDEr_mat_regs_qr_decomp_(p_desc190_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_desc191_p_O_FDEr_mat_regs_qr_decomp_(p_desc191_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_),.p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_(p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_),.p_desc739_p_O_FDEvec_sub_qr_decomp_(p_desc739_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc740_p_O_FDEvec_sub_qr_decomp_(p_desc740_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc741_p_O_FDEvec_sub_qr_decomp_(p_desc741_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc742_p_O_FDEvec_sub_qr_decomp_(p_desc742_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc743_p_O_FDEvec_sub_qr_decomp_(p_desc743_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc744_p_O_FDEvec_sub_qr_decomp_(p_desc744_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc745_p_O_FDEvec_sub_qr_decomp_(p_desc745_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc746_p_O_FDEvec_sub_qr_decomp_(p_desc746_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc747_p_O_FDEvec_sub_qr_decomp_(p_desc747_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc748_p_O_FDEvec_sub_qr_decomp_(p_desc748_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc749_p_O_FDEvec_sub_qr_decomp_(p_desc749_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc750_p_O_FDEvec_sub_qr_decomp_(p_desc750_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc751_p_O_FDEvec_sub_qr_decomp_(p_desc751_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc752_p_O_FDEvec_sub_qr_decomp_(p_desc752_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc753_p_O_FDEvec_sub_qr_decomp_(p_desc753_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc754_p_O_FDEvec_sub_qr_decomp_(p_desc754_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc755_p_O_FDEvec_sub_qr_decomp_(p_desc755_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc756_p_O_FDEvec_sub_qr_decomp_(p_desc756_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc757_p_O_FDEvec_sub_qr_decomp_(p_desc757_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc758_p_O_FDEvec_sub_qr_decomp_(p_desc758_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc759_p_O_FDEvec_sub_qr_decomp_(p_desc759_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc760_p_O_FDEvec_sub_qr_decomp_(p_desc760_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc761_p_O_FDEvec_sub_qr_decomp_(p_desc761_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc762_p_O_FDEvec_sub_qr_decomp_(p_desc762_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc763_p_O_FDEvec_sub_qr_decomp_(p_desc763_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc764_p_O_FDEvec_sub_qr_decomp_(p_desc764_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc765_p_O_FDEvec_sub_qr_decomp_(p_desc765_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc766_p_O_FDEvec_sub_qr_decomp_(p_desc766_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc767_p_O_FDEvec_sub_qr_decomp_(p_desc767_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc768_p_O_FDEvec_sub_qr_decomp_(p_desc768_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc769_p_O_FDEvec_sub_qr_decomp_(p_desc769_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc770_p_O_FDEvec_sub_qr_decomp_(p_desc770_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc771_p_O_FDEvec_sub_qr_decomp_(p_desc771_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc772_p_O_FDEvec_sub_qr_decomp_(p_desc772_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc773_p_O_FDEvec_sub_qr_decomp_(p_desc773_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc774_p_O_FDEvec_sub_qr_decomp_(p_desc774_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc775_p_O_FDEvec_sub_qr_decomp_(p_desc775_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc776_p_O_FDEvec_sub_qr_decomp_(p_desc776_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc777_p_O_FDEvec_sub_qr_decomp_(p_desc777_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc778_p_O_FDEvec_sub_qr_decomp_(p_desc778_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc779_p_O_FDEvec_sub_qr_decomp_(p_desc779_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc780_p_O_FDEvec_sub_qr_decomp_(p_desc780_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc781_p_O_FDEvec_sub_qr_decomp_(p_desc781_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc782_p_O_FDEvec_sub_qr_decomp_(p_desc782_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc783_p_O_FDEvec_sub_qr_decomp_(p_desc783_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc784_p_O_FDEvec_sub_qr_decomp_(p_desc784_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc785_p_O_FDEvec_sub_qr_decomp_(p_desc785_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc786_p_O_FDEvec_sub_qr_decomp_(p_desc786_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc787_p_O_FDEvec_sub_qr_decomp_(p_desc787_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc788_p_O_FDEvec_sub_qr_decomp_(p_desc788_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc789_p_O_FDEvec_sub_qr_decomp_(p_desc789_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc790_p_O_FDEvec_sub_qr_decomp_(p_desc790_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc791_p_O_FDEvec_sub_qr_decomp_(p_desc791_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc792_p_O_FDEvec_sub_qr_decomp_(p_desc792_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc793_p_O_FDEvec_sub_qr_decomp_(p_desc793_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc794_p_O_FDEvec_sub_qr_decomp_(p_desc794_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc795_p_O_FDEvec_sub_qr_decomp_(p_desc795_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc796_p_O_FDEvec_sub_qr_decomp_(p_desc796_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc797_p_O_FDEvec_sub_qr_decomp_(p_desc797_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc798_p_O_FDEvec_sub_qr_decomp_(p_desc798_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc799_p_O_FDEvec_sub_qr_decomp_(p_desc799_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc800_p_O_FDEvec_sub_qr_decomp_(p_desc800_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc801_p_O_FDEvec_sub_qr_decomp_(p_desc801_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc802_p_O_FDEvec_sub_qr_decomp_(p_desc802_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc803_p_O_FDEvec_sub_qr_decomp_(p_desc803_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc804_p_O_FDEvec_sub_qr_decomp_(p_desc804_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc805_p_O_FDEvec_sub_qr_decomp_(p_desc805_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc806_p_O_FDEvec_sub_qr_decomp_(p_desc806_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc807_p_O_FDEvec_sub_qr_decomp_(p_desc807_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc808_p_O_FDEvec_sub_qr_decomp_(p_desc808_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc809_p_O_FDEvec_sub_qr_decomp_(p_desc809_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc810_p_O_FDEvec_sub_qr_decomp_(p_desc810_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc811_p_O_FDEvec_sub_qr_decomp_(p_desc811_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc812_p_O_FDEvec_sub_qr_decomp_(p_desc812_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc813_p_O_FDEvec_sub_qr_decomp_(p_desc813_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc814_p_O_FDEvec_sub_qr_decomp_(p_desc814_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc815_p_O_FDEvec_sub_qr_decomp_(p_desc815_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc816_p_O_FDEvec_sub_qr_decomp_(p_desc816_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc817_p_O_FDEvec_sub_qr_decomp_(p_desc817_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc818_p_O_FDEvec_sub_qr_decomp_(p_desc818_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc819_p_O_FDEvec_sub_qr_decomp_(p_desc819_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc820_p_O_FDEvec_sub_qr_decomp_(p_desc820_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc821_p_O_FDEvec_sub_qr_decomp_(p_desc821_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc822_p_O_FDEvec_sub_qr_decomp_(p_desc822_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc823_p_O_FDEvec_sub_qr_decomp_(p_desc823_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc824_p_O_FDEvec_sub_qr_decomp_(p_desc824_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc825_p_O_FDEvec_sub_qr_decomp_(p_desc825_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc826_p_O_FDEvec_sub_qr_decomp_(p_desc826_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc827_p_O_FDEvec_sub_qr_decomp_(p_desc827_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc828_p_O_FDEvec_sub_qr_decomp_(p_desc828_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc829_p_O_FDEvec_sub_qr_decomp_(p_desc829_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc830_p_O_FDEvec_sub_qr_decomp_(p_desc830_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc831_p_O_FDEvec_sub_qr_decomp_(p_desc831_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc832_p_O_FDEvec_sub_qr_decomp_(p_desc832_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc833_p_O_FDEvec_sub_qr_decomp_(p_desc833_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_desc834_p_O_FDEvec_sub_qr_decomp_(p_desc834_p_O_FDEvec_sub_qr_decomp_qr_wrapper_),.p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_(p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_),.p_desc318_p_O_FDCinner_prod_qr_decomp_(p_desc318_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc319_p_O_FDCinner_prod_qr_decomp_(p_desc319_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc320_p_O_FDCinner_prod_qr_decomp_(p_desc320_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc321_p_O_FDCinner_prod_qr_decomp_(p_desc321_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc322_p_O_FDCinner_prod_qr_decomp_(p_desc322_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_(p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_done_Z_p_O_FDCinner_prod_qr_decomp_(p_done_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_(p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc325_p_O_FDCinner_prod_qr_decomp_(p_desc325_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc326_p_O_FDCinner_prod_qr_decomp_(p_desc326_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc327_p_O_FDCinner_prod_qr_decomp_(p_desc327_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc328_p_O_FDCinner_prod_qr_decomp_(p_desc328_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc329_p_O_FDCinner_prod_qr_decomp_(p_desc329_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc330_p_O_FDCinner_prod_qr_decomp_(p_desc330_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc331_p_O_FDCinner_prod_qr_decomp_(p_desc331_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc332_p_O_FDCinner_prod_qr_decomp_(p_desc332_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc333_p_O_FDCinner_prod_qr_decomp_(p_desc333_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc334_p_O_FDCinner_prod_qr_decomp_(p_desc334_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc335_p_O_FDCinner_prod_qr_decomp_(p_desc335_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc336_p_O_FDCinner_prod_qr_decomp_(p_desc336_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc337_p_O_FDCinner_prod_qr_decomp_(p_desc337_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc338_p_O_FDCinner_prod_qr_decomp_(p_desc338_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc339_p_O_FDCinner_prod_qr_decomp_(p_desc339_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc340_p_O_FDCinner_prod_qr_decomp_(p_desc340_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc341_p_O_FDCinner_prod_qr_decomp_(p_desc341_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc342_p_O_FDCinner_prod_qr_decomp_(p_desc342_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc343_p_O_FDCinner_prod_qr_decomp_(p_desc343_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc344_p_O_FDCinner_prod_qr_decomp_(p_desc344_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc345_p_O_FDCinner_prod_qr_decomp_(p_desc345_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc346_p_O_FDCinner_prod_qr_decomp_(p_desc346_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc347_p_O_FDCinner_prod_qr_decomp_(p_desc347_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc348_p_O_FDCinner_prod_qr_decomp_(p_desc348_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc349_p_O_FDCinner_prod_qr_decomp_(p_desc349_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc350_p_O_FDCinner_prod_qr_decomp_(p_desc350_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc375_p_O_FDCinner_prod_qr_decomp_(p_desc375_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc376_p_O_FDCinner_prod_qr_decomp_(p_desc376_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc377_p_O_FDCinner_prod_qr_decomp_(p_desc377_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc378_p_O_FDCinner_prod_qr_decomp_(p_desc378_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc379_p_O_FDCinner_prod_qr_decomp_(p_desc379_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc380_p_O_FDCinner_prod_qr_decomp_(p_desc380_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc381_p_O_FDCinner_prod_qr_decomp_(p_desc381_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc382_p_O_FDCinner_prod_qr_decomp_(p_desc382_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc383_p_O_FDCinner_prod_qr_decomp_(p_desc383_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc384_p_O_FDCinner_prod_qr_decomp_(p_desc384_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc385_p_O_FDCinner_prod_qr_decomp_(p_desc385_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc386_p_O_FDCinner_prod_qr_decomp_(p_desc386_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc387_p_O_FDCinner_prod_qr_decomp_(p_desc387_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc388_p_O_FDCinner_prod_qr_decomp_(p_desc388_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc389_p_O_FDCinner_prod_qr_decomp_(p_desc389_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc390_p_O_FDCinner_prod_qr_decomp_(p_desc390_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc391_p_O_FDCinner_prod_qr_decomp_(p_desc391_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc392_p_O_FDCinner_prod_qr_decomp_(p_desc392_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc393_p_O_FDCinner_prod_qr_decomp_(p_desc393_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc394_p_O_FDCinner_prod_qr_decomp_(p_desc394_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc395_p_O_FDCinner_prod_qr_decomp_(p_desc395_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc396_p_O_FDCinner_prod_qr_decomp_(p_desc396_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc397_p_O_FDCinner_prod_qr_decomp_(p_desc397_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_desc398_p_O_FDCinner_prod_qr_decomp_(p_desc398_p_O_FDCinner_prod_qr_decomp_qr_wrapper_),.p_done_Z_p_O_FDCinv_sqrt_qr_decomp_(p_done_Z_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc946_p_O_FDCinv_sqrt_qr_decomp_(p_desc946_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc947_p_O_FDCinv_sqrt_qr_decomp_(p_desc947_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc948_p_O_FDCinv_sqrt_qr_decomp_(p_desc948_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc949_p_O_FDCinv_sqrt_qr_decomp_(p_desc949_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc950_p_O_FDCinv_sqrt_qr_decomp_(p_desc950_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_),.p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_(p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_(p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_start_QR_Z_p_O_FDC(p_start_QR_Z_p_O_FDCqr_wrapper_),.p_wr_A_QR_Z_p_O_FDC(p_wr_A_QR_Z_p_O_FDCqr_wrapper_),.p_valid_out_Z_p_O_FDC(p_valid_out_Z_p_O_FDCqr_wrapper_),.p_ready_Z_p_O_FDC(p_ready_Z_p_O_FDCqr_wrapper_),.p_red_mat_reg_Z_p_O_FDC(p_red_mat_reg_Z_p_O_FDCqr_wrapper_),.p_desc1317_p_O_FDC(p_desc1317_p_O_FDCqr_wrapper_),.p_desc1318_p_O_FDC(p_desc1318_p_O_FDCqr_wrapper_),.p_desc1319_p_O_FDC(p_desc1319_p_O_FDCqr_wrapper_),.p_desc1320_p_O_FDC(p_desc1320_p_O_FDCqr_wrapper_),.p_desc1321_p_O_FDC(p_desc1321_p_O_FDCqr_wrapper_),.p_desc1322_p_O_FDC(p_desc1322_p_O_FDCqr_wrapper_),.p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_(p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_qr_wrapper_),.p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_(p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_(p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_(p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc324_p_O_FDCEinner_prod_qr_decomp_(p_desc324_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc351_p_O_FDCEinner_prod_qr_decomp_(p_desc351_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc352_p_O_FDCEinner_prod_qr_decomp_(p_desc352_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc353_p_O_FDCEinner_prod_qr_decomp_(p_desc353_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc354_p_O_FDCEinner_prod_qr_decomp_(p_desc354_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc355_p_O_FDCEinner_prod_qr_decomp_(p_desc355_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc356_p_O_FDCEinner_prod_qr_decomp_(p_desc356_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc357_p_O_FDCEinner_prod_qr_decomp_(p_desc357_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc358_p_O_FDCEinner_prod_qr_decomp_(p_desc358_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc359_p_O_FDCEinner_prod_qr_decomp_(p_desc359_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc360_p_O_FDCEinner_prod_qr_decomp_(p_desc360_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc361_p_O_FDCEinner_prod_qr_decomp_(p_desc361_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc362_p_O_FDCEinner_prod_qr_decomp_(p_desc362_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc363_p_O_FDCEinner_prod_qr_decomp_(p_desc363_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc364_p_O_FDCEinner_prod_qr_decomp_(p_desc364_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc365_p_O_FDCEinner_prod_qr_decomp_(p_desc365_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc366_p_O_FDCEinner_prod_qr_decomp_(p_desc366_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc367_p_O_FDCEinner_prod_qr_decomp_(p_desc367_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc368_p_O_FDCEinner_prod_qr_decomp_(p_desc368_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc369_p_O_FDCEinner_prod_qr_decomp_(p_desc369_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc370_p_O_FDCEinner_prod_qr_decomp_(p_desc370_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc371_p_O_FDCEinner_prod_qr_decomp_(p_desc371_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc372_p_O_FDCEinner_prod_qr_decomp_(p_desc372_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc373_p_O_FDCEinner_prod_qr_decomp_(p_desc373_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc374_p_O_FDCEinner_prod_qr_decomp_(p_desc374_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_),.p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_),.p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_(p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_));
assign out_R_i[0:0]=GND;
assign out_R_i[1:1]=GND;
assign out_R_i[2:2]=GND;
assign out_R_i[3:3]=GND;
assign out_R_i[4:4]=GND;
assign out_R_i[5:5]=GND;
assign out_R_i[6:6]=GND;
assign out_R_i[7:7]=GND;
assign out_R_i[8:8]=GND;
assign out_R_i[9:9]=GND;
assign out_R_i[10:10]=GND;
assign out_R_i[11:11]=GND;
assign permut[0:0]=GND;
assign permut[1:1]=GND;
assign permut[2:2]=GND;
assign permut[3:3]=GND;
assign permut[4:4]=GND;
assign permut[5:5]=GND;
assign permut[6:6]=GND;
assign permut[7:7]=GND;
endmodule
module r_mat_regs_inj (row_sel_R,col_sel_R_mux_i_m3_lut6_2_O6,col_sel_R_mux_i_m3_lut6_2_O5,single_in_r_R_mux,wr_en_AQ_sel,col_sel_R,col_sel_R_int,out_R_i,out_R_r,wr_en_R,N_28_i,clk,N_30_i,N_32_i,N_34_i,N_383_i,N_384_i,N_385_i,N_386_i,N_387_i,N_388_i,N_389_i,N_390_i,N_391_i,N_392_i,N_393_i,N_394_i,N_395_i,N_396_i,N_397_i,N_398_i,N_399_i,N_400_i,N_401_i,p_desc48_p_O_FDE,p_desc49_p_O_FDE,p_desc50_p_O_FDE,p_desc51_p_O_FDE,p_desc52_p_O_FDE,p_desc53_p_O_FDE,p_desc54_p_O_FDE,p_desc55_p_O_FDE,p_desc56_p_O_FDE,p_desc57_p_O_FDE,p_desc58_p_O_FDE,p_desc59_p_O_FDE,p_desc60_p_O_FDE,p_desc61_p_O_FDE,p_desc62_p_O_FDE,p_desc63_p_O_FDE,p_desc64_p_O_FDE,p_desc65_p_O_FDE,p_desc66_p_O_FDE,p_desc67_p_O_FDE,p_desc68_p_O_FDE,p_desc69_p_O_FDE,p_desc70_p_O_FDE,p_desc71_p_O_FDE,p_desc72_p_O_FDE,p_desc73_p_O_FDE,p_desc74_p_O_FDE,p_desc75_p_O_FDE,p_desc76_p_O_FDE,p_desc77_p_O_FDE,p_desc78_p_O_FDE,p_desc79_p_O_FDE,p_desc80_p_O_FDE,p_desc81_p_O_FDE,p_desc82_p_O_FDE,p_desc83_p_O_FDE,p_desc84_p_O_FDE,p_desc85_p_O_FDE,p_desc86_p_O_FDE,p_desc87_p_O_FDE,p_desc88_p_O_FDE,p_desc89_p_O_FDE,p_desc90_p_O_FDE,p_desc91_p_O_FDE,p_desc92_p_O_FDE,p_desc93_p_O_FDE,p_desc94_p_O_FDE,p_desc95_p_O_FDE,p_desc96_p_O_FDE,p_desc97_p_O_FDE,p_desc98_p_O_FDE,p_desc99_p_O_FDE,p_desc100_p_O_FDE,p_desc101_p_O_FDE,p_desc102_p_O_FDE,p_desc103_p_O_FDE,p_desc104_p_O_FDE,p_desc105_p_O_FDE,p_desc106_p_O_FDE,p_desc107_p_O_FDE,p_desc108_p_O_FDE,p_desc109_p_O_FDE,p_desc110_p_O_FDE,p_desc111_p_O_FDE,p_desc112_p_O_FDE,p_desc113_p_O_FDE,p_desc114_p_O_FDE,p_desc115_p_O_FDE,p_desc116_p_O_FDE,p_desc117_p_O_FDE,p_desc118_p_O_FDE,p_desc119_p_O_FDE,p_desc120_p_O_FDE,p_desc121_p_O_FDE,p_desc122_p_O_FDE,p_desc123_p_O_FDE,p_desc124_p_O_FDE,p_desc125_p_O_FDE,p_desc126_p_O_FDE,p_desc127_p_O_FDE,p_desc128_p_O_FDE,p_desc129_p_O_FDE,p_desc130_p_O_FDE,p_desc131_p_O_FDE,p_desc132_p_O_FDE,p_desc133_p_O_FDE,p_desc134_p_O_FDE,p_desc135_p_O_FDE,p_desc136_p_O_FDE,p_desc137_p_O_FDE,p_desc138_p_O_FDE,p_desc139_p_O_FDE,p_desc140_p_O_FDE,p_desc141_p_O_FDE,p_desc142_p_O_FDE,p_desc143_p_O_FDE,p_desc144_p_O_FDE,p_desc145_p_O_FDE,p_desc146_p_O_FDE,p_desc147_p_O_FDE,p_desc148_p_O_FDE,p_desc149_p_O_FDE,p_desc150_p_O_FDE,p_desc151_p_O_FDE,p_desc152_p_O_FDE,p_desc153_p_O_FDE,p_desc154_p_O_FDE,p_desc155_p_O_FDE,p_desc156_p_O_FDE,p_desc157_p_O_FDE,p_desc158_p_O_FDE,p_desc159_p_O_FDE,p_desc160_p_O_FDE,p_desc161_p_O_FDE,p_desc162_p_O_FDE,p_desc163_p_O_FDE,p_desc164_p_O_FDE,p_desc165_p_O_FDE,p_desc166_p_O_FDE,p_desc167_p_O_FDE,p_desc168_p_O_FDE,p_desc169_p_O_FDE,p_desc170_p_O_FDE,p_desc171_p_O_FDE,p_desc172_p_O_FDE,p_desc173_p_O_FDE,p_desc174_p_O_FDE,p_desc175_p_O_FDE,p_desc176_p_O_FDE,p_desc177_p_O_FDE,p_desc178_p_O_FDE,p_desc179_p_O_FDE,p_desc180_p_O_FDE,p_desc181_p_O_FDE,p_desc182_p_O_FDE,p_desc183_p_O_FDE,p_desc184_p_O_FDE,p_desc185_p_O_FDE,p_desc186_p_O_FDE,p_desc187_p_O_FDE,p_desc188_p_O_FDE,p_desc189_p_O_FDE,p_desc190_p_O_FDE,p_desc191_p_O_FDE);
input [1:0] row_sel_R ;
input col_sel_R_mux_i_m3_lut6_2_O6 ;
input col_sel_R_mux_i_m3_lut6_2_O5 ;
input [11:11] single_in_r_R_mux ;
input wr_en_AQ_sel ;
input [1:0] col_sel_R ;
input [1:0] col_sel_R_int ;
output [47:12] out_R_i ;
output [47:0] out_R_r ;
input wr_en_R ;
input N_28_i ;
input clk ;
input N_30_i ;
input N_32_i ;
input N_34_i ;
input N_383_i ;
input N_384_i ;
input N_385_i ;
input N_386_i ;
input N_387_i ;
input N_388_i ;
input N_389_i ;
input N_390_i ;
input N_391_i ;
input N_392_i ;
input N_393_i ;
input N_394_i ;
input N_395_i ;
input N_396_i ;
input N_397_i ;
input N_398_i ;
input N_399_i ;
input N_400_i ;
input N_401_i ;
wire wr_en_R ;
wire N_28_i ;
wire clk ;
wire N_30_i ;
wire N_32_i ;
wire N_34_i ;
wire N_383_i ;
wire N_384_i ;
wire N_385_i ;
wire N_386_i ;
wire N_387_i ;
wire N_388_i ;
wire N_389_i ;
wire N_390_i ;
wire N_391_i ;
wire N_392_i ;
wire N_393_i ;
wire N_394_i ;
wire N_395_i ;
wire N_396_i ;
wire N_397_i ;
wire N_398_i ;
wire N_399_i ;
wire N_400_i ;
wire N_401_i ;
wire [11:0] mat_r_reg_3_3 ;
wire [11:0] mat_r_reg_3_2 ;
wire [11:0] mat_r_reg_3_1 ;
wire [11:0] mat_r_reg_2_2 ;
wire [11:0] mat_r_reg_2_1 ;
wire [11:0] mat_r_reg_1_1 ;
wire [11:0] mat_i_reg_3_2 ;
wire [11:0] mat_i_reg_3_1 ;
wire [11:0] mat_i_reg_3_0 ;
wire [11:0] mat_i_reg_2_1 ;
wire [11:0] mat_i_reg_2_0 ;
wire [11:0] mat_i_reg_1_0 ;
wire VCC ;
wire mat_i_reg_1_0_1_sqmuxa ;
wire mat_i_reg_3_0_1_sqmuxa ;
wire mat_r_reg_1_1_1_sqmuxa ;
wire mat_i_reg_3_1_1_sqmuxa ;
wire mat_i_reg_2_0_1_sqmuxa ;
wire mat_i_reg_3_2_1_sqmuxa ;
wire mat_r_reg_2_2_1_sqmuxa ;
wire mat_r_reg_3_3_1_sqmuxa ;
wire mat_i_reg_2_1_1_sqmuxa ;
wire mat_i_reg_2_1_1_sqmuxa_lut6_2_O5 ;
wire GND ;
input p_desc48_p_O_FDE ;
input p_desc49_p_O_FDE ;
input p_desc50_p_O_FDE ;
input p_desc51_p_O_FDE ;
input p_desc52_p_O_FDE ;
input p_desc53_p_O_FDE ;
input p_desc54_p_O_FDE ;
input p_desc55_p_O_FDE ;
input p_desc56_p_O_FDE ;
input p_desc57_p_O_FDE ;
input p_desc58_p_O_FDE ;
input p_desc59_p_O_FDE ;
input p_desc60_p_O_FDE ;
input p_desc61_p_O_FDE ;
input p_desc62_p_O_FDE ;
input p_desc63_p_O_FDE ;
input p_desc64_p_O_FDE ;
input p_desc65_p_O_FDE ;
input p_desc66_p_O_FDE ;
input p_desc67_p_O_FDE ;
input p_desc68_p_O_FDE ;
input p_desc69_p_O_FDE ;
input p_desc70_p_O_FDE ;
input p_desc71_p_O_FDE ;
input p_desc72_p_O_FDE ;
input p_desc73_p_O_FDE ;
input p_desc74_p_O_FDE ;
input p_desc75_p_O_FDE ;
input p_desc76_p_O_FDE ;
input p_desc77_p_O_FDE ;
input p_desc78_p_O_FDE ;
input p_desc79_p_O_FDE ;
input p_desc80_p_O_FDE ;
input p_desc81_p_O_FDE ;
input p_desc82_p_O_FDE ;
input p_desc83_p_O_FDE ;
input p_desc84_p_O_FDE ;
input p_desc85_p_O_FDE ;
input p_desc86_p_O_FDE ;
input p_desc87_p_O_FDE ;
input p_desc88_p_O_FDE ;
input p_desc89_p_O_FDE ;
input p_desc90_p_O_FDE ;
input p_desc91_p_O_FDE ;
input p_desc92_p_O_FDE ;
input p_desc93_p_O_FDE ;
input p_desc94_p_O_FDE ;
input p_desc95_p_O_FDE ;
input p_desc96_p_O_FDE ;
input p_desc97_p_O_FDE ;
input p_desc98_p_O_FDE ;
input p_desc99_p_O_FDE ;
input p_desc100_p_O_FDE ;
input p_desc101_p_O_FDE ;
input p_desc102_p_O_FDE ;
input p_desc103_p_O_FDE ;
input p_desc104_p_O_FDE ;
input p_desc105_p_O_FDE ;
input p_desc106_p_O_FDE ;
input p_desc107_p_O_FDE ;
input p_desc108_p_O_FDE ;
input p_desc109_p_O_FDE ;
input p_desc110_p_O_FDE ;
input p_desc111_p_O_FDE ;
input p_desc112_p_O_FDE ;
input p_desc113_p_O_FDE ;
input p_desc114_p_O_FDE ;
input p_desc115_p_O_FDE ;
input p_desc116_p_O_FDE ;
input p_desc117_p_O_FDE ;
input p_desc118_p_O_FDE ;
input p_desc119_p_O_FDE ;
input p_desc120_p_O_FDE ;
input p_desc121_p_O_FDE ;
input p_desc122_p_O_FDE ;
input p_desc123_p_O_FDE ;
input p_desc124_p_O_FDE ;
input p_desc125_p_O_FDE ;
input p_desc126_p_O_FDE ;
input p_desc127_p_O_FDE ;
input p_desc128_p_O_FDE ;
input p_desc129_p_O_FDE ;
input p_desc130_p_O_FDE ;
input p_desc131_p_O_FDE ;
input p_desc132_p_O_FDE ;
input p_desc133_p_O_FDE ;
input p_desc134_p_O_FDE ;
input p_desc135_p_O_FDE ;
input p_desc136_p_O_FDE ;
input p_desc137_p_O_FDE ;
input p_desc138_p_O_FDE ;
input p_desc139_p_O_FDE ;
input p_desc140_p_O_FDE ;
input p_desc141_p_O_FDE ;
input p_desc142_p_O_FDE ;
input p_desc143_p_O_FDE ;
input p_desc144_p_O_FDE ;
input p_desc145_p_O_FDE ;
input p_desc146_p_O_FDE ;
input p_desc147_p_O_FDE ;
input p_desc148_p_O_FDE ;
input p_desc149_p_O_FDE ;
input p_desc150_p_O_FDE ;
input p_desc151_p_O_FDE ;
input p_desc152_p_O_FDE ;
input p_desc153_p_O_FDE ;
input p_desc154_p_O_FDE ;
input p_desc155_p_O_FDE ;
input p_desc156_p_O_FDE ;
input p_desc157_p_O_FDE ;
input p_desc158_p_O_FDE ;
input p_desc159_p_O_FDE ;
input p_desc160_p_O_FDE ;
input p_desc161_p_O_FDE ;
input p_desc162_p_O_FDE ;
input p_desc163_p_O_FDE ;
input p_desc164_p_O_FDE ;
input p_desc165_p_O_FDE ;
input p_desc166_p_O_FDE ;
input p_desc167_p_O_FDE ;
input p_desc168_p_O_FDE ;
input p_desc169_p_O_FDE ;
input p_desc170_p_O_FDE ;
input p_desc171_p_O_FDE ;
input p_desc172_p_O_FDE ;
input p_desc173_p_O_FDE ;
input p_desc174_p_O_FDE ;
input p_desc175_p_O_FDE ;
input p_desc176_p_O_FDE ;
input p_desc177_p_O_FDE ;
input p_desc178_p_O_FDE ;
input p_desc179_p_O_FDE ;
input p_desc180_p_O_FDE ;
input p_desc181_p_O_FDE ;
input p_desc182_p_O_FDE ;
input p_desc183_p_O_FDE ;
input p_desc184_p_O_FDE ;
input p_desc185_p_O_FDE ;
input p_desc186_p_O_FDE ;
input p_desc187_p_O_FDE ;
input p_desc188_p_O_FDE ;
input p_desc189_p_O_FDE ;
input p_desc190_p_O_FDE ;
input p_desc191_p_O_FDE ;
// instances
  p_O_FDE desc48(.Q(mat_r_reg_3_3[0:0]),.D(N_28_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc48_p_O_FDE));
  p_O_FDE desc49(.Q(mat_r_reg_3_3[1:1]),.D(N_30_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc49_p_O_FDE));
  p_O_FDE desc50(.Q(mat_r_reg_3_3[2:2]),.D(N_32_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc50_p_O_FDE));
  p_O_FDE desc51(.Q(mat_r_reg_3_3[3:3]),.D(N_34_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc51_p_O_FDE));
  p_O_FDE desc52(.Q(mat_r_reg_3_3[4:4]),.D(N_383_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc52_p_O_FDE));
  p_O_FDE desc53(.Q(mat_r_reg_3_3[5:5]),.D(N_384_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc53_p_O_FDE));
  p_O_FDE desc54(.Q(mat_r_reg_3_3[6:6]),.D(N_385_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc54_p_O_FDE));
  p_O_FDE desc55(.Q(mat_r_reg_3_3[7:7]),.D(N_386_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc55_p_O_FDE));
  p_O_FDE desc56(.Q(mat_r_reg_3_3[8:8]),.D(N_387_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc56_p_O_FDE));
  p_O_FDE desc57(.Q(mat_r_reg_3_3[9:9]),.D(N_388_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc57_p_O_FDE));
  p_O_FDE desc58(.Q(mat_r_reg_3_3[10:10]),.D(N_389_i),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc58_p_O_FDE));
  p_O_FDE desc59(.Q(mat_r_reg_3_3[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_r_reg_3_3_1_sqmuxa),.E(p_desc59_p_O_FDE));
  p_O_FDE desc60(.Q(mat_r_reg_3_2[0:0]),.D(N_28_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc60_p_O_FDE));
  p_O_FDE desc61(.Q(mat_r_reg_3_2[1:1]),.D(N_30_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc61_p_O_FDE));
  p_O_FDE desc62(.Q(mat_r_reg_3_2[2:2]),.D(N_32_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc62_p_O_FDE));
  p_O_FDE desc63(.Q(mat_r_reg_3_2[3:3]),.D(N_34_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc63_p_O_FDE));
  p_O_FDE desc64(.Q(mat_r_reg_3_2[4:4]),.D(N_383_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc64_p_O_FDE));
  p_O_FDE desc65(.Q(mat_r_reg_3_2[5:5]),.D(N_384_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc65_p_O_FDE));
  p_O_FDE desc66(.Q(mat_r_reg_3_2[6:6]),.D(N_385_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc66_p_O_FDE));
  p_O_FDE desc67(.Q(mat_r_reg_3_2[7:7]),.D(N_386_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc67_p_O_FDE));
  p_O_FDE desc68(.Q(mat_r_reg_3_2[8:8]),.D(N_387_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc68_p_O_FDE));
  p_O_FDE desc69(.Q(mat_r_reg_3_2[9:9]),.D(N_388_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc69_p_O_FDE));
  p_O_FDE desc70(.Q(mat_r_reg_3_2[10:10]),.D(N_389_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc70_p_O_FDE));
  p_O_FDE desc71(.Q(mat_r_reg_3_2[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc71_p_O_FDE));
  p_O_FDE desc72(.Q(mat_r_reg_3_1[0:0]),.D(N_28_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc72_p_O_FDE));
  p_O_FDE desc73(.Q(mat_r_reg_3_1[1:1]),.D(N_30_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc73_p_O_FDE));
  p_O_FDE desc74(.Q(mat_r_reg_3_1[2:2]),.D(N_32_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc74_p_O_FDE));
  p_O_FDE desc75(.Q(mat_r_reg_3_1[3:3]),.D(N_34_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc75_p_O_FDE));
  p_O_FDE desc76(.Q(mat_r_reg_3_1[4:4]),.D(N_383_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc76_p_O_FDE));
  p_O_FDE desc77(.Q(mat_r_reg_3_1[5:5]),.D(N_384_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc77_p_O_FDE));
  p_O_FDE desc78(.Q(mat_r_reg_3_1[6:6]),.D(N_385_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc78_p_O_FDE));
  p_O_FDE desc79(.Q(mat_r_reg_3_1[7:7]),.D(N_386_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc79_p_O_FDE));
  p_O_FDE desc80(.Q(mat_r_reg_3_1[8:8]),.D(N_387_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc80_p_O_FDE));
  p_O_FDE desc81(.Q(mat_r_reg_3_1[9:9]),.D(N_388_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc81_p_O_FDE));
  p_O_FDE desc82(.Q(mat_r_reg_3_1[10:10]),.D(N_389_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc82_p_O_FDE));
  p_O_FDE desc83(.Q(mat_r_reg_3_1[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc83_p_O_FDE));
  p_O_FDE desc84(.Q(mat_r_reg_2_2[0:0]),.D(N_28_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc84_p_O_FDE));
  p_O_FDE desc85(.Q(mat_r_reg_2_2[1:1]),.D(N_30_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc85_p_O_FDE));
  p_O_FDE desc86(.Q(mat_r_reg_2_2[2:2]),.D(N_32_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc86_p_O_FDE));
  p_O_FDE desc87(.Q(mat_r_reg_2_2[3:3]),.D(N_34_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc87_p_O_FDE));
  p_O_FDE desc88(.Q(mat_r_reg_2_2[4:4]),.D(N_383_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc88_p_O_FDE));
  p_O_FDE desc89(.Q(mat_r_reg_2_2[5:5]),.D(N_384_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc89_p_O_FDE));
  p_O_FDE desc90(.Q(mat_r_reg_2_2[6:6]),.D(N_385_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc90_p_O_FDE));
  p_O_FDE desc91(.Q(mat_r_reg_2_2[7:7]),.D(N_386_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc91_p_O_FDE));
  p_O_FDE desc92(.Q(mat_r_reg_2_2[8:8]),.D(N_387_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc92_p_O_FDE));
  p_O_FDE desc93(.Q(mat_r_reg_2_2[9:9]),.D(N_388_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc93_p_O_FDE));
  p_O_FDE desc94(.Q(mat_r_reg_2_2[10:10]),.D(N_389_i),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc94_p_O_FDE));
  p_O_FDE desc95(.Q(mat_r_reg_2_2[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_r_reg_2_2_1_sqmuxa),.E(p_desc95_p_O_FDE));
  p_O_FDE desc96(.Q(mat_r_reg_2_1[0:0]),.D(N_28_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc96_p_O_FDE));
  p_O_FDE desc97(.Q(mat_r_reg_2_1[1:1]),.D(N_30_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc97_p_O_FDE));
  p_O_FDE desc98(.Q(mat_r_reg_2_1[2:2]),.D(N_32_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc98_p_O_FDE));
  p_O_FDE desc99(.Q(mat_r_reg_2_1[3:3]),.D(N_34_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc99_p_O_FDE));
  p_O_FDE desc100(.Q(mat_r_reg_2_1[4:4]),.D(N_383_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc100_p_O_FDE));
  p_O_FDE desc101(.Q(mat_r_reg_2_1[5:5]),.D(N_384_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc101_p_O_FDE));
  p_O_FDE desc102(.Q(mat_r_reg_2_1[6:6]),.D(N_385_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc102_p_O_FDE));
  p_O_FDE desc103(.Q(mat_r_reg_2_1[7:7]),.D(N_386_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc103_p_O_FDE));
  p_O_FDE desc104(.Q(mat_r_reg_2_1[8:8]),.D(N_387_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc104_p_O_FDE));
  p_O_FDE desc105(.Q(mat_r_reg_2_1[9:9]),.D(N_388_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc105_p_O_FDE));
  p_O_FDE desc106(.Q(mat_r_reg_2_1[10:10]),.D(N_389_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc106_p_O_FDE));
  p_O_FDE desc107(.Q(mat_r_reg_2_1[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc107_p_O_FDE));
  p_O_FDE desc108(.Q(mat_r_reg_1_1[0:0]),.D(N_28_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc108_p_O_FDE));
  p_O_FDE desc109(.Q(mat_r_reg_1_1[1:1]),.D(N_30_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc109_p_O_FDE));
  p_O_FDE desc110(.Q(mat_r_reg_1_1[2:2]),.D(N_32_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc110_p_O_FDE));
  p_O_FDE desc111(.Q(mat_r_reg_1_1[3:3]),.D(N_34_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc111_p_O_FDE));
  p_O_FDE desc112(.Q(mat_r_reg_1_1[4:4]),.D(N_383_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc112_p_O_FDE));
  p_O_FDE desc113(.Q(mat_r_reg_1_1[5:5]),.D(N_384_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc113_p_O_FDE));
  p_O_FDE desc114(.Q(mat_r_reg_1_1[6:6]),.D(N_385_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc114_p_O_FDE));
  p_O_FDE desc115(.Q(mat_r_reg_1_1[7:7]),.D(N_386_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc115_p_O_FDE));
  p_O_FDE desc116(.Q(mat_r_reg_1_1[8:8]),.D(N_387_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc116_p_O_FDE));
  p_O_FDE desc117(.Q(mat_r_reg_1_1[9:9]),.D(N_388_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc117_p_O_FDE));
  p_O_FDE desc118(.Q(mat_r_reg_1_1[10:10]),.D(N_389_i),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc118_p_O_FDE));
  p_O_FDE desc119(.Q(mat_r_reg_1_1[11:11]),.D(single_in_r_R_mux[11:11]),.C(clk),.CE(mat_r_reg_1_1_1_sqmuxa),.E(p_desc119_p_O_FDE));
  p_O_FDE desc120(.Q(mat_i_reg_3_2[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc120_p_O_FDE));
  p_O_FDE desc121(.Q(mat_i_reg_3_2[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc121_p_O_FDE));
  p_O_FDE desc122(.Q(mat_i_reg_3_2[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc122_p_O_FDE));
  p_O_FDE desc123(.Q(mat_i_reg_3_2[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc123_p_O_FDE));
  p_O_FDE desc124(.Q(mat_i_reg_3_2[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc124_p_O_FDE));
  p_O_FDE desc125(.Q(mat_i_reg_3_2[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc125_p_O_FDE));
  p_O_FDE desc126(.Q(mat_i_reg_3_2[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc126_p_O_FDE));
  p_O_FDE desc127(.Q(mat_i_reg_3_2[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc127_p_O_FDE));
  p_O_FDE desc128(.Q(mat_i_reg_3_2[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc128_p_O_FDE));
  p_O_FDE desc129(.Q(mat_i_reg_3_2[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc129_p_O_FDE));
  p_O_FDE desc130(.Q(mat_i_reg_3_2[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc130_p_O_FDE));
  p_O_FDE desc131(.Q(mat_i_reg_3_2[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_3_2_1_sqmuxa),.E(p_desc131_p_O_FDE));
  p_O_FDE desc132(.Q(mat_i_reg_3_1[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc132_p_O_FDE));
  p_O_FDE desc133(.Q(mat_i_reg_3_1[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc133_p_O_FDE));
  p_O_FDE desc134(.Q(mat_i_reg_3_1[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc134_p_O_FDE));
  p_O_FDE desc135(.Q(mat_i_reg_3_1[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc135_p_O_FDE));
  p_O_FDE desc136(.Q(mat_i_reg_3_1[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc136_p_O_FDE));
  p_O_FDE desc137(.Q(mat_i_reg_3_1[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc137_p_O_FDE));
  p_O_FDE desc138(.Q(mat_i_reg_3_1[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc138_p_O_FDE));
  p_O_FDE desc139(.Q(mat_i_reg_3_1[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc139_p_O_FDE));
  p_O_FDE desc140(.Q(mat_i_reg_3_1[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc140_p_O_FDE));
  p_O_FDE desc141(.Q(mat_i_reg_3_1[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc141_p_O_FDE));
  p_O_FDE desc142(.Q(mat_i_reg_3_1[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc142_p_O_FDE));
  p_O_FDE desc143(.Q(mat_i_reg_3_1[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_3_1_1_sqmuxa),.E(p_desc143_p_O_FDE));
  p_O_FDE desc144(.Q(mat_i_reg_3_0[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc144_p_O_FDE));
  p_O_FDE desc145(.Q(mat_i_reg_3_0[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc145_p_O_FDE));
  p_O_FDE desc146(.Q(mat_i_reg_3_0[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc146_p_O_FDE));
  p_O_FDE desc147(.Q(mat_i_reg_3_0[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc147_p_O_FDE));
  p_O_FDE desc148(.Q(mat_i_reg_3_0[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc148_p_O_FDE));
  p_O_FDE desc149(.Q(mat_i_reg_3_0[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc149_p_O_FDE));
  p_O_FDE desc150(.Q(mat_i_reg_3_0[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc150_p_O_FDE));
  p_O_FDE desc151(.Q(mat_i_reg_3_0[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc151_p_O_FDE));
  p_O_FDE desc152(.Q(mat_i_reg_3_0[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc152_p_O_FDE));
  p_O_FDE desc153(.Q(mat_i_reg_3_0[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc153_p_O_FDE));
  p_O_FDE desc154(.Q(mat_i_reg_3_0[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc154_p_O_FDE));
  p_O_FDE desc155(.Q(mat_i_reg_3_0[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_3_0_1_sqmuxa),.E(p_desc155_p_O_FDE));
  p_O_FDE desc156(.Q(mat_i_reg_2_1[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc156_p_O_FDE));
  p_O_FDE desc157(.Q(mat_i_reg_2_1[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc157_p_O_FDE));
  p_O_FDE desc158(.Q(mat_i_reg_2_1[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc158_p_O_FDE));
  p_O_FDE desc159(.Q(mat_i_reg_2_1[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc159_p_O_FDE));
  p_O_FDE desc160(.Q(mat_i_reg_2_1[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc160_p_O_FDE));
  p_O_FDE desc161(.Q(mat_i_reg_2_1[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc161_p_O_FDE));
  p_O_FDE desc162(.Q(mat_i_reg_2_1[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc162_p_O_FDE));
  p_O_FDE desc163(.Q(mat_i_reg_2_1[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc163_p_O_FDE));
  p_O_FDE desc164(.Q(mat_i_reg_2_1[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc164_p_O_FDE));
  p_O_FDE desc165(.Q(mat_i_reg_2_1[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc165_p_O_FDE));
  p_O_FDE desc166(.Q(mat_i_reg_2_1[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc166_p_O_FDE));
  p_O_FDE desc167(.Q(mat_i_reg_2_1[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_2_1_1_sqmuxa),.E(p_desc167_p_O_FDE));
  p_O_FDE desc168(.Q(mat_i_reg_2_0[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc168_p_O_FDE));
  p_O_FDE desc169(.Q(mat_i_reg_2_0[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc169_p_O_FDE));
  p_O_FDE desc170(.Q(mat_i_reg_2_0[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc170_p_O_FDE));
  p_O_FDE desc171(.Q(mat_i_reg_2_0[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc171_p_O_FDE));
  p_O_FDE desc172(.Q(mat_i_reg_2_0[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc172_p_O_FDE));
  p_O_FDE desc173(.Q(mat_i_reg_2_0[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc173_p_O_FDE));
  p_O_FDE desc174(.Q(mat_i_reg_2_0[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc174_p_O_FDE));
  p_O_FDE desc175(.Q(mat_i_reg_2_0[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc175_p_O_FDE));
  p_O_FDE desc176(.Q(mat_i_reg_2_0[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc176_p_O_FDE));
  p_O_FDE desc177(.Q(mat_i_reg_2_0[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc177_p_O_FDE));
  p_O_FDE desc178(.Q(mat_i_reg_2_0[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc178_p_O_FDE));
  p_O_FDE desc179(.Q(mat_i_reg_2_0[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_2_0_1_sqmuxa),.E(p_desc179_p_O_FDE));
  p_O_FDE desc180(.Q(mat_i_reg_1_0[0:0]),.D(N_390_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc180_p_O_FDE));
  p_O_FDE desc181(.Q(mat_i_reg_1_0[1:1]),.D(N_391_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc181_p_O_FDE));
  p_O_FDE desc182(.Q(mat_i_reg_1_0[2:2]),.D(N_392_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc182_p_O_FDE));
  p_O_FDE desc183(.Q(mat_i_reg_1_0[3:3]),.D(N_393_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc183_p_O_FDE));
  p_O_FDE desc184(.Q(mat_i_reg_1_0[4:4]),.D(N_394_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc184_p_O_FDE));
  p_O_FDE desc185(.Q(mat_i_reg_1_0[5:5]),.D(N_395_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc185_p_O_FDE));
  p_O_FDE desc186(.Q(mat_i_reg_1_0[6:6]),.D(N_396_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc186_p_O_FDE));
  p_O_FDE desc187(.Q(mat_i_reg_1_0[7:7]),.D(N_397_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc187_p_O_FDE));
  p_O_FDE desc188(.Q(mat_i_reg_1_0[8:8]),.D(N_398_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc188_p_O_FDE));
  p_O_FDE desc189(.Q(mat_i_reg_1_0[9:9]),.D(N_399_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc189_p_O_FDE));
  p_O_FDE desc190(.Q(mat_i_reg_1_0[10:10]),.D(N_400_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc190_p_O_FDE));
  p_O_FDE desc191(.Q(mat_i_reg_1_0[11:11]),.D(N_401_i),.C(clk),.CE(mat_i_reg_1_0_1_sqmuxa),.E(p_desc191_p_O_FDE));
  LUT6 desc192(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[0:0]),.I3(mat_r_reg_3_2[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[12:12]));
defparam desc192.INIT=64'hFC300000A820A820;
  LUT6 desc193(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[11:11]),.I3(mat_i_reg_3_1[11:11]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[35:35]));
defparam desc193.INIT=64'hFC300000A820A820;
  LUT6 desc194(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[10:10]),.I3(mat_i_reg_3_1[10:10]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[34:34]));
defparam desc194.INIT=64'hFC300000A820A820;
  LUT6 desc195(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[9:9]),.I3(mat_i_reg_3_1[9:9]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[33:33]));
defparam desc195.INIT=64'hFC300000A820A820;
  LUT6 desc196(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[6:6]),.I3(mat_i_reg_3_1[6:6]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[30:30]));
defparam desc196.INIT=64'hFC300000A820A820;
  LUT6 desc197(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[5:5]),.I3(mat_i_reg_3_1[5:5]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[29:29]));
defparam desc197.INIT=64'hFC300000A820A820;
  LUT6 desc198(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[4:4]),.I3(mat_i_reg_3_1[4:4]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[28:28]));
defparam desc198.INIT=64'hFC300000A820A820;
  LUT6 desc199(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[3:3]),.I3(mat_i_reg_3_1[3:3]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[27:27]));
defparam desc199.INIT=64'hFC300000A820A820;
  LUT6 desc200(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[2:2]),.I3(mat_i_reg_3_1[2:2]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[26:26]));
defparam desc200.INIT=64'hFC300000A820A820;
  LUT6 desc201(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[1:1]),.I3(mat_i_reg_3_1[1:1]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[25:25]));
defparam desc201.INIT=64'hFC300000A820A820;
  LUT6 desc202(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[0:0]),.I3(mat_i_reg_3_1[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[24:24]));
defparam desc202.INIT=64'hFC300000A820A820;
  LUT6 desc203(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[1:1]),.I3(mat_r_reg_3_2[1:1]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[13:13]));
defparam desc203.INIT=64'hFC300000A820A820;
  LUT6 desc204(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[3:3]),.I3(mat_r_reg_3_2[3:3]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[15:15]));
defparam desc204.INIT=64'hFC300000A820A820;
  LUT6 desc205(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[2:2]),.I3(mat_r_reg_3_2[2:2]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[14:14]));
defparam desc205.INIT=64'hFC300000A820A820;
  LUT6 desc206(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[5:5]),.I3(mat_r_reg_3_2[5:5]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[17:17]));
defparam desc206.INIT=64'hFC300000A820A820;
  LUT6 desc207(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[7:7]),.I3(mat_r_reg_3_2[7:7]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[19:19]));
defparam desc207.INIT=64'hFC300000A820A820;
  LUT6 desc208(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[6:6]),.I3(mat_r_reg_3_2[6:6]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[18:18]));
defparam desc208.INIT=64'hFC300000A820A820;
  LUT6 desc209(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[9:9]),.I3(mat_r_reg_3_2[9:9]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[21:21]));
defparam desc209.INIT=64'hFC300000A820A820;
  LUT6 desc210(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[8:8]),.I3(mat_r_reg_3_2[8:8]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[20:20]));
defparam desc210.INIT=64'hFC300000A820A820;
  LUT6 desc211(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[11:11]),.I3(mat_r_reg_3_2[11:11]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[23:23]));
defparam desc211.INIT=64'hFC300000A820A820;
  LUT6 desc212(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[10:10]),.I3(mat_r_reg_3_2[10:10]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[22:22]));
defparam desc212.INIT=64'hFC300000A820A820;
  LUT6 desc213(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[7:7]),.I3(mat_i_reg_3_1[7:7]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[31:31]));
defparam desc213.INIT=64'hFC300000A820A820;
  LUT6 desc214(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_r_reg_2_2[4:4]),.I3(mat_r_reg_3_2[4:4]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[16:16]));
defparam desc214.INIT=64'hFC300000A820A820;
  LUT6 desc215(.I0(col_sel_R[1:1]),.I1(col_sel_R_mux_i_m3_lut6_2_O6),.I2(mat_i_reg_2_1[8:8]),.I3(mat_i_reg_3_1[8:8]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[32:32]));
defparam desc215.INIT=64'hFC300000A820A820;
  LUT6 desc216(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[4:4]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[4:4]));
defparam desc216.INIT=64'hF000000080808080;
  LUT6 desc217(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[3:3]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[3:3]));
defparam desc217.INIT=64'hF000000080808080;
  LUT6 desc218(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[1:1]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[1:1]));
defparam desc218.INIT=64'hF000000080808080;
  LUT6 desc219(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[0:0]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[0:0]));
defparam desc219.INIT=64'hF000000080808080;
  LUT6 desc220(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[11:11]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[23:23]));
defparam desc220.INIT=64'hF000000080808080;
  LUT6 desc221(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[10:10]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[22:22]));
defparam desc221.INIT=64'hF000000080808080;
  LUT6 desc222(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[9:9]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[21:21]));
defparam desc222.INIT=64'hF000000080808080;
  LUT6 desc223(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[8:8]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[8:8]));
defparam desc223.INIT=64'hF000000080808080;
  LUT6 desc224(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[10:10]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[10:10]));
defparam desc224.INIT=64'hF000000080808080;
  LUT6 desc225(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[9:9]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[9:9]));
defparam desc225.INIT=64'hF000000080808080;
  LUT6 desc226(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[7:7]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[7:7]));
defparam desc226.INIT=64'hF000000080808080;
  LUT6 desc227(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[6:6]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[6:6]));
defparam desc227.INIT=64'hF000000080808080;
  LUT6 desc228(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[5:5]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[5:5]));
defparam desc228.INIT=64'hF000000080808080;
  LUT6 desc229(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[2:2]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[14:14]));
defparam desc229.INIT=64'hF000000080808080;
  LUT6 desc230(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[2:2]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[2:2]));
defparam desc230.INIT=64'hF000000080808080;
  LUT6 desc231(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[8:8]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[20:20]));
defparam desc231.INIT=64'hF000000080808080;
  LUT6 desc232(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[7:7]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[19:19]));
defparam desc232.INIT=64'hF000000080808080;
  LUT6 desc233(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[6:6]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[18:18]));
defparam desc233.INIT=64'hF000000080808080;
  LUT6 desc234(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[5:5]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[17:17]));
defparam desc234.INIT=64'hF000000080808080;
  LUT6 desc235(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[4:4]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[16:16]));
defparam desc235.INIT=64'hF000000080808080;
  LUT6 desc236(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[3:3]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[15:15]));
defparam desc236.INIT=64'hF000000080808080;
  LUT6 desc237(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[1:1]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[13:13]));
defparam desc237.INIT=64'hF000000080808080;
  LUT6 desc238(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_i_reg_3_2[0:0]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_i[12:12]));
defparam desc238.INIT=64'hF000000080808080;
  LUT6 desc239(.I0(col_sel_R[0:0]),.I1(col_sel_R[1:1]),.I2(mat_r_reg_3_3[11:11]),.I3(col_sel_R_int[0:0]),.I4(col_sel_R_int[1:1]),.I5(wr_en_AQ_sel),.O(out_R_r[11:11]));
defparam desc239.INIT=64'hF000000080808080;
  LUT5 desc240(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[2:2]),.I3(mat_i_reg_2_0[2:2]),.I4(mat_i_reg_3_0[2:2]),.O(out_R_i[38:38]));
defparam desc240.INIT=32'hECA86420;
  LUT5 desc241(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[1:1]),.I3(mat_i_reg_2_0[1:1]),.I4(mat_i_reg_3_0[1:1]),.O(out_R_i[37:37]));
defparam desc241.INIT=32'hECA86420;
  LUT5 desc242(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[4:4]),.I3(mat_i_reg_2_0[4:4]),.I4(mat_i_reg_3_0[4:4]),.O(out_R_i[40:40]));
defparam desc242.INIT=32'hECA86420;
  LUT5 desc243(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[3:3]),.I3(mat_i_reg_2_0[3:3]),.I4(mat_i_reg_3_0[3:3]),.O(out_R_i[39:39]));
defparam desc243.INIT=32'hECA86420;
  LUT5 desc244(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[6:6]),.I3(mat_i_reg_2_0[6:6]),.I4(mat_i_reg_3_0[6:6]),.O(out_R_i[42:42]));
defparam desc244.INIT=32'hECA86420;
  LUT5 desc245(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[5:5]),.I3(mat_i_reg_2_0[5:5]),.I4(mat_i_reg_3_0[5:5]),.O(out_R_i[41:41]));
defparam desc245.INIT=32'hECA86420;
  LUT5 desc246(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[8:8]),.I3(mat_i_reg_2_0[8:8]),.I4(mat_i_reg_3_0[8:8]),.O(out_R_i[44:44]));
defparam desc246.INIT=32'hECA86420;
  LUT5 desc247(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[7:7]),.I3(mat_i_reg_2_0[7:7]),.I4(mat_i_reg_3_0[7:7]),.O(out_R_i[43:43]));
defparam desc247.INIT=32'hECA86420;
  LUT5 desc248(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[10:10]),.I3(mat_i_reg_2_0[10:10]),.I4(mat_i_reg_3_0[10:10]),.O(out_R_i[46:46]));
defparam desc248.INIT=32'hECA86420;
  LUT5 desc249(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[9:9]),.I3(mat_i_reg_2_0[9:9]),.I4(mat_i_reg_3_0[9:9]),.O(out_R_i[45:45]));
defparam desc249.INIT=32'hECA86420;
  LUT5 desc250(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[11:11]),.I3(mat_i_reg_2_0[11:11]),.I4(mat_i_reg_3_0[11:11]),.O(out_R_i[47:47]));
defparam desc250.INIT=32'hECA86420;
  LUT5 desc251(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[11:11]),.I3(mat_r_reg_2_1[11:11]),.I4(mat_r_reg_3_1[11:11]),.O(out_R_r[35:35]));
defparam desc251.INIT=32'hECA86420;
  LUT5 desc252(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[8:8]),.I3(mat_r_reg_2_1[8:8]),.I4(mat_r_reg_3_1[8:8]),.O(out_R_r[32:32]));
defparam desc252.INIT=32'hECA86420;
  LUT5 desc253(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[9:9]),.I3(mat_r_reg_2_1[9:9]),.I4(mat_r_reg_3_1[9:9]),.O(out_R_r[33:33]));
defparam desc253.INIT=32'hECA86420;
  LUT5 desc254(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[10:10]),.I3(mat_r_reg_2_1[10:10]),.I4(mat_r_reg_3_1[10:10]),.O(out_R_r[34:34]));
defparam desc254.INIT=32'hECA86420;
  LUT5 desc255(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[5:5]),.I3(mat_r_reg_2_1[5:5]),.I4(mat_r_reg_3_1[5:5]),.O(out_R_r[29:29]));
defparam desc255.INIT=32'hECA86420;
  LUT5 desc256(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[6:6]),.I3(mat_r_reg_2_1[6:6]),.I4(mat_r_reg_3_1[6:6]),.O(out_R_r[30:30]));
defparam desc256.INIT=32'hECA86420;
  LUT5 desc257(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[7:7]),.I3(mat_r_reg_2_1[7:7]),.I4(mat_r_reg_3_1[7:7]),.O(out_R_r[31:31]));
defparam desc257.INIT=32'hECA86420;
  LUT5 desc258(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[2:2]),.I3(mat_r_reg_2_1[2:2]),.I4(mat_r_reg_3_1[2:2]),.O(out_R_r[26:26]));
defparam desc258.INIT=32'hECA86420;
  LUT5 desc259(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[3:3]),.I3(mat_r_reg_2_1[3:3]),.I4(mat_r_reg_3_1[3:3]),.O(out_R_r[27:27]));
defparam desc259.INIT=32'hECA86420;
  LUT5 desc260(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[4:4]),.I3(mat_r_reg_2_1[4:4]),.I4(mat_r_reg_3_1[4:4]),.O(out_R_r[28:28]));
defparam desc260.INIT=32'hECA86420;
  LUT5 desc261(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_i_reg_1_0[0:0]),.I3(mat_i_reg_2_0[0:0]),.I4(mat_i_reg_3_0[0:0]),.O(out_R_i[36:36]));
defparam desc261.INIT=32'hECA86420;
  LUT5 desc262(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[0:0]),.I3(mat_r_reg_2_1[0:0]),.I4(mat_r_reg_3_1[0:0]),.O(out_R_r[24:24]));
defparam desc262.INIT=32'hECA86420;
  LUT5 desc263(.I0(col_sel_R_mux_i_m3_lut6_2_O6),.I1(col_sel_R_mux_i_m3_lut6_2_O5),.I2(mat_r_reg_1_1[1:1]),.I3(mat_r_reg_2_1[1:1]),.I4(mat_r_reg_3_1[1:1]),.O(out_R_r[25:25]));
defparam desc263.INIT=32'hECA86420;
  RAM32X1S mat_r_reg_0_mat_r_reg_0_11_0(.O(out_R_r[47:47]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(single_in_r_R_mux[11:11]),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_10_0(.O(out_R_r[46:46]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_389_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_9_0(.O(out_R_r[45:45]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_388_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_8_0(.O(out_R_r[44:44]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_387_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_7_0(.O(out_R_r[43:43]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_386_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_6_0(.O(out_R_r[42:42]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_385_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_5_0(.O(out_R_r[41:41]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_384_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_4_0(.O(out_R_r[40:40]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_383_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_3_0(.O(out_R_r[39:39]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_34_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_2_0(.O(out_R_r[38:38]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_32_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_1_0(.O(out_R_r[37:37]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_30_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  RAM32X1S mat_r_reg_0_mat_r_reg_0_0_0(.O(out_R_r[36:36]),.A0(col_sel_R_mux_i_m3_lut6_2_O6),.A1(col_sel_R_mux_i_m3_lut6_2_O5),.A2(GND),.A3(GND),.A4(GND),.D(N_28_i),.WCLK(clk),.WE(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT5 mat_i_reg_2_1_1_sqmuxa_lut6_2_o6(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_2_1_1_sqmuxa));
defparam mat_i_reg_2_1_1_sqmuxa_lut6_2_o6.INIT=32'h00200000;
  LUT3 mat_i_reg_2_1_1_sqmuxa_lut6_2_o5(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.O(mat_i_reg_2_1_1_sqmuxa_lut6_2_O5));
defparam mat_i_reg_2_1_1_sqmuxa_lut6_2_o5.INIT=8'h10;
  LUT5 mat_r_reg_2_2_1_sqmuxa_lut6_2_o6(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_r_reg_2_2_1_sqmuxa));
defparam mat_r_reg_2_2_1_sqmuxa_lut6_2_o6.INIT=32'h00400000;
  LUT5 mat_r_reg_2_2_1_sqmuxa_lut6_2_o5(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_r_reg_3_3_1_sqmuxa));
defparam mat_r_reg_2_2_1_sqmuxa_lut6_2_o5.INIT=32'h80000000;
  LUT5 mat_i_reg_2_0_1_sqmuxa_lut6_2_o6(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_2_0_1_sqmuxa));
defparam mat_i_reg_2_0_1_sqmuxa_lut6_2_o6.INIT=32'h00100000;
  LUT5 mat_i_reg_2_0_1_sqmuxa_lut6_2_o5(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_3_2_1_sqmuxa));
defparam mat_i_reg_2_0_1_sqmuxa_lut6_2_o5.INIT=32'h40000000;
  LUT5 mat_r_reg_1_1_1_sqmuxa_lut6_2_o6(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_r_reg_1_1_1_sqmuxa));
defparam mat_r_reg_1_1_1_sqmuxa_lut6_2_o6.INIT=32'h00002000;
  LUT5 mat_r_reg_1_1_1_sqmuxa_lut6_2_o5(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_3_1_1_sqmuxa));
defparam mat_r_reg_1_1_1_sqmuxa_lut6_2_o5.INIT=32'h20000000;
  LUT5 mat_i_reg_1_0_1_sqmuxa_lut6_2_o6(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_1_0_1_sqmuxa));
defparam mat_i_reg_1_0_1_sqmuxa_lut6_2_o6.INIT=32'h00001000;
  LUT5 mat_i_reg_1_0_1_sqmuxa_lut6_2_o5(.I0(row_sel_R[0:0]),.I1(row_sel_R[1:1]),.I2(wr_en_R),.I3(col_sel_R_mux_i_m3_lut6_2_O6),.I4(col_sel_R_mux_i_m3_lut6_2_O5),.O(mat_i_reg_3_0_1_sqmuxa));
defparam mat_i_reg_1_0_1_sqmuxa_lut6_2_o5.INIT=32'h10000000;
endmodule
module shifterZ0_inj (input_reg,shift_amount_1,un14_pos_output,ret_val,un11_output_6_d_0,out_shift_amount,un7_output_2_0_0,un7_output_2_1,output_d,shift_amount_1_i,un11_output_1,un11_output_2,un20_output_2,pre_output,done_inv_sqrt,un4_overflow_0,output_reg_pipe_12_RNIPJ901_O6,un9_0_axb_8,un9_0_s_6,un9_0_s_7,N_414,N_33,clk,N_420,un3_shift_right,N_410,un9_0_s_5,un9_0_s_8,N_79,N_50,un9_0_s_4,un9_0_s_3,N_13_0,N_100_i,N_31,N_18_0,N_378,N_33_0,N_80,N_51,un9_0_s_0,un9_0_s_1,m9_0_0,N_417,N_62,N_454,SUM1_0_i_1_1,N_56,N_434_i,N_431_i,N_428_i,N_425_i,un9_0_s_2,N_419,N_49,N_413,un20_output_0_0_a2_0_0_lut6_2_O5,un1_apply_nrlt8_1,un1_apply_nrlt7,p_output_reg_pipe_13_Z_p_O_FD,p_output_reg_pipe_12_Z_p_O_FD,p_output_reg_pipe_Z_p_O_FD,p_output_reg_pipe_1_Z_p_O_FDE,p_output_reg_pipe_4_Z_p_O_FDE,p_output_reg_pipe_5_Z_p_O_FDE,p_output_reg_pipe_6_Z_p_O_FDE,p_output_reg_pipe_9_Z_p_O_FDE,p_output_reg_pipe_10_Z_p_O_FDE,p_output_reg_pipe_11_Z_p_O_FDE,p_output_reg_pipe_14_Z_p_O_FDE,p_output_reg_pipe_15_Z_p_O_FDE,p_output_reg_pipe_16_Z_p_O_FDE,p_output_reg_pipe_19_Z_p_O_FDE);
input [11:10] input_reg ;
input [1:1] shift_amount_1 ;
input [6:3] un14_pos_output ;
input [3:1] ret_val ;
output [9:9] un11_output_6_d_0 ;
input [1:1] out_shift_amount ;
output [6:6] un7_output_2_0_0 ;
output [6:5] un7_output_2_1 ;
output [4:4] output_d ;
input [2:2] shift_amount_1_i ;
output un11_output_1 ;
output un11_output_2 ;
input [14:14] un20_output_2 ;
output [11:1] pre_output ;
input done_inv_sqrt ;
input un4_overflow_0 ;
output output_reg_pipe_12_RNIPJ901_O6 ;
input un9_0_axb_8 ;
input un9_0_s_6 ;
input un9_0_s_7 ;
output N_414 ;
output N_33 ;
input clk ;
output N_420 ;
input un3_shift_right ;
output N_410 ;
input un9_0_s_5 ;
input un9_0_s_8 ;
output N_79 ;
output N_50 ;
input un9_0_s_4 ;
input un9_0_s_3 ;
output N_13_0 ;
input N_100_i ;
output N_31 ;
output N_18_0 ;
input N_378 ;
output N_33_0 ;
output N_80 ;
output N_51 ;
input un9_0_s_0 ;
input un9_0_s_1 ;
output m9_0_0 ;
output N_417 ;
output N_62 ;
input N_454 ;
input SUM1_0_i_1_1 ;
output N_56 ;
output N_434_i ;
output N_431_i ;
output N_428_i ;
output N_425_i ;
input un9_0_s_2 ;
input N_419 ;
output N_49 ;
output N_413 ;
input un20_output_0_0_a2_0_0_lut6_2_O5 ;
input un1_apply_nrlt8_1 ;
input un1_apply_nrlt7 ;
wire un11_output_1 ;
wire un11_output_2 ;
wire done_inv_sqrt ;
wire un4_overflow_0 ;
wire output_reg_pipe_12_RNIPJ901_O6 ;
wire un9_0_axb_8 ;
wire un9_0_s_6 ;
wire un9_0_s_7 ;
wire N_414 ;
wire N_33 ;
wire clk ;
wire N_420 ;
wire un3_shift_right ;
wire N_410 ;
wire un9_0_s_5 ;
wire un9_0_s_8 ;
wire N_79 ;
wire N_50 ;
wire un9_0_s_4 ;
wire un9_0_s_3 ;
wire N_13_0 ;
wire N_100_i ;
wire N_31 ;
wire N_18_0 ;
wire N_378 ;
wire N_33_0 ;
wire N_80 ;
wire N_51 ;
wire un9_0_s_0 ;
wire un9_0_s_1 ;
wire m9_0_0 ;
wire N_417 ;
wire N_62 ;
wire N_454 ;
wire SUM1_0_i_1_1 ;
wire N_56 ;
wire N_434_i ;
wire N_431_i ;
wire N_428_i ;
wire N_425_i ;
wire un9_0_s_2 ;
wire N_419 ;
wire N_49 ;
wire N_413 ;
wire un20_output_0_0_a2_0_0_lut6_2_O5 ;
wire un1_apply_nrlt8_1 ;
wire un1_apply_nrlt7 ;
wire [6:3] un14_pos_outputf ;
wire [6:3] pre_outputf ;
wire [4:4] un11_output ;
wire [6:4] un11_output_1_Z ;
wire un4_overflow_if ;
wire VCC ;
wire un4_overflow_i_0 ;
wire output_reg_pipe_13 ;
wire m41 ;
wire output_reg_pipe ;
wire m44 ;
wire output_reg_pipe_5 ;
wire N_427 ;
wire output_reg_pipe_10 ;
wire N_430 ;
wire output_reg_pipe_15 ;
wire N_433 ;
wire m25_0_1 ;
wire m25_0_0 ;
wire m17_0_2 ;
wire GND ;
input p_output_reg_pipe_13_Z_p_O_FD ;
input p_output_reg_pipe_12_Z_p_O_FD ;
input p_output_reg_pipe_Z_p_O_FD ;
input p_output_reg_pipe_1_Z_p_O_FDE ;
input p_output_reg_pipe_4_Z_p_O_FDE ;
input p_output_reg_pipe_5_Z_p_O_FDE ;
input p_output_reg_pipe_6_Z_p_O_FDE ;
input p_output_reg_pipe_9_Z_p_O_FDE ;
input p_output_reg_pipe_10_Z_p_O_FDE ;
input p_output_reg_pipe_11_Z_p_O_FDE ;
input p_output_reg_pipe_14_Z_p_O_FDE ;
input p_output_reg_pipe_15_Z_p_O_FDE ;
input p_output_reg_pipe_16_Z_p_O_FDE ;
input p_output_reg_pipe_19_Z_p_O_FDE ;
// instances
  p_O_FD output_reg_pipe_13_Z(.Q(output_reg_pipe_13),.D(m41),.C(clk),.E(p_output_reg_pipe_13_Z_p_O_FD));
  p_O_FD output_reg_pipe_12_Z(.Q(un4_overflow_if),.D(un4_overflow_i_0),.C(clk),.E(p_output_reg_pipe_12_Z_p_O_FD));
  p_O_FD output_reg_pipe_Z(.Q(output_reg_pipe),.D(m44),.C(clk),.E(p_output_reg_pipe_Z_p_O_FD));
  LUT5 output_reg_pipe_RNO(.I0(un4_overflow_0),.I1(pre_output[3:3]),.I2(N_420),.I3(output_reg_pipe),.I4(done_inv_sqrt),.O(m44));
defparam output_reg_pipe_RNO.INIT=32'h0101FF00;
  LUT6 output_reg_pipe_13_RNO(.I0(input_reg[10:10]),.I1(input_reg[11:11]),.I2(un4_overflow_0),.I3(N_420),.I4(output_reg_pipe_13),.I5(done_inv_sqrt),.O(m41));
defparam output_reg_pipe_13_RNO.INIT=64'hEF00EF00FFFF0000;
  p_O_FDE output_reg_pipe_1_Z(.Q(un14_pos_outputf[3:3]),.D(un14_pos_output[3:3]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_1_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_4_Z(.Q(pre_outputf[3:3]),.D(pre_output[3:3]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_4_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_5_Z(.Q(output_reg_pipe_5),.D(N_427),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_5_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_6_Z(.Q(un14_pos_outputf[4:4]),.D(un14_pos_output[4:4]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_6_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_9_Z(.Q(pre_outputf[4:4]),.D(pre_output[4:4]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_9_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_10_Z(.Q(output_reg_pipe_10),.D(N_430),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_10_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_11_Z(.Q(un14_pos_outputf[5:5]),.D(un14_pos_output[5:5]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_11_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_14_Z(.Q(pre_outputf[5:5]),.D(pre_output[5:5]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_14_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_15_Z(.Q(output_reg_pipe_15),.D(N_433),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_15_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_16_Z(.Q(un14_pos_outputf[6:6]),.D(un14_pos_output[6:6]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_16_Z_p_O_FDE));
  p_O_FDE output_reg_pipe_19_Z(.Q(pre_outputf[6:6]),.D(pre_output[6:6]),.C(clk),.CE(done_inv_sqrt),.E(p_output_reg_pipe_19_Z_p_O_FDE));
  LUT3 desc883(.I0(un3_shift_right),.I1(un7_output_2_1[5:5]),.I2(un11_output_1),.O(pre_output[5:5]));
defparam desc883.INIT=8'hD8;
  LUT4 m26(.I0(ret_val[3:3]),.I1(N_410),.I2(m25_0_1),.I3(m25_0_0),.O(pre_output[8:8]));
defparam m26.INIT=16'hFFD8;
  LUT5 desc884(.I0(ret_val[3:3]),.I1(ret_val[1:1]),.I2(shift_amount_1[1:1]),.I3(un9_0_s_5),.I4(un9_0_s_8),.O(un11_output_6_d_0[9:9]));
defparam desc884.INIT=32'hF8F00800;
  LUT5 desc885(.I0(ret_val[3:3]),.I1(ret_val[1:1]),.I2(un3_shift_right),.I3(N_79),.I4(N_50),.O(pre_output[2:2]));
defparam desc885.INIT=32'hFFF00700;
  LUT4 m19(.I0(ret_val[2:2]),.I1(un9_0_axb_8),.I2(shift_amount_1[1:1]),.I3(un9_0_s_4),.O(N_410));
defparam m19.INIT=16'h0600;
  LUT4 m12(.I0(ret_val[2:2]),.I1(un9_0_axb_8),.I2(shift_amount_1[1:1]),.I3(un9_0_s_3),.O(N_13_0));
defparam m12.INIT=16'h0600;
  LUT3 m31(.I0(N_100_i),.I1(un9_0_s_6),.I2(N_31),.O(pre_output[10:10]));
defparam m31.INIT=8'hE4;
  LUT3 m18(.I0(N_100_i),.I1(un9_0_s_3),.I2(N_18_0),.O(pre_output[7:7]));
defparam m18.INIT=8'hE4;
  LUT5 desc886(.I0(N_378),.I1(un3_shift_right),.I2(un9_0_s_6),.I3(N_33_0),.I4(un11_output[4:4]),.O(pre_output[4:4]));
defparam desc886.INIT=32'hF733CC80;
  LUT5 desc887(.I0(ret_val[3:3]),.I1(ret_val[1:1]),.I2(un9_0_axb_8),.I3(out_shift_amount[1:1]),.I4(un9_0_s_8),.O(un7_output_2_0_0[6:6]));
defparam desc887.INIT=32'h437F007F;
  LUT6 desc888(.I0(ret_val[3:3]),.I1(ret_val[1:1]),.I2(un9_0_axb_8),.I3(un3_shift_right),.I4(N_80),.I5(N_51),.O(pre_output[3:3]));
defparam desc888.INIT=64'hFF7FFF00007F0000;
  LUT6 m25_0_1_cZ(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un3_shift_right),.I4(un9_0_s_8),.I5(un9_0_s_7),.O(m25_0_1));
defparam m25_0_1_cZ.INIT=64'h090F000609090000;
  LUT6 m30(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un3_shift_right),.I4(un9_0_s_8),.I5(un9_0_s_7),.O(N_31));
defparam m30.INIT=64'h00F0006000900000;
  LUT5 desc889(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un9_0_s_6),.I4(un9_0_s_7),.O(un7_output_2_1[5:5]));
defparam desc889.INIT=32'hFF990F09;
  LUT5 desc890(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un9_0_s_6),.I4(un9_0_s_7),.O(un7_output_2_1[6:6]));
defparam desc890.INIT=32'hFFF69990;
  LUT6 m25_0_0_cZ(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un3_shift_right),.I4(un9_0_s_5),.I5(un9_0_s_6),.O(m25_0_0));
defparam m25_0_0_cZ.INIT=64'h00F0009000600000;
  LUT5 desc891(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(un3_shift_right),.I3(un9_0_s_6),.I4(un11_output[4:4]),.O(output_d[4:4]));
defparam desc891.INIT=32'h9F0F9000;
  LUT6 m9_0_0_c(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(out_shift_amount[1:1]),.I3(un3_shift_right),.I4(un9_0_s_0),.I5(un9_0_s_1),.O(m9_0_0));
defparam m9_0_0_c.INIT=64'h0F09060009090000;
  LUT4 m33(.I0(ret_val[2:2]),.I1(shift_amount_1[1:1]),.I2(un3_shift_right),.I3(un9_0_s_8),.O(N_417));
defparam m33.INIT=16'h0400;
  LUT4 desc892(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(un9_0_s_6),.I3(un9_0_s_7),.O(N_62));
defparam desc892.INIT=16'hF960;
  LUT6 desc893(.I0(N_454),.I1(SUM1_0_i_1_1),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.I4(un9_0_s_0),.I5(un9_0_s_1),.O(N_56));
defparam desc893.INIT=64'hFFFF3013CFEC0000;
  LUT4 desc894(.I0(ret_val[1:1]),.I1(un9_0_axb_8),.I2(un9_0_s_4),.I3(un9_0_s_5),.O(N_33_0));
defparam desc894.INIT=16'hF690;
  LUT5 output_reg_pipe_15_RNIJLNH1(.I0(un14_pos_outputf[6:6]),.I1(output_reg_pipe_15),.I2(pre_outputf[6:6]),.I3(un4_overflow_if),.I4(output_reg_pipe_13),.O(N_434_i));
defparam output_reg_pipe_15_RNIJLNH1.INIT=32'h22277277;
  LUT5 output_reg_pipe_10_RNI4LNH1(.I0(un14_pos_outputf[5:5]),.I1(output_reg_pipe_10),.I2(pre_outputf[5:5]),.I3(un4_overflow_if),.I4(output_reg_pipe_13),.O(N_431_i));
defparam output_reg_pipe_10_RNI4LNH1.INIT=32'h22277277;
  LUT5 output_reg_pipe_5_RNI0B2S(.I0(un14_pos_outputf[4:4]),.I1(output_reg_pipe_5),.I2(pre_outputf[4:4]),.I3(un4_overflow_if),.I4(output_reg_pipe_13),.O(N_428_i));
defparam output_reg_pipe_5_RNI0B2S.INIT=32'h22277277;
  LUT5 output_reg_pipe_1_RNI23E61(.I0(un14_pos_outputf[3:3]),.I1(output_reg_pipe),.I2(pre_outputf[3:3]),.I3(un4_overflow_if),.I4(output_reg_pipe_13),.O(N_425_i));
defparam output_reg_pipe_1_RNI23E61.INIT=32'h22277277;
  LUT5 desc895(.I0(shift_amount_1_i[2:2]),.I1(shift_amount_1[1:1]),.I2(un9_0_s_0),.I3(un9_0_s_1),.I4(un9_0_s_2),.O(N_79));
defparam desc895.INIT=32'hBA329810;
  LUT5 desc896(.I0(shift_amount_1_i[2:2]),.I1(shift_amount_1[1:1]),.I2(un9_0_s_2),.I3(N_56),.I4(un9_0_s_3),.O(N_80));
defparam desc896.INIT=32'hF7A2D580;
  LUT6_L desc897(.I0(shift_amount_1_i[2:2]),.I1(N_100_i),.I2(shift_amount_1[1:1]),.I3(un9_0_s_1),.I4(un9_0_s_2),.I5(un9_0_s_3),.LO(un11_output_1_Z[5:5]));
defparam desc897.INIT=64'h4644060442400200;
  LUT6_L desc898(.I0(shift_amount_1_i[2:2]),.I1(N_100_i),.I2(shift_amount_1[1:1]),.I3(un9_0_s_0),.I4(un9_0_s_1),.I5(un9_0_s_2),.LO(un11_output_1_Z[4:4]));
defparam desc898.INIT=64'h4644060442400200;
  LUT6 desc899(.I0(N_419),.I1(N_378),.I2(N_100_i),.I3(un9_0_s_1),.I4(un9_0_s_2),.I5(un9_0_s_3),.O(N_49));
defparam desc899.INIT=64'hEA62C840AA228800;
  LUT6 desc900(.I0(N_419),.I1(N_378),.I2(N_100_i),.I3(un9_0_s_2),.I4(un9_0_s_3),.I5(un9_0_s_4),.O(N_50));
defparam desc900.INIT=64'hEA62C840AA228800;
  LUT6_L desc901(.I0(N_378),.I1(N_100_i),.I2(out_shift_amount[1:1]),.I3(un9_0_s_2),.I4(un9_0_s_3),.I5(un9_0_s_4),.LO(un11_output_1_Z[6:6]));
defparam desc901.INIT=64'hC2C0828042400200;
  LUT6_L m17_0_2_cZ(.I0(N_378),.I1(out_shift_amount[1:1]),.I2(un3_shift_right),.I3(un9_0_s_4),.I4(un9_0_s_5),.I5(un9_0_s_8),.LO(m17_0_2));
defparam m17_0_2_cZ.INIT=64'h1C1814100C080400;
  LUT6 m25_0(.I0(N_378),.I1(out_shift_amount[1:1]),.I2(un3_shift_right),.I3(un9_0_s_8),.I4(un9_0_s_7),.I5(m25_0_0),.O(N_413));
defparam m25_0.INIT=64'hFFFFFFFF23012200;
  LUT6 desc902(.I0(shift_amount_1_i[2:2]),.I1(N_378),.I2(N_100_i),.I3(un9_0_s_4),.I4(un9_0_s_5),.I5(un11_output_1_Z[5:5]),.O(un11_output_1));
defparam desc902.INIT=64'hFFFFFFFFA0802000;
  LUT6 desc903(.I0(shift_amount_1_i[2:2]),.I1(N_378),.I2(N_100_i),.I3(un9_0_s_3),.I4(un9_0_s_4),.I5(un11_output_1_Z[4:4]),.O(un11_output[4:4]));
defparam desc903.INIT=64'hFFFFFFFFA0802000;
  LUT6 desc904(.I0(un20_output_0_0_a2_0_0_lut6_2_O5),.I1(N_378),.I2(un3_shift_right),.I3(un9_0_s_6),.I4(un9_0_s_7),.I5(un11_output_6_d_0[9:9]),.O(pre_output[9:9]));
defparam desc904.INIT=64'h0F0D07050A080200;
  LUT6 m34(.I0(N_100_i),.I1(out_shift_amount[1:1]),.I2(shift_amount_1[1:1]),.I3(un3_shift_right),.I4(un9_0_s_8),.I5(un9_0_s_7),.O(pre_output[11:11]));
defparam m34.INIT=64'h0081000100800000;
  LUT6 desc905(.I0(N_378),.I1(N_100_i),.I2(out_shift_amount[1:1]),.I3(un9_0_s_3),.I4(un9_0_s_4),.I5(un9_0_s_5),.O(N_51));
defparam desc905.INIT=64'h8C8488800C040800;
  LUT6 m17_0(.I0(N_378),.I1(out_shift_amount[1:1]),.I2(un3_shift_right),.I3(un9_0_s_6),.I4(un9_0_s_7),.I5(m17_0_2),.O(N_18_0));
defparam m17_0.INIT=64'hFFFFFFFF23220100;
  LUT6 desc906(.I0(N_378),.I1(N_100_i),.I2(out_shift_amount[1:1]),.I3(un9_0_s_5),.I4(un9_0_s_6),.I5(un11_output_1_Z[6:6]),.O(un11_output_2));
defparam desc906.INIT=64'hFFFFFFFF0C080400;
  LUT6 desc907(.I0(pre_output[11:11]),.I1(pre_output[10:10]),.I2(pre_output[9:9]),.I3(pre_output[8:8]),.I4(un1_apply_nrlt8_1),.I5(un1_apply_nrlt7),.O(N_420));
defparam desc907.INIT=64'h0101011101110111;
  LUT5_L output_reg_pipe_5_RNO(.I0(input_reg[10:10]),.I1(input_reg[11:11]),.I2(un4_overflow_0),.I3(pre_output[4:4]),.I4(N_420),.LO(N_427));
defparam output_reg_pipe_5_RNO.INIT=32'h000000EF;
  LUT5_L output_reg_pipe_10_RNO(.I0(input_reg[10:10]),.I1(input_reg[11:11]),.I2(un4_overflow_0),.I3(pre_output[5:5]),.I4(N_420),.LO(N_430));
defparam output_reg_pipe_10_RNO.INIT=32'h000000EF;
  LUT5_L output_reg_pipe_15_RNO(.I0(input_reg[10:10]),.I1(input_reg[11:11]),.I2(un4_overflow_0),.I3(pre_output[6:6]),.I4(N_420),.LO(N_433));
defparam output_reg_pipe_15_RNO.INIT=32'h000000EF;
  LUT4 desc908(.I0(un20_output_2[14:14]),.I1(un3_shift_right),.I2(N_56),.I3(N_49),.O(pre_output[1:1]));
defparam desc908.INIT=16'hEC20;
  LUT4 desc909(.I0(un3_shift_right),.I1(un7_output_2_0_0[6:6]),.I2(un7_output_2_1[6:6]),.I3(un11_output_2),.O(pre_output[6:6]));
defparam desc909.INIT=16'hD580;
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT4 m27_lut6_2_o6(.I0(ret_val[2:2]),.I1(un9_0_axb_8),.I2(shift_amount_1[1:1]),.I3(un9_0_s_6),.O(N_414));
defparam m27_lut6_2_o6.INIT=16'h0600;
  LUT4 m27_lut6_2_o5(.I0(ret_val[2:2]),.I1(un9_0_axb_8),.I2(shift_amount_1[1:1]),.I3(un9_0_s_7),.O(N_33));
defparam m27_lut6_2_o5.INIT=16'h0600;
  LUT4 output_reg_pipe_12_RNIPJ901_o6(.I0(input_reg[10:10]),.I1(input_reg[11:11]),.I2(done_inv_sqrt),.I3(un4_overflow_0),.O(output_reg_pipe_12_RNIPJ901_O6));
defparam output_reg_pipe_12_RNIPJ901_o6.INIT=16'h1000;
  LUT5 output_reg_pipe_12_RNIPJ901_o5(.I0(un4_overflow_if),.I1(input_reg[10:10]),.I2(input_reg[11:11]),.I3(done_inv_sqrt),.I4(un4_overflow_0),.O(un4_overflow_i_0));
defparam output_reg_pipe_12_RNIPJ901_o5.INIT=32'hFCAAFFAA;
endmodule
module shifterZ1_inj (ret_val,un20_output_2,ret_val_m2,shift_amount_1,un26_output_0_iv_3,ret_val_d_a1,ret_val_d_a0,un26_output_6,un26_output_2,un26_output_4,un26_output_3,un26_output_0,un1_poly_odd_i,input_reg,un26_output_0_iv_2_0_1,input_shifted_4,input_shifted_0,input_shifted_3,un1_input_shifted,un1_poly_odd,un9_0_axb_8,un20_output_0_0_a2_0_0_lut6_2_O5,N_100_i,N_65,un3_shift_right,N_2502_i,un4_overflow_2,N_454,N_72,ret_val_ss0,N_458,N_45,N_70,N_73,N_71,N_441,un9_0_axb_4);
input [3:1] ret_val ;
output [14:14] un20_output_2 ;
input [3:3] ret_val_m2 ;
input [1:1] shift_amount_1 ;
output [6:6] un26_output_0_iv_3 ;
input [1:1] ret_val_d_a1 ;
input [1:1] ret_val_d_a0 ;
output un26_output_6 ;
output un26_output_2 ;
output un26_output_4 ;
output un26_output_3 ;
output un26_output_0 ;
output [6:6] un1_poly_odd_i ;
input [11:0] input_reg ;
output un26_output_0_iv_2_0_1 ;
output input_shifted_4 ;
output input_shifted_0 ;
output input_shifted_3 ;
input [4:4] un1_input_shifted ;
input [8:8] un1_poly_odd ;
input un9_0_axb_8 ;
output un20_output_0_0_a2_0_0_lut6_2_O5 ;
output N_100_i ;
output N_65 ;
input un3_shift_right ;
output N_2502_i ;
input un4_overflow_2 ;
input N_454 ;
output N_72 ;
input ret_val_ss0 ;
input N_458 ;
output N_45 ;
output N_70 ;
output N_73 ;
output N_71 ;
input N_441 ;
output un9_0_axb_4 ;
wire un26_output_6 ;
wire un26_output_2 ;
wire un26_output_4 ;
wire un26_output_3 ;
wire un26_output_0 ;
wire un26_output_0_iv_2_0_1 ;
wire input_shifted_4 ;
wire input_shifted_0 ;
wire input_shifted_3 ;
wire un9_0_axb_8 ;
wire un20_output_0_0_a2_0_0_lut6_2_O5 ;
wire N_100_i ;
wire N_65 ;
wire un3_shift_right ;
wire N_2502_i ;
wire un4_overflow_2 ;
wire N_454 ;
wire N_72 ;
wire ret_val_ss0 ;
wire N_458 ;
wire N_45 ;
wire N_70 ;
wire N_73 ;
wire N_71 ;
wire N_441 ;
wire un9_0_axb_4 ;
wire [4:4] input_m_s ;
wire [5:5] un26_output_0_iv_2_0 ;
wire [3:3] input_m_0 ;
wire [2:2] output_a1_0 ;
wire [3:3] un26_output_0_iv_0 ;
wire [4:4] un26_output_0_iv_2_a0 ;
wire [1:0] input_m_4 ;
wire input_m_2 ;
wire [2:2] input_m_3 ;
wire [7:7] un26_output_0_iv_0_a2_xx ;
wire [7:7] un26_output_0_iv_0_a2_yy ;
wire input_m_4_a0_0 ;
wire [2:2] output_0_2 ;
wire GND ;
wire VCC ;
wire un20_output_0_0_a2_0_0 ;
wire N_47 ;
wire un20_output_0_2_a0_0 ;
wire un20_output_3_0_0_a2_s ;
wire un26_m3_i_0 ;
wire N_46 ;
wire N_443 ;
wire N_445 ;
// instances
  LUT4 desc845(.I0(N_65),.I1(un26_output_6),.I2(un3_shift_right),.I3(un9_0_axb_8),.O(N_2502_i));
defparam desc845.INIT=16'h00AC;
  LUT4 un20_output_0(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(un20_output_0_2_a0_0),.I3(ret_val[3:3]),.O(un20_output_2[14:14]));
defparam un20_output_0.INIT=16'h00DF;
  LUT5 un20_output_1_0_0_a2_0(.I0(input_reg[3:3]),.I1(un4_overflow_2),.I2(ret_val_m2[3:3]),.I3(N_454),.I4(un9_0_axb_8),.O(un20_output_3_0_0_a2_s));
defparam un20_output_1_0_0_a2_0.INIT=32'h000037FF;
  LUT5 desc846(.I0(input_reg[3:3]),.I1(input_reg[6:6]),.I2(un9_0_axb_8),.I3(input_m_s[4:4]),.I4(shift_amount_1[1:1]),.O(un26_output_0_iv_3[6:6]));
defparam desc846.INIT=32'hFF0ACCC0;
  LUT3 desc847(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(un9_0_axb_8),.O(un26_output_0_iv_2_0[5:5]));
defparam desc847.INIT=8'hCA;
  LUT4 desc848(.I0(input_reg[3:3]),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(input_m_0[3:3]));
defparam desc848.INIT=16'h2A00;
  LUT5 desc849(.I0(input_reg[8:8]),.I1(input_reg[7:7]),.I2(un9_0_axb_8),.I3(N_47),.I4(shift_amount_1[1:1]),.O(N_72));
defparam desc849.INIT=32'hCACAFF00;
  LUT6 desc850(.I0(input_reg[2:2]),.I1(ret_val_ss0),.I2(ret_val_d_a1[1:1]),.I3(N_458),.I4(ret_val_d_a0[1:1]),.I5(N_454),.O(output_a1_0[2:2]));
defparam desc850.INIT=64'h1155115055555050;
  LUT6 desc851(.I0(input_reg[2:2]),.I1(un9_0_axb_8),.I2(un20_output_2[14:14]),.I3(input_m_0[3:3]),.I4(shift_amount_1[1:1]),.I5(un26_output_0_iv_0[3:3]),.O(un26_output_2));
defparam desc851.INIT=64'hFFFFFFFF0000FF20;
  LUT6 desc852(.I0(input_reg[2:2]),.I1(un9_0_axb_8),.I2(un26_output_0_iv_2_0[5:5]),.I3(un26_m3_i_0),.I4(input_m_0[3:3]),.I5(shift_amount_1[1:1]),.O(un26_output_4));
defparam desc852.INIT=64'hFFFFFF22FFF0FFF0;
  LUT6 desc853(.I0(input_reg[3:3]),.I1(un9_0_axb_8),.I2(un20_output_2[14:14]),.I3(input_m_s[4:4]),.I4(un26_output_0_iv_2_a0[4:4]),.I5(shift_amount_1[1:1]),.O(un26_output_3));
defparam desc853.INIT=64'h0000FFFFFF20FF2F;
  LUT6 desc854(.I0(input_reg[5:5]),.I1(input_reg[6:6]),.I2(un9_0_axb_8),.I3(un20_output_2[14:14]),.I4(N_45),.I5(shift_amount_1[1:1]),.O(N_70));
defparam desc854.INIT=64'hAC00AC00FF000000;
  LUT6 desc855(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[7:7]),.I3(input_reg[6:6]),.I4(un9_0_axb_8),.I5(shift_amount_1[1:1]),.O(N_73));
defparam desc855.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc856(.I0(input_reg[7:7]),.I1(input_reg[6:6]),.I2(un9_0_axb_8),.I3(un20_output_2[14:14]),.I4(N_46),.I5(shift_amount_1[1:1]),.O(N_71));
defparam desc856.INIT=64'hCACACACAFF000000;
  LUT4 desc857(.I0(input_reg[1:1]),.I1(ret_val[3:3]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(input_m_4[1:1]));
defparam desc857.INIT=16'h0008;
  LUT4 desc858(.I0(input_reg[4:4]),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(input_m_s[4:4]));
defparam desc858.INIT=16'h2A00;
  LUT4_L desc859(.I0(input_reg[0:0]),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.LO(input_m_2));
defparam desc859.INIT=16'h8000;
  LUT4 desc860(.I0(input_reg[2:2]),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(input_m_3[2:2]));
defparam desc860.INIT=16'h8000;
  LUT5_L desc861(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(un9_0_axb_8),.I3(un20_output_2[14:14]),.I4(shift_amount_1[1:1]),.LO(un26_output_0_iv_0[3:3]));
defparam desc861.INIT=32'hCA000000;
  LUT5 desc862(.I0(input_reg[1:1]),.I1(input_reg[2:2]),.I2(un9_0_axb_8),.I3(un20_output_2[14:14]),.I4(input_m_2),.O(un26_output_0_iv_2_a0[4:4]));
defparam desc862.INIT=32'h000035FF;
  LUT5 desc863(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(un9_0_axb_8),.I3(un20_output_0_0_a2_0_0),.I4(shift_amount_1[1:1]),.O(un26_output_0));
defparam desc863.INIT=32'h0000CA00;
  LUT5 desc864(.I0(N_443),.I1(N_445),.I2(un26_output_0_iv_0_a2_xx[7:7]),.I3(un26_output_0_iv_0_a2_yy[7:7]),.I4(shift_amount_1[1:1]),.O(un26_output_6));
defparam desc864.INIT=32'hFFAAFCFC;
  LUT5 desc865(.I0(un9_0_axb_8),.I1(un3_shift_right),.I2(N_65),.I3(un26_output_6),.I4(input_shifted_4),.O(un1_poly_odd_i[6:6]));
defparam desc865.INIT=32'hF7D5A280;
  LUT3 desc866(.I0(input_reg[3:3]),.I1(input_reg[4:4]),.I2(un9_0_axb_8),.O(N_45));
defparam desc866.INIT=8'hAC;
  LUT3 desc867(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(un9_0_axb_8),.O(N_46));
defparam desc867.INIT=8'hAC;
  LUT3 desc868(.I0(input_reg[7:7]),.I1(input_reg[6:6]),.I2(un9_0_axb_8),.O(N_445));
defparam desc868.INIT=8'hAC;
  LUT3 desc869(.I0(input_reg[4:4]),.I1(input_reg[5:5]),.I2(un9_0_axb_8),.O(N_443));
defparam desc869.INIT=8'hCA;
  LUT6 un20_output_0_2_a0_0_0(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[7:7]),.I3(input_reg[10:10]),.I4(input_reg[11:11]),.I5(input_reg[6:6]),.O(un20_output_0_2_a0_0));
defparam un20_output_0_2_a0_0_0.INIT=64'h0000000000000001;
  LUT6 desc870(.I0(input_reg[0:0]),.I1(input_reg[7:7]),.I2(input_reg[11:11]),.I3(input_reg[6:6]),.I4(un4_overflow_2),.I5(N_441),.O(input_m_4_a0_0));
defparam desc870.INIT=64'hAAAAAAAAA0A2A0A0;
  LUT4 desc871(.I0(input_m_4_a0_0),.I1(ret_val[3:3]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(input_m_4[0:0]));
defparam desc871.INIT=16'h0800;
  LUT6 desc872(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(ret_val[2:2]),.I3(output_a1_0[2:2]),.I4(ret_val[3:3]),.I5(un9_0_axb_8),.O(output_0_2[2:2]));
defparam desc872.INIT=64'h000000AF0000CFCF;
  LUT6 un26_m3_i_0_cZ(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(ret_val[2:2]),.I3(ret_val[3:3]),.I4(ret_val[1:1]),.I5(un9_0_axb_8),.O(un26_m3_i_0));
defparam un26_m3_i_0_cZ.INIT=64'h00C0000000000A00;
  LUT6 desc873(.I0(input_reg[0:0]),.I1(input_reg[1:1]),.I2(ret_val[2:2]),.I3(ret_val[3:3]),.I4(ret_val[1:1]),.I5(un9_0_axb_8),.O(un26_output_0_iv_0_a2_yy[7:7]));
defparam desc873.INIT=64'h00C00C000A000A00;
  LUT6 desc874(.I0(input_reg[2:2]),.I1(input_reg[3:3]),.I2(ret_val[2:2]),.I3(ret_val[3:3]),.I4(ret_val[1:1]),.I5(un9_0_axb_8),.O(un26_output_0_iv_0_a2_xx[7:7]));
defparam desc874.INIT=64'h00C00C000A000A00;
  LUT6 desc875(.I0(input_reg[9:9]),.I1(input_reg[8:8]),.I2(input_reg[7:7]),.I3(input_reg[10:10]),.I4(un9_0_axb_8),.I5(shift_amount_1[1:1]),.O(N_65));
defparam desc875.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc876(.I0(input_reg[3:3]),.I1(ret_val[2:2]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.I4(output_0_2[2:2]),.I5(N_46),.O(input_shifted_0));
defparam desc876.INIT=64'h3F2F00003C2C0000;
  LUT6 desc877(.I0(input_reg[5:5]),.I1(un20_output_3_0_0_a2_s),.I2(input_m_3[2:2]),.I3(input_m_4[0:0]),.I4(input_m_4[1:1]),.I5(shift_amount_1[1:1]),.O(un26_output_0_iv_2_0_1));
defparam desc877.INIT=64'hFFFFFFF0FFFFFFF8;
  LUT3 desc878(.I0(un3_shift_right),.I1(N_72),.I2(un26_output_4),.O(input_shifted_3));
defparam desc878.INIT=8'hD8;
  LUT4 desc879(.I0(un3_shift_right),.I1(N_73),.I2(un26_output_0_iv_3[6:6]),.I3(un26_output_0_iv_2_0_1),.O(input_shifted_4));
defparam desc879.INIT=16'hDDD8;
  LUT5 desc880(.I0(un9_0_axb_8),.I1(input_shifted_3),.I2(un1_input_shifted[4:4]),.I3(un1_poly_odd[8:8]),.I4(input_shifted_4),.O(un9_0_axb_4));
defparam desc880.INIT=32'hEBB1411B;
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT3 desc881(.I0(input_reg[5:5]),.I1(input_reg[6:6]),.I2(un9_0_axb_8),.O(N_47));
defparam desc881.INIT=8'hAC;
  LUT3 desc882(.I0(ret_val[3:3]),.I1(ret_val[1:1]),.I2(un9_0_axb_8),.O(N_100_i));
defparam desc882.INIT=8'h7F;
  LUT3 un20_output_0_0_a2_0_0_lut6_2_o6(.I0(ret_val[2:2]),.I1(ret_val[3:3]),.I2(ret_val[1:1]),.O(un20_output_0_0_a2_0_0));
defparam un20_output_0_0_a2_0_0_lut6_2_o6.INIT=8'h13;
  LUT4 un20_output_0_0_a2_0_0_lut6_2_o5(.I0(ret_val[2:2]),.I1(ret_val[3:3]),.I2(ret_val[1:1]),.I3(un9_0_axb_8),.O(un20_output_0_0_a2_0_0_lut6_2_O5));
defparam un20_output_0_0_a2_0_0_lut6_2_o5.INIT=16'h2444;
endmodule
module vec_mult_inj (in_b_vec_mult_sel,out_inner_prod_i,out_i_vec_mult_2,out_r_vec_mult_2,out_inner_prod_r,vec_out_r_AQ_2,out_inv_sqrt_0,out_inv_sqrt_1,out_inv_sqrt_2,out_inv_sqrt_7,out_inv_sqrt_8,out_inv_sqrt_9,out_inv_sqrt_10,out_inv_sqrt_11,vec_out_i_AQ_2,out_i_vec_mult_1,out_r_vec_mult_1,vec_out_r_AQ_1,vec_out_i_AQ_1,out_i_vec_mult_0,out_r_vec_mult_0,vec_out_r_AQ_0,vec_out_i_AQ_0,out_i_vec_mult_3,out_r_vec_mult_3,vec_out_r_AQ_3,vec_out_i_AQ_3,clk,N_425_i,N_428_i,N_431_i,N_434_i);
input in_b_vec_mult_sel ;
input [11:0] out_inner_prod_i ;
output [11:0] out_i_vec_mult_2 ;
output [11:0] out_r_vec_mult_2 ;
input [11:0] out_inner_prod_r ;
input [11:0] vec_out_r_AQ_2 ;
input out_inv_sqrt_0 ;
input out_inv_sqrt_1 ;
input out_inv_sqrt_2 ;
input out_inv_sqrt_7 ;
input out_inv_sqrt_8 ;
input out_inv_sqrt_9 ;
input out_inv_sqrt_10 ;
input out_inv_sqrt_11 ;
input [11:0] vec_out_i_AQ_2 ;
output [11:0] out_i_vec_mult_1 ;
output [11:0] out_r_vec_mult_1 ;
input [11:0] vec_out_r_AQ_1 ;
input [11:0] vec_out_i_AQ_1 ;
output [11:0] out_i_vec_mult_0 ;
output [11:0] out_r_vec_mult_0 ;
input [11:0] vec_out_r_AQ_0 ;
input [11:0] vec_out_i_AQ_0 ;
output [11:0] out_i_vec_mult_3 ;
output [11:0] out_r_vec_mult_3 ;
input [11:0] vec_out_r_AQ_3 ;
input [11:0] vec_out_i_AQ_3 ;
input clk ;
input N_425_i ;
input N_428_i ;
input N_431_i ;
input N_434_i ;
wire out_inv_sqrt_0 ;
wire out_inv_sqrt_1 ;
wire out_inv_sqrt_2 ;
wire out_inv_sqrt_7 ;
wire out_inv_sqrt_8 ;
wire out_inv_sqrt_9 ;
wire out_inv_sqrt_10 ;
wire out_inv_sqrt_11 ;
wire clk ;
wire N_425_i ;
wire N_428_i ;
wire N_431_i ;
wire N_434_i ;
wire [11:0] in_b_i_reg ;
wire GND ;
wire VCC ;
// instances
  FDR desc695(.Q(in_b_i_reg[11:11]),.D(out_inner_prod_i[11:11]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc696(.Q(in_b_i_reg[10:10]),.D(out_inner_prod_i[10:10]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc697(.Q(in_b_i_reg[9:9]),.D(out_inner_prod_i[9:9]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc698(.Q(in_b_i_reg[8:8]),.D(out_inner_prod_i[8:8]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc699(.Q(in_b_i_reg[7:7]),.D(out_inner_prod_i[7:7]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc700(.Q(in_b_i_reg[6:6]),.D(out_inner_prod_i[6:6]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc701(.Q(in_b_i_reg[5:5]),.D(out_inner_prod_i[5:5]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc702(.Q(in_b_i_reg[4:4]),.D(out_inner_prod_i[4:4]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc703(.Q(in_b_i_reg[3:3]),.D(out_inner_prod_i[3:3]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc704(.Q(in_b_i_reg[2:2]),.D(out_inner_prod_i[2:2]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc705(.Q(in_b_i_reg[1:1]),.D(out_inner_prod_i[1:1]),.C(clk),.R(in_b_vec_mult_sel));
  FDR desc706(.Q(in_b_i_reg[0:0]),.D(out_inner_prod_i[0:0]),.C(clk),.R(in_b_vec_mult_sel));
  desc481_inj desc707(.out_i_vec_mult_2(out_i_vec_mult_2[11:0]),.out_r_vec_mult_2(out_r_vec_mult_2[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_2(vec_out_r_AQ_2[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.vec_out_i_AQ_2(vec_out_i_AQ_2[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  desc536_inj desc708(.out_i_vec_mult_1(out_i_vec_mult_1[11:0]),.out_r_vec_mult_1(out_r_vec_mult_1[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_1(vec_out_r_AQ_1[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.vec_out_i_AQ_1(vec_out_i_AQ_1[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  desc591_inj desc709(.out_i_vec_mult_0(out_i_vec_mult_0[11:0]),.out_r_vec_mult_0(out_r_vec_mult_0[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_0(vec_out_r_AQ_0[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.vec_out_i_AQ_0(vec_out_i_AQ_0[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  desc646_inj desc710(.out_i_vec_mult_3(out_i_vec_mult_3[11:0]),.out_r_vec_mult_3(out_r_vec_mult_3[11:0]),.out_inner_prod_r(out_inner_prod_r[11:0]),.vec_out_r_AQ_3(vec_out_r_AQ_3[11:0]),.out_inv_sqrt_0(out_inv_sqrt_0),.out_inv_sqrt_1(out_inv_sqrt_1),.out_inv_sqrt_2(out_inv_sqrt_2),.out_inv_sqrt_7(out_inv_sqrt_7),.out_inv_sqrt_8(out_inv_sqrt_8),.out_inv_sqrt_9(out_inv_sqrt_9),.out_inv_sqrt_10(out_inv_sqrt_10),.out_inv_sqrt_11(out_inv_sqrt_11),.in_b_vec_mult_sel(in_b_vec_mult_sel),.vec_out_i_AQ_3(vec_out_i_AQ_3[11:0]),.out_inner_prod_i(out_inner_prod_i[11:0]),.in_b_i_reg(in_b_i_reg[11:0]),.clk(clk),.N_425_i(N_425_i),.N_428_i(N_428_i),.N_431_i(N_431_i),.N_434_i(N_434_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
module vec_sub_inj (in_a_r_reg_3_11,in_a_r_reg_2_11,in_a_r_reg_1_11,in_a_r_reg_0_0,in_a_r_reg_0_11,out_Q_r,in_a_i_reg_3_11,in_a_i_reg_2_11,in_a_i_reg_1_11,in_a_i_reg_0_11,out_Q_i,out_r_vec_mult_0,out_r_vec_mult_1,out_r_vec_mult_2,pre_out,out_r_vec_mult_3,pre_out_i_m_1,pre_out_0,output_iv,output_iv_0_0,output_iv_0_1,output_iv_0_2,output_iv_0_3,output_iv_0_4,output_iv_0_6,output_iv_0_7,output_iv_0_8,output_iv_0_9,out_i_vec_sub_0,out_i_vec_mult_0,pre_out_i_m_2,out_i_vec_mult_1,pre_out_1,pre_out_4,pre_out_i_m_3,out_i_vec_mult_2,pre_out_2,pre_out_5,out_i_vec_mult_3,pre_out_i_m,pre_out_i_m_0_0,pre_out_i_m_0_1,pre_out_i_m_0_6,pre_out_i_m_0_4,pre_out_i_m_4,pre_out_6,pre_out_3_9,pre_out_3_0,pre_out_3_1,pre_out_3_3,pre_out_3_5,pre_out_3_7,pre_out_3_8,pre_out_3_6,clk,w_in_a_vec_sub,N_500,un5_output,un5_output_0,un5_output_1,un5_output_2,un5_output_3,un5_output_4,p_desc739_p_O_FDE,p_desc740_p_O_FDE,p_desc741_p_O_FDE,p_desc742_p_O_FDE,p_desc743_p_O_FDE,p_desc744_p_O_FDE,p_desc745_p_O_FDE,p_desc746_p_O_FDE,p_desc747_p_O_FDE,p_desc748_p_O_FDE,p_desc749_p_O_FDE,p_desc750_p_O_FDE,p_desc751_p_O_FDE,p_desc752_p_O_FDE,p_desc753_p_O_FDE,p_desc754_p_O_FDE,p_desc755_p_O_FDE,p_desc756_p_O_FDE,p_desc757_p_O_FDE,p_desc758_p_O_FDE,p_desc759_p_O_FDE,p_desc760_p_O_FDE,p_desc761_p_O_FDE,p_desc762_p_O_FDE,p_desc763_p_O_FDE,p_desc764_p_O_FDE,p_desc765_p_O_FDE,p_desc766_p_O_FDE,p_desc767_p_O_FDE,p_desc768_p_O_FDE,p_desc769_p_O_FDE,p_desc770_p_O_FDE,p_desc771_p_O_FDE,p_desc772_p_O_FDE,p_desc773_p_O_FDE,p_desc774_p_O_FDE,p_desc775_p_O_FDE,p_desc776_p_O_FDE,p_desc777_p_O_FDE,p_desc778_p_O_FDE,p_desc779_p_O_FDE,p_desc780_p_O_FDE,p_desc781_p_O_FDE,p_desc782_p_O_FDE,p_desc783_p_O_FDE,p_desc784_p_O_FDE,p_desc785_p_O_FDE,p_desc786_p_O_FDE,p_desc787_p_O_FDE,p_desc788_p_O_FDE,p_desc789_p_O_FDE,p_desc790_p_O_FDE,p_desc791_p_O_FDE,p_desc792_p_O_FDE,p_desc793_p_O_FDE,p_desc794_p_O_FDE,p_desc795_p_O_FDE,p_desc796_p_O_FDE,p_desc797_p_O_FDE,p_desc798_p_O_FDE,p_desc799_p_O_FDE,p_desc800_p_O_FDE,p_desc801_p_O_FDE,p_desc802_p_O_FDE,p_desc803_p_O_FDE,p_desc804_p_O_FDE,p_desc805_p_O_FDE,p_desc806_p_O_FDE,p_desc807_p_O_FDE,p_desc808_p_O_FDE,p_desc809_p_O_FDE,p_desc810_p_O_FDE,p_desc811_p_O_FDE,p_desc812_p_O_FDE,p_desc813_p_O_FDE,p_desc814_p_O_FDE,p_desc815_p_O_FDE,p_desc816_p_O_FDE,p_desc817_p_O_FDE,p_desc818_p_O_FDE,p_desc819_p_O_FDE,p_desc820_p_O_FDE,p_desc821_p_O_FDE,p_desc822_p_O_FDE,p_desc823_p_O_FDE,p_desc824_p_O_FDE,p_desc825_p_O_FDE,p_desc826_p_O_FDE,p_desc827_p_O_FDE,p_desc828_p_O_FDE,p_desc829_p_O_FDE,p_desc830_p_O_FDE,p_desc831_p_O_FDE,p_desc832_p_O_FDE,p_desc833_p_O_FDE,p_desc834_p_O_FDE);
output in_a_r_reg_3_11 ;
output in_a_r_reg_2_11 ;
output in_a_r_reg_1_11 ;
output in_a_r_reg_0_0 ;
output in_a_r_reg_0_11 ;
input [47:0] out_Q_r ;
output in_a_i_reg_3_11 ;
output in_a_i_reg_2_11 ;
output in_a_i_reg_1_11 ;
output in_a_i_reg_0_11 ;
input [47:0] out_Q_i ;
input [11:0] out_r_vec_mult_0 ;
input [11:0] out_r_vec_mult_1 ;
input [11:0] out_r_vec_mult_2 ;
output [11:1] pre_out ;
input [11:0] out_r_vec_mult_3 ;
output pre_out_i_m_1 ;
output [11:1] pre_out_0 ;
output [10:0] output_iv ;
output output_iv_0_0 ;
output output_iv_0_1 ;
output output_iv_0_2 ;
output output_iv_0_3 ;
output output_iv_0_4 ;
output output_iv_0_6 ;
output output_iv_0_7 ;
output output_iv_0_8 ;
output output_iv_0_9 ;
output [11:11] out_i_vec_sub_0 ;
input [11:0] out_i_vec_mult_0 ;
output pre_out_i_m_2 ;
input [11:0] out_i_vec_mult_1 ;
output [11:1] pre_out_1 ;
output [11:11] pre_out_4 ;
output pre_out_i_m_3 ;
input [11:0] out_i_vec_mult_2 ;
output [11:1] pre_out_2 ;
output [11:11] pre_out_5 ;
input [11:0] out_i_vec_mult_3 ;
output [10:0] pre_out_i_m ;
output pre_out_i_m_0_0 ;
output pre_out_i_m_0_1 ;
output pre_out_i_m_0_6 ;
output pre_out_i_m_0_4 ;
output pre_out_i_m_4 ;
output [11:11] pre_out_6 ;
output pre_out_3_9 ;
output pre_out_3_0 ;
output pre_out_3_1 ;
output pre_out_3_3 ;
output pre_out_3_5 ;
output pre_out_3_7 ;
output pre_out_3_8 ;
output pre_out_3_6 ;
input clk ;
input w_in_a_vec_sub ;
output N_500 ;
output un5_output ;
output un5_output_0 ;
output un5_output_1 ;
output un5_output_2 ;
output un5_output_3 ;
output un5_output_4 ;
wire in_a_r_reg_3_11 ;
wire in_a_r_reg_2_11 ;
wire in_a_r_reg_1_11 ;
wire in_a_r_reg_0_0 ;
wire in_a_r_reg_0_11 ;
wire in_a_i_reg_3_11 ;
wire in_a_i_reg_2_11 ;
wire in_a_i_reg_1_11 ;
wire in_a_i_reg_0_11 ;
wire output_iv_0_0 ;
wire output_iv_0_1 ;
wire output_iv_0_2 ;
wire output_iv_0_3 ;
wire output_iv_0_4 ;
wire output_iv_0_6 ;
wire output_iv_0_7 ;
wire output_iv_0_8 ;
wire output_iv_0_9 ;
wire pre_out_i_m_0_0 ;
wire pre_out_i_m_0_1 ;
wire pre_out_i_m_0_6 ;
wire pre_out_i_m_0_4 ;
wire pre_out_3_9 ;
wire pre_out_3_0 ;
wire pre_out_3_1 ;
wire pre_out_3_3 ;
wire pre_out_3_5 ;
wire pre_out_3_7 ;
wire pre_out_3_8 ;
wire pre_out_3_6 ;
wire clk ;
wire w_in_a_vec_sub ;
wire N_500 ;
wire un5_output ;
wire un5_output_0 ;
wire un5_output_1 ;
wire un5_output_2 ;
wire un5_output_3 ;
wire un5_output_4 ;
wire [10:0] in_a_r_reg_3 ;
wire [10:0] in_a_r_reg_2 ;
wire [10:0] in_a_r_reg_1 ;
wire [10:1] in_a_r_reg_0 ;
wire [10:0] in_a_i_reg_3 ;
wire [10:0] in_a_i_reg_2 ;
wire [10:0] in_a_i_reg_1 ;
wire [10:0] in_a_i_reg_0 ;
wire GND ;
wire VCC ;
input p_desc739_p_O_FDE ;
input p_desc740_p_O_FDE ;
input p_desc741_p_O_FDE ;
input p_desc742_p_O_FDE ;
input p_desc743_p_O_FDE ;
input p_desc744_p_O_FDE ;
input p_desc745_p_O_FDE ;
input p_desc746_p_O_FDE ;
input p_desc747_p_O_FDE ;
input p_desc748_p_O_FDE ;
input p_desc749_p_O_FDE ;
input p_desc750_p_O_FDE ;
input p_desc751_p_O_FDE ;
input p_desc752_p_O_FDE ;
input p_desc753_p_O_FDE ;
input p_desc754_p_O_FDE ;
input p_desc755_p_O_FDE ;
input p_desc756_p_O_FDE ;
input p_desc757_p_O_FDE ;
input p_desc758_p_O_FDE ;
input p_desc759_p_O_FDE ;
input p_desc760_p_O_FDE ;
input p_desc761_p_O_FDE ;
input p_desc762_p_O_FDE ;
input p_desc763_p_O_FDE ;
input p_desc764_p_O_FDE ;
input p_desc765_p_O_FDE ;
input p_desc766_p_O_FDE ;
input p_desc767_p_O_FDE ;
input p_desc768_p_O_FDE ;
input p_desc769_p_O_FDE ;
input p_desc770_p_O_FDE ;
input p_desc771_p_O_FDE ;
input p_desc772_p_O_FDE ;
input p_desc773_p_O_FDE ;
input p_desc774_p_O_FDE ;
input p_desc775_p_O_FDE ;
input p_desc776_p_O_FDE ;
input p_desc777_p_O_FDE ;
input p_desc778_p_O_FDE ;
input p_desc779_p_O_FDE ;
input p_desc780_p_O_FDE ;
input p_desc781_p_O_FDE ;
input p_desc782_p_O_FDE ;
input p_desc783_p_O_FDE ;
input p_desc784_p_O_FDE ;
input p_desc785_p_O_FDE ;
input p_desc786_p_O_FDE ;
input p_desc787_p_O_FDE ;
input p_desc788_p_O_FDE ;
input p_desc789_p_O_FDE ;
input p_desc790_p_O_FDE ;
input p_desc791_p_O_FDE ;
input p_desc792_p_O_FDE ;
input p_desc793_p_O_FDE ;
input p_desc794_p_O_FDE ;
input p_desc795_p_O_FDE ;
input p_desc796_p_O_FDE ;
input p_desc797_p_O_FDE ;
input p_desc798_p_O_FDE ;
input p_desc799_p_O_FDE ;
input p_desc800_p_O_FDE ;
input p_desc801_p_O_FDE ;
input p_desc802_p_O_FDE ;
input p_desc803_p_O_FDE ;
input p_desc804_p_O_FDE ;
input p_desc805_p_O_FDE ;
input p_desc806_p_O_FDE ;
input p_desc807_p_O_FDE ;
input p_desc808_p_O_FDE ;
input p_desc809_p_O_FDE ;
input p_desc810_p_O_FDE ;
input p_desc811_p_O_FDE ;
input p_desc812_p_O_FDE ;
input p_desc813_p_O_FDE ;
input p_desc814_p_O_FDE ;
input p_desc815_p_O_FDE ;
input p_desc816_p_O_FDE ;
input p_desc817_p_O_FDE ;
input p_desc818_p_O_FDE ;
input p_desc819_p_O_FDE ;
input p_desc820_p_O_FDE ;
input p_desc821_p_O_FDE ;
input p_desc822_p_O_FDE ;
input p_desc823_p_O_FDE ;
input p_desc824_p_O_FDE ;
input p_desc825_p_O_FDE ;
input p_desc826_p_O_FDE ;
input p_desc827_p_O_FDE ;
input p_desc828_p_O_FDE ;
input p_desc829_p_O_FDE ;
input p_desc830_p_O_FDE ;
input p_desc831_p_O_FDE ;
input p_desc832_p_O_FDE ;
input p_desc833_p_O_FDE ;
input p_desc834_p_O_FDE ;
// instances
  p_O_FDE desc739(.Q(in_a_r_reg_3[0:0]),.D(out_Q_r[0:0]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc739_p_O_FDE));
  p_O_FDE desc740(.Q(in_a_r_reg_3[1:1]),.D(out_Q_r[1:1]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc740_p_O_FDE));
  p_O_FDE desc741(.Q(in_a_r_reg_3[2:2]),.D(out_Q_r[2:2]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc741_p_O_FDE));
  p_O_FDE desc742(.Q(in_a_r_reg_3[3:3]),.D(out_Q_r[3:3]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc742_p_O_FDE));
  p_O_FDE desc743(.Q(in_a_r_reg_3[4:4]),.D(out_Q_r[4:4]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc743_p_O_FDE));
  p_O_FDE desc744(.Q(in_a_r_reg_3[5:5]),.D(out_Q_r[5:5]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc744_p_O_FDE));
  p_O_FDE desc745(.Q(in_a_r_reg_3[6:6]),.D(out_Q_r[6:6]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc745_p_O_FDE));
  p_O_FDE desc746(.Q(in_a_r_reg_3[7:7]),.D(out_Q_r[7:7]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc746_p_O_FDE));
  p_O_FDE desc747(.Q(in_a_r_reg_3[8:8]),.D(out_Q_r[8:8]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc747_p_O_FDE));
  p_O_FDE desc748(.Q(in_a_r_reg_3[9:9]),.D(out_Q_r[9:9]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc748_p_O_FDE));
  p_O_FDE desc749(.Q(in_a_r_reg_3[10:10]),.D(out_Q_r[10:10]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc749_p_O_FDE));
  p_O_FDE desc750(.Q(in_a_r_reg_3_11),.D(out_Q_r[11:11]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc750_p_O_FDE));
  p_O_FDE desc751(.Q(in_a_r_reg_2[0:0]),.D(out_Q_r[12:12]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc751_p_O_FDE));
  p_O_FDE desc752(.Q(in_a_r_reg_2[1:1]),.D(out_Q_r[13:13]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc752_p_O_FDE));
  p_O_FDE desc753(.Q(in_a_r_reg_2[2:2]),.D(out_Q_r[14:14]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc753_p_O_FDE));
  p_O_FDE desc754(.Q(in_a_r_reg_2[3:3]),.D(out_Q_r[15:15]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc754_p_O_FDE));
  p_O_FDE desc755(.Q(in_a_r_reg_2[4:4]),.D(out_Q_r[16:16]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc755_p_O_FDE));
  p_O_FDE desc756(.Q(in_a_r_reg_2[5:5]),.D(out_Q_r[17:17]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc756_p_O_FDE));
  p_O_FDE desc757(.Q(in_a_r_reg_2[6:6]),.D(out_Q_r[18:18]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc757_p_O_FDE));
  p_O_FDE desc758(.Q(in_a_r_reg_2[7:7]),.D(out_Q_r[19:19]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc758_p_O_FDE));
  p_O_FDE desc759(.Q(in_a_r_reg_2[8:8]),.D(out_Q_r[20:20]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc759_p_O_FDE));
  p_O_FDE desc760(.Q(in_a_r_reg_2[9:9]),.D(out_Q_r[21:21]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc760_p_O_FDE));
  p_O_FDE desc761(.Q(in_a_r_reg_2[10:10]),.D(out_Q_r[22:22]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc761_p_O_FDE));
  p_O_FDE desc762(.Q(in_a_r_reg_2_11),.D(out_Q_r[23:23]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc762_p_O_FDE));
  p_O_FDE desc763(.Q(in_a_r_reg_1[0:0]),.D(out_Q_r[24:24]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc763_p_O_FDE));
  p_O_FDE desc764(.Q(in_a_r_reg_1[1:1]),.D(out_Q_r[25:25]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc764_p_O_FDE));
  p_O_FDE desc765(.Q(in_a_r_reg_1[2:2]),.D(out_Q_r[26:26]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc765_p_O_FDE));
  p_O_FDE desc766(.Q(in_a_r_reg_1[3:3]),.D(out_Q_r[27:27]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc766_p_O_FDE));
  p_O_FDE desc767(.Q(in_a_r_reg_1[4:4]),.D(out_Q_r[28:28]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc767_p_O_FDE));
  p_O_FDE desc768(.Q(in_a_r_reg_1[5:5]),.D(out_Q_r[29:29]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc768_p_O_FDE));
  p_O_FDE desc769(.Q(in_a_r_reg_1[6:6]),.D(out_Q_r[30:30]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc769_p_O_FDE));
  p_O_FDE desc770(.Q(in_a_r_reg_1[7:7]),.D(out_Q_r[31:31]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc770_p_O_FDE));
  p_O_FDE desc771(.Q(in_a_r_reg_1[8:8]),.D(out_Q_r[32:32]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc771_p_O_FDE));
  p_O_FDE desc772(.Q(in_a_r_reg_1[9:9]),.D(out_Q_r[33:33]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc772_p_O_FDE));
  p_O_FDE desc773(.Q(in_a_r_reg_1[10:10]),.D(out_Q_r[34:34]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc773_p_O_FDE));
  p_O_FDE desc774(.Q(in_a_r_reg_1_11),.D(out_Q_r[35:35]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc774_p_O_FDE));
  p_O_FDE desc775(.Q(in_a_r_reg_0_0),.D(out_Q_r[36:36]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc775_p_O_FDE));
  p_O_FDE desc776(.Q(in_a_r_reg_0[1:1]),.D(out_Q_r[37:37]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc776_p_O_FDE));
  p_O_FDE desc777(.Q(in_a_r_reg_0[2:2]),.D(out_Q_r[38:38]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc777_p_O_FDE));
  p_O_FDE desc778(.Q(in_a_r_reg_0[3:3]),.D(out_Q_r[39:39]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc778_p_O_FDE));
  p_O_FDE desc779(.Q(in_a_r_reg_0[4:4]),.D(out_Q_r[40:40]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc779_p_O_FDE));
  p_O_FDE desc780(.Q(in_a_r_reg_0[5:5]),.D(out_Q_r[41:41]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc780_p_O_FDE));
  p_O_FDE desc781(.Q(in_a_r_reg_0[6:6]),.D(out_Q_r[42:42]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc781_p_O_FDE));
  p_O_FDE desc782(.Q(in_a_r_reg_0[7:7]),.D(out_Q_r[43:43]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc782_p_O_FDE));
  p_O_FDE desc783(.Q(in_a_r_reg_0[8:8]),.D(out_Q_r[44:44]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc783_p_O_FDE));
  p_O_FDE desc784(.Q(in_a_r_reg_0[9:9]),.D(out_Q_r[45:45]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc784_p_O_FDE));
  p_O_FDE desc785(.Q(in_a_r_reg_0[10:10]),.D(out_Q_r[46:46]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc785_p_O_FDE));
  p_O_FDE desc786(.Q(in_a_r_reg_0_11),.D(out_Q_r[47:47]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc786_p_O_FDE));
  p_O_FDE desc787(.Q(in_a_i_reg_3[0:0]),.D(out_Q_i[0:0]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc787_p_O_FDE));
  p_O_FDE desc788(.Q(in_a_i_reg_3[1:1]),.D(out_Q_i[1:1]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc788_p_O_FDE));
  p_O_FDE desc789(.Q(in_a_i_reg_3[2:2]),.D(out_Q_i[2:2]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc789_p_O_FDE));
  p_O_FDE desc790(.Q(in_a_i_reg_3[3:3]),.D(out_Q_i[3:3]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc790_p_O_FDE));
  p_O_FDE desc791(.Q(in_a_i_reg_3[4:4]),.D(out_Q_i[4:4]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc791_p_O_FDE));
  p_O_FDE desc792(.Q(in_a_i_reg_3[5:5]),.D(out_Q_i[5:5]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc792_p_O_FDE));
  p_O_FDE desc793(.Q(in_a_i_reg_3[6:6]),.D(out_Q_i[6:6]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc793_p_O_FDE));
  p_O_FDE desc794(.Q(in_a_i_reg_3[7:7]),.D(out_Q_i[7:7]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc794_p_O_FDE));
  p_O_FDE desc795(.Q(in_a_i_reg_3[8:8]),.D(out_Q_i[8:8]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc795_p_O_FDE));
  p_O_FDE desc796(.Q(in_a_i_reg_3[9:9]),.D(out_Q_i[9:9]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc796_p_O_FDE));
  p_O_FDE desc797(.Q(in_a_i_reg_3[10:10]),.D(out_Q_i[10:10]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc797_p_O_FDE));
  p_O_FDE desc798(.Q(in_a_i_reg_3_11),.D(out_Q_i[11:11]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc798_p_O_FDE));
  p_O_FDE desc799(.Q(in_a_i_reg_2[0:0]),.D(out_Q_i[12:12]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc799_p_O_FDE));
  p_O_FDE desc800(.Q(in_a_i_reg_2[1:1]),.D(out_Q_i[13:13]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc800_p_O_FDE));
  p_O_FDE desc801(.Q(in_a_i_reg_2[2:2]),.D(out_Q_i[14:14]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc801_p_O_FDE));
  p_O_FDE desc802(.Q(in_a_i_reg_2[3:3]),.D(out_Q_i[15:15]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc802_p_O_FDE));
  p_O_FDE desc803(.Q(in_a_i_reg_2[4:4]),.D(out_Q_i[16:16]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc803_p_O_FDE));
  p_O_FDE desc804(.Q(in_a_i_reg_2[5:5]),.D(out_Q_i[17:17]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc804_p_O_FDE));
  p_O_FDE desc805(.Q(in_a_i_reg_2[6:6]),.D(out_Q_i[18:18]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc805_p_O_FDE));
  p_O_FDE desc806(.Q(in_a_i_reg_2[7:7]),.D(out_Q_i[19:19]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc806_p_O_FDE));
  p_O_FDE desc807(.Q(in_a_i_reg_2[8:8]),.D(out_Q_i[20:20]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc807_p_O_FDE));
  p_O_FDE desc808(.Q(in_a_i_reg_2[9:9]),.D(out_Q_i[21:21]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc808_p_O_FDE));
  p_O_FDE desc809(.Q(in_a_i_reg_2[10:10]),.D(out_Q_i[22:22]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc809_p_O_FDE));
  p_O_FDE desc810(.Q(in_a_i_reg_2_11),.D(out_Q_i[23:23]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc810_p_O_FDE));
  p_O_FDE desc811(.Q(in_a_i_reg_1[0:0]),.D(out_Q_i[24:24]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc811_p_O_FDE));
  p_O_FDE desc812(.Q(in_a_i_reg_1[1:1]),.D(out_Q_i[25:25]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc812_p_O_FDE));
  p_O_FDE desc813(.Q(in_a_i_reg_1[2:2]),.D(out_Q_i[26:26]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc813_p_O_FDE));
  p_O_FDE desc814(.Q(in_a_i_reg_1[3:3]),.D(out_Q_i[27:27]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc814_p_O_FDE));
  p_O_FDE desc815(.Q(in_a_i_reg_1[4:4]),.D(out_Q_i[28:28]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc815_p_O_FDE));
  p_O_FDE desc816(.Q(in_a_i_reg_1[5:5]),.D(out_Q_i[29:29]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc816_p_O_FDE));
  p_O_FDE desc817(.Q(in_a_i_reg_1[6:6]),.D(out_Q_i[30:30]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc817_p_O_FDE));
  p_O_FDE desc818(.Q(in_a_i_reg_1[7:7]),.D(out_Q_i[31:31]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc818_p_O_FDE));
  p_O_FDE desc819(.Q(in_a_i_reg_1[8:8]),.D(out_Q_i[32:32]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc819_p_O_FDE));
  p_O_FDE desc820(.Q(in_a_i_reg_1[9:9]),.D(out_Q_i[33:33]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc820_p_O_FDE));
  p_O_FDE desc821(.Q(in_a_i_reg_1[10:10]),.D(out_Q_i[34:34]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc821_p_O_FDE));
  p_O_FDE desc822(.Q(in_a_i_reg_1_11),.D(out_Q_i[35:35]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc822_p_O_FDE));
  p_O_FDE desc823(.Q(in_a_i_reg_0[0:0]),.D(out_Q_i[36:36]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc823_p_O_FDE));
  p_O_FDE desc824(.Q(in_a_i_reg_0[1:1]),.D(out_Q_i[37:37]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc824_p_O_FDE));
  p_O_FDE desc825(.Q(in_a_i_reg_0[2:2]),.D(out_Q_i[38:38]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc825_p_O_FDE));
  p_O_FDE desc826(.Q(in_a_i_reg_0[3:3]),.D(out_Q_i[39:39]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc826_p_O_FDE));
  p_O_FDE desc827(.Q(in_a_i_reg_0[4:4]),.D(out_Q_i[40:40]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc827_p_O_FDE));
  p_O_FDE desc828(.Q(in_a_i_reg_0[5:5]),.D(out_Q_i[41:41]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc828_p_O_FDE));
  p_O_FDE desc829(.Q(in_a_i_reg_0[6:6]),.D(out_Q_i[42:42]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc829_p_O_FDE));
  p_O_FDE desc830(.Q(in_a_i_reg_0[7:7]),.D(out_Q_i[43:43]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc830_p_O_FDE));
  p_O_FDE desc831(.Q(in_a_i_reg_0[8:8]),.D(out_Q_i[44:44]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc831_p_O_FDE));
  p_O_FDE desc832(.Q(in_a_i_reg_0[9:9]),.D(out_Q_i[45:45]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc832_p_O_FDE));
  p_O_FDE desc833(.Q(in_a_i_reg_0[10:10]),.D(out_Q_i[46:46]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc833_p_O_FDE));
  p_O_FDE desc834(.Q(in_a_i_reg_0_11),.D(out_Q_i[47:47]),.C(clk),.CE(w_in_a_vec_sub),.E(p_desc834_p_O_FDE));
  add_subZ3_inj desc835(.pre_out_10(pre_out[11:11]),.output_iv_0(output_iv[1:1]),.output_iv_1(output_iv[2:2]),.output_iv_9(output_iv[10:10]),.output_iv_8(output_iv[9:9]),.output_iv_6(output_iv[7:7]),.output_iv_7(output_iv[8:8]),.output_iv_2(output_iv[3:3]),.output_iv_3(output_iv[4:4]),.output_iv_4(output_iv[5:5]),.out_r_vec_mult_0(out_r_vec_mult_0[11:0]),.in_a_r_reg_0({in_a_r_reg_0_11,in_a_r_reg_0[10:1],in_a_r_reg_0_0}),.N_500(N_500));
  add_subZ3_1_inj desc836(.pre_out_i_m_8(pre_out_i_m[8:8]),.pre_out_i_m_4(pre_out_i_m[4:4]),.pre_out_i_m_0(pre_out_i_m[0:0]),.out_r_vec_mult_1(out_r_vec_mult_1[11:0]),.in_a_r_reg_1({in_a_r_reg_1_11,in_a_r_reg_1[10:0]}),.pre_out_10(pre_out_0[11:11]),.pre_out_9(pre_out[10:10]),.pre_out_8(pre_out[9:9]),.pre_out_6(pre_out[7:7]),.pre_out_5(pre_out[6:6]),.pre_out_4(pre_out[5:5]),.pre_out_2(pre_out[3:3]),.pre_out_1(pre_out[2:2]),.pre_out_0(pre_out[1:1]),.un5_output(un5_output));
  add_subZ3_2_inj desc837(.out_r_vec_mult_2(out_r_vec_mult_2[11:0]),.in_a_r_reg_2({in_a_r_reg_2_11,in_a_r_reg_2[10:0]}),.pre_out_i_m_6(pre_out_i_m[6:6]),.pre_out_i_m_0(pre_out_i_m_0_0),.pre_out_10(pre_out_1[11:11]),.pre_out_9(pre_out_0[10:10]),.pre_out_8(pre_out_0[9:9]),.pre_out_7(pre_out[8:8]),.pre_out_6(pre_out_0[7:7]),.pre_out_4(pre_out_0[5:5]),.pre_out_3(pre_out[4:4]),.pre_out_2(pre_out_0[3:3]),.pre_out_1(pre_out_0[2:2]),.pre_out_0(pre_out_0[1:1]),.un5_output(un5_output_0));
  add_subZ3_3_inj desc838(.out_r_vec_mult_3(out_r_vec_mult_3[11:0]),.in_a_r_reg_3({in_a_r_reg_3_11,in_a_r_reg_3[10:0]}),.pre_out_i_m({pre_out_i_m[1:1],pre_out_i_m_1}),.pre_out_10(pre_out_2[11:11]),.pre_out_9(pre_out_1[10:10]),.pre_out_8(pre_out_1[9:9]),.pre_out_7(pre_out_0[8:8]),.pre_out_6(pre_out_1[7:7]),.pre_out_5(pre_out_0[6:6]),.pre_out_4(pre_out_1[5:5]),.pre_out_3(pre_out_0[4:4]),.pre_out_2(pre_out_1[3:3]),.pre_out_1(pre_out_1[2:2]),.un5_output(un5_output_1));
  add_subZ3_4_inj desc839(.pre_out_10(pre_out_3_9),.output_iv({output_iv_0_9,output_iv_0_8,output_iv_0_7,output_iv_0_6,output_iv[6:6],output_iv_0_4,output_iv_0_3,output_iv_0_2,output_iv_0_1,output_iv_0_0,output_iv[0:0]}),.out_i_vec_sub_0(out_i_vec_sub_0[11:11]),.out_i_vec_mult_0(out_i_vec_mult_0[11:0]),.in_a_i_reg_0({in_a_i_reg_0_11,in_a_i_reg_0[10:0]}));
  add_subZ3_5_inj desc840(.pre_out_i_m(pre_out_i_m_2),.out_i_vec_mult_1(out_i_vec_mult_1[11:0]),.in_a_i_reg_1({in_a_i_reg_1_11,in_a_i_reg_1[10:0]}),.pre_out({pre_out_4[11:11],pre_out_2[10:9],pre_out_1[8:8],pre_out_2[7:7],pre_out_1[6:6],pre_out_2[5:5],pre_out_1[4:4],pre_out_2[3:2],pre_out_1[1:1]}),.un5_output(un5_output_2));
  add_subZ3_6_inj desc841(.pre_out_i_m(pre_out_i_m_3),.out_i_vec_mult_2(out_i_vec_mult_2[11:0]),.in_a_i_reg_2({in_a_i_reg_2_11,in_a_i_reg_2[10:0]}),.pre_out({pre_out_5[11:11],pre_out_3_8,pre_out_3_7,pre_out_2[8:8],pre_out_3_5,pre_out_2[6:6],pre_out_3_3,pre_out_2[4:4],pre_out_3_1,pre_out_3_0,pre_out_2[1:1]}),.un5_output(un5_output_3));
  add_subZ3_7_inj desc842(.out_i_vec_mult_3(out_i_vec_mult_3[11:0]),.in_a_i_reg_3({in_a_i_reg_3_11,in_a_i_reg_3[10:0]}),.pre_out_i_m_1(pre_out_i_m_0_1),.pre_out_i_m_5(pre_out_i_m[5:5]),.pre_out_i_m_2(pre_out_i_m[2:2]),.pre_out_i_m_10(pre_out_i_m[10:10]),.pre_out_i_m_9(pre_out_i_m[9:9]),.pre_out_i_m_6(pre_out_i_m_0_6),.pre_out_i_m_7(pre_out_i_m[7:7]),.pre_out_i_m_3(pre_out_i_m[3:3]),.pre_out_i_m_4(pre_out_i_m_0_4),.pre_out_i_m_0(pre_out_i_m_4),.pre_out_10(pre_out_6[11:11]),.pre_out_7(pre_out_3_6),.un5_output(un5_output_4));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
endmodule
