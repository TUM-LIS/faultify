`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[18:0] testVector;
output[18:0] resultVector;
input[345:0] injectionVector;
IIR_Biquad_inj toplevel_instance (
.clk(clk),
.n_reset(rst),
.sample_trig(testVector[0]),
.X_in(testVector [18:1]),
.filter_done(resultVector[0]),
.Y_out(resultVector [18:1]),
.p_desc86_p_O_FDE(injectionVector[0]),
.p_desc87_p_O_FDE(injectionVector[1]),
.p_desc88_p_O_FDE(injectionVector[2]),
.p_desc89_p_O_FDE(injectionVector[3]),
.p_desc90_p_O_FDE(injectionVector[4]),
.p_desc91_p_O_FDE(injectionVector[5]),
.p_desc92_p_O_FDE(injectionVector[6]),
.p_desc93_p_O_FDE(injectionVector[7]),
.p_desc94_p_O_FDE(injectionVector[8]),
.p_desc95_p_O_FDE(injectionVector[9]),
.p_desc96_p_O_FDE(injectionVector[10]),
.p_desc97_p_O_FDE(injectionVector[11]),
.p_desc98_p_O_FDE(injectionVector[12]),
.p_desc99_p_O_FDE(injectionVector[13]),
.p_desc100_p_O_FDE(injectionVector[14]),
.p_desc101_p_O_FDE(injectionVector[15]),
.p_desc102_p_O_FDE(injectionVector[16]),
.p_desc103_p_O_FDE(injectionVector[17]),
.p_desc104_p_O_FDE(injectionVector[18]),
.p_desc105_p_O_FDE(injectionVector[19]),
.p_desc106_p_O_FDE(injectionVector[20]),
.p_desc107_p_O_FDE(injectionVector[21]),
.p_desc108_p_O_FDE(injectionVector[22]),
.p_desc109_p_O_FDE(injectionVector[23]),
.p_desc110_p_O_FDE(injectionVector[24]),
.p_desc111_p_O_FDE(injectionVector[25]),
.p_desc112_p_O_FDE(injectionVector[26]),
.p_desc113_p_O_FDE(injectionVector[27]),
.p_desc114_p_O_FDE(injectionVector[28]),
.p_desc115_p_O_FDE(injectionVector[29]),
.p_desc116_p_O_FDE(injectionVector[30]),
.p_desc117_p_O_FDE(injectionVector[31]),
.p_desc118_p_O_FDE(injectionVector[32]),
.p_desc119_p_O_FDE(injectionVector[33]),
.p_desc120_p_O_FDE(injectionVector[34]),
.p_desc121_p_O_FDE(injectionVector[35]),
.p_desc162_p_O_FDE(injectionVector[36]),
.p_desc163_p_O_FDE(injectionVector[37]),
.p_desc164_p_O_FDE(injectionVector[38]),
.p_desc165_p_O_FDE(injectionVector[39]),
.p_desc166_p_O_FDE(injectionVector[40]),
.p_desc167_p_O_FDE(injectionVector[41]),
.p_desc168_p_O_FDE(injectionVector[42]),
.p_desc169_p_O_FDE(injectionVector[43]),
.p_desc170_p_O_FDE(injectionVector[44]),
.p_desc171_p_O_FDE(injectionVector[45]),
.p_desc172_p_O_FDE(injectionVector[46]),
.p_desc173_p_O_FDE(injectionVector[47]),
.p_desc174_p_O_FDE(injectionVector[48]),
.p_desc175_p_O_FDE(injectionVector[49]),
.p_desc176_p_O_FDE(injectionVector[50]),
.p_desc177_p_O_FDE(injectionVector[51]),
.p_desc178_p_O_FDE(injectionVector[52]),
.p_desc179_p_O_FDE(injectionVector[53]),
.p_desc198_p_O_FDE(injectionVector[54]),
.p_desc199_p_O_FDE(injectionVector[55]),
.p_desc200_p_O_FDE(injectionVector[56]),
.p_desc201_p_O_FDE(injectionVector[57]),
.p_desc202_p_O_FDE(injectionVector[58]),
.p_desc203_p_O_FDE(injectionVector[59]),
.p_desc204_p_O_FDE(injectionVector[60]),
.p_desc205_p_O_FDE(injectionVector[61]),
.p_desc206_p_O_FDE(injectionVector[62]),
.p_desc207_p_O_FDE(injectionVector[63]),
.p_desc208_p_O_FDE(injectionVector[64]),
.p_desc209_p_O_FDE(injectionVector[65]),
.p_desc210_p_O_FDE(injectionVector[66]),
.p_desc211_p_O_FDE(injectionVector[67]),
.p_desc212_p_O_FDE(injectionVector[68]),
.p_desc213_p_O_FDE(injectionVector[69]),
.p_desc214_p_O_FDE(injectionVector[70]),
.p_desc215_p_O_FDE(injectionVector[71]),
.p_desc216_p_O_FDE(injectionVector[72]),
.p_desc217_p_O_FDE(injectionVector[73]),
.p_desc218_p_O_FDE(injectionVector[74]),
.p_desc219_p_O_FDE(injectionVector[75]),
.p_desc220_p_O_FDE(injectionVector[76]),
.p_desc221_p_O_FDE(injectionVector[77]),
.p_desc222_p_O_FDE(injectionVector[78]),
.p_desc223_p_O_FDE(injectionVector[79]),
.p_desc224_p_O_FDE(injectionVector[80]),
.p_desc225_p_O_FDE(injectionVector[81]),
.p_desc226_p_O_FDE(injectionVector[82]),
.p_desc227_p_O_FDE(injectionVector[83]),
.p_desc228_p_O_FDE(injectionVector[84]),
.p_desc229_p_O_FDE(injectionVector[85]),
.p_desc230_p_O_FDE(injectionVector[86]),
.p_desc231_p_O_FDE(injectionVector[87]),
.p_desc232_p_O_FDE(injectionVector[88]),
.p_desc233_p_O_FDE(injectionVector[89]),
.p_desc234_p_O_FDE(injectionVector[90]),
.p_desc235_p_O_FDE(injectionVector[91]),
.p_desc236_p_O_FDE(injectionVector[92]),
.p_desc237_p_O_FDE(injectionVector[93]),
.p_desc238_p_O_FDE(injectionVector[94]),
.p_desc239_p_O_FDE(injectionVector[95]),
.p_desc240_p_O_FDE(injectionVector[96]),
.p_desc241_p_O_FDE(injectionVector[97]),
.p_desc242_p_O_FDE(injectionVector[98]),
.p_desc243_p_O_FDE(injectionVector[99]),
.p_desc244_p_O_FDE(injectionVector[100]),
.p_desc245_p_O_FDE(injectionVector[101]),
.p_desc246_p_O_FDE(injectionVector[102]),
.p_desc247_p_O_FDE(injectionVector[103]),
.p_desc248_p_O_FDE(injectionVector[104]),
.p_desc249_p_O_FDE(injectionVector[105]),
.p_desc250_p_O_FDE(injectionVector[106]),
.p_desc251_p_O_FDE(injectionVector[107]),
.p_desc252_p_O_FDE(injectionVector[108]),
.p_desc253_p_O_FDE(injectionVector[109]),
.p_desc254_p_O_FDE(injectionVector[110]),
.p_desc255_p_O_FDE(injectionVector[111]),
.p_desc256_p_O_FDE(injectionVector[112]),
.p_desc257_p_O_FDE(injectionVector[113]),
.p_desc258_p_O_FDE(injectionVector[114]),
.p_desc259_p_O_FDE(injectionVector[115]),
.p_desc260_p_O_FDE(injectionVector[116]),
.p_desc261_p_O_FDE(injectionVector[117]),
.p_desc262_p_O_FDE(injectionVector[118]),
.p_desc263_p_O_FDE(injectionVector[119]),
.p_desc264_p_O_FDE(injectionVector[120]),
.p_desc334_p_O_FDC(injectionVector[121]),
.p_desc335_p_O_FDC(injectionVector[122]),
.p_desc336_p_O_FDC(injectionVector[123]),
.p_desc337_p_O_FDC(injectionVector[124]),
.p_state_reg_ret_5_Z_p_O_FDC(injectionVector[125]),
.p_state_reg_ret_Z_p_O_FDP(injectionVector[126]),
.p_state_reg_ret_1_Z_p_O_FDP(injectionVector[127]),
.p_state_reg_ret_2_Z_p_O_FDP(injectionVector[128]),
.p_state_reg_ret_4_Z_p_O_FDP(injectionVector[129]),
.p_desc180_p_O_FDCE(injectionVector[130]),
.p_desc181_p_O_FDCE(injectionVector[131]),
.p_desc182_p_O_FDCE(injectionVector[132]),
.p_desc183_p_O_FDCE(injectionVector[133]),
.p_desc184_p_O_FDCE(injectionVector[134]),
.p_desc185_p_O_FDCE(injectionVector[135]),
.p_desc186_p_O_FDCE(injectionVector[136]),
.p_desc187_p_O_FDCE(injectionVector[137]),
.p_desc188_p_O_FDCE(injectionVector[138]),
.p_desc189_p_O_FDCE(injectionVector[139]),
.p_desc190_p_O_FDCE(injectionVector[140]),
.p_desc191_p_O_FDCE(injectionVector[141]),
.p_desc192_p_O_FDCE(injectionVector[142]),
.p_desc193_p_O_FDCE(injectionVector[143]),
.p_desc194_p_O_FDCE(injectionVector[144]),
.p_desc195_p_O_FDCE(injectionVector[145]),
.p_desc196_p_O_FDCE(injectionVector[146]),
.p_desc197_p_O_FDCE(injectionVector[147]),
.p_desc265_p_O_FDCE(injectionVector[148]),
.p_desc266_p_O_FDCE(injectionVector[149]),
.p_desc267_p_O_FDCE(injectionVector[150]),
.p_desc268_p_O_FDCE(injectionVector[151]),
.p_desc269_p_O_FDCE(injectionVector[152]),
.p_desc270_p_O_FDCE(injectionVector[153]),
.p_desc271_p_O_FDCE(injectionVector[154]),
.p_desc272_p_O_FDCE(injectionVector[155]),
.p_desc273_p_O_FDCE(injectionVector[156]),
.p_desc274_p_O_FDCE(injectionVector[157]),
.p_desc275_p_O_FDCE(injectionVector[158]),
.p_desc276_p_O_FDCE(injectionVector[159]),
.p_desc277_p_O_FDCE(injectionVector[160]),
.p_desc278_p_O_FDCE(injectionVector[161]),
.p_desc279_p_O_FDCE(injectionVector[162]),
.p_desc280_p_O_FDCE(injectionVector[163]),
.p_desc281_p_O_FDCE(injectionVector[164]),
.p_desc282_p_O_FDCE(injectionVector[165]),
.p_desc283_p_O_FDCE(injectionVector[166]),
.p_desc284_p_O_FDCE(injectionVector[167]),
.p_desc285_p_O_FDCE(injectionVector[168]),
.p_desc286_p_O_FDCE(injectionVector[169]),
.p_desc287_p_O_FDCE(injectionVector[170]),
.p_desc288_p_O_FDCE(injectionVector[171]),
.p_desc289_p_O_FDCE(injectionVector[172]),
.p_desc290_p_O_FDCE(injectionVector[173]),
.p_desc291_p_O_FDCE(injectionVector[174]),
.p_desc292_p_O_FDCE(injectionVector[175]),
.p_desc293_p_O_FDCE(injectionVector[176]),
.p_desc294_p_O_FDCE(injectionVector[177]),
.p_desc295_p_O_FDCE(injectionVector[178]),
.p_desc296_p_O_FDCE(injectionVector[179]),
.p_desc297_p_O_FDCE(injectionVector[180]),
.p_desc298_p_O_FDCE(injectionVector[181]),
.p_desc299_p_O_FDCE(injectionVector[182]),
.p_desc300_p_O_FDCE(injectionVector[183]),
.p_desc301_p_O_FDCE(injectionVector[184]),
.p_desc302_p_O_FDCE(injectionVector[185]),
.p_desc303_p_O_FDCE(injectionVector[186]),
.p_desc304_p_O_FDCE(injectionVector[187]),
.p_desc305_p_O_FDCE(injectionVector[188]),
.p_desc306_p_O_FDCE(injectionVector[189]),
.p_desc307_p_O_FDCE(injectionVector[190]),
.p_desc308_p_O_FDCE(injectionVector[191]),
.p_desc309_p_O_FDCE(injectionVector[192]),
.p_desc310_p_O_FDCE(injectionVector[193]),
.p_desc311_p_O_FDCE(injectionVector[194]),
.p_desc312_p_O_FDCE(injectionVector[195]),
.p_desc313_p_O_FDCE(injectionVector[196]),
.p_desc314_p_O_FDCE(injectionVector[197]),
.p_desc315_p_O_FDCE(injectionVector[198]),
.p_desc316_p_O_FDCE(injectionVector[199]),
.p_desc317_p_O_FDCE(injectionVector[200]),
.p_desc318_p_O_FDCE(injectionVector[201]),
.p_desc319_p_O_FDCE(injectionVector[202]),
.p_desc320_p_O_FDCE(injectionVector[203]),
.p_desc321_p_O_FDCE(injectionVector[204]),
.p_desc322_p_O_FDCE(injectionVector[205]),
.p_desc323_p_O_FDCE(injectionVector[206]),
.p_desc324_p_O_FDCE(injectionVector[207]),
.p_desc325_p_O_FDCE(injectionVector[208]),
.p_desc326_p_O_FDCE(injectionVector[209]),
.p_desc327_p_O_FDCE(injectionVector[210]),
.p_desc328_p_O_FDCE(injectionVector[211]),
.p_desc329_p_O_FDCE(injectionVector[212]),
.p_desc330_p_O_FDCE(injectionVector[213]),
.p_desc331_p_O_FDCE(injectionVector[214]),
.p_desc332_p_O_FDCE(injectionVector[215]),
.p_desc333_p_O_FDCE(injectionVector[216]),
.p_desc338_p_O_FDCE(injectionVector[217]),
.p_ZFF_Y1_0_rep1_Z_p_O_FDCE(injectionVector[218]),
.p_desc339_p_O_FDCE(injectionVector[219]),
.p_ZFF_Y1_15_rep1_Z_p_O_FDCE(injectionVector[220]),
.p_desc340_p_O_FDCE(injectionVector[221]),
.p_ZFF_X0_7_rep1_Z_p_O_FDCE(injectionVector[222]),
.p_desc341_p_O_FDCE(injectionVector[223]),
.p_desc342_p_O_FDCE(injectionVector[224]),
.p_desc343_p_O_FDCE(injectionVector[225]),
.p_desc344_p_O_FDCE(injectionVector[226]),
.p_ZFF_Y1_16_rep1_Z_p_O_FDCE(injectionVector[227]),
.p_desc345_p_O_FDCE(injectionVector[228]),
.p_ZFF_X0_6_rep1_Z_p_O_FDCE(injectionVector[229]),
.p_desc346_p_O_FDCE(injectionVector[230]),
.p_desc347_p_O_FDCE(injectionVector[231]),
.p_ZFF_Y1_2_rep1_Z_p_O_FDCE(injectionVector[232]),
.p_desc348_p_O_FDCE(injectionVector[233]),
.p_desc349_p_O_FDCE(injectionVector[234]),
.p_ZFF_X0_10_rep1_Z_p_O_FDCE(injectionVector[235]),
.p_desc350_p_O_FDCE(injectionVector[236]),
.p_ZFF_X0_11_rep1_Z_p_O_FDCE(injectionVector[237]),
.p_desc351_p_O_FDCE(injectionVector[238]),
.p_ZFF_X0_12_rep1_Z_p_O_FDCE(injectionVector[239]),
.p_desc352_p_O_FDCE(injectionVector[240]),
.p_ZFF_X2_6_rep1_Z_p_O_FDCE(injectionVector[241]),
.p_desc353_p_O_FDCE(injectionVector[242]),
.p_ZFF_X0_4_rep1_Z_p_O_FDCE(injectionVector[243]),
.p_desc354_p_O_FDCE(injectionVector[244]),
.p_desc355_p_O_FDCE(injectionVector[245]),
.p_desc356_p_O_FDCE(injectionVector[246]),
.p_desc357_p_O_FDCE(injectionVector[247]),
.p_ZFF_X2_10_rep1_Z_p_O_FDCE(injectionVector[248]),
.p_desc358_p_O_FDCE(injectionVector[249]),
.p_ZFF_X0_2_rep1_Z_p_O_FDCE(injectionVector[250]),
.p_desc359_p_O_FDCE(injectionVector[251]),
.p_ZFF_X0_1_rep1_Z_p_O_FDCE(injectionVector[252]),
.p_desc360_p_O_FDCE(injectionVector[253]),
.p_ZFF_Y1_1_rep1_Z_p_O_FDCE(injectionVector[254]),
.p_desc361_p_O_FDCE(injectionVector[255]),
.p_desc362_p_O_FDCE(injectionVector[256]),
.p_desc363_p_O_FDCE(injectionVector[257]),
.p_desc364_p_O_FDCE(injectionVector[258]),
.p_ZFF_X2_2_rep1_Z_p_O_FDCE(injectionVector[259]),
.p_desc365_p_O_FDCE(injectionVector[260]),
.p_ZFF_X0_3_rep1_Z_p_O_FDCE(injectionVector[261]),
.p_desc366_p_O_FDCE(injectionVector[262]),
.p_desc367_p_O_FDCE(injectionVector[263]),
.p_ZFF_X2_3_rep1_Z_p_O_FDCE(injectionVector[264]),
.p_desc368_p_O_FDCE(injectionVector[265]),
.p_ZFF_Y1_4_rep1_Z_p_O_FDCE(injectionVector[266]),
.p_desc369_p_O_FDCE(injectionVector[267]),
.p_desc370_p_O_FDCE(injectionVector[268]),
.p_ZFF_Y1_3_rep1_Z_p_O_FDCE(injectionVector[269]),
.p_desc371_p_O_FDCE(injectionVector[270]),
.p_desc372_p_O_FDCE(injectionVector[271]),
.p_desc373_p_O_FDCE(injectionVector[272]),
.p_ZFF_Y1_5_rep1_Z_p_O_FDCE(injectionVector[273]),
.p_desc374_p_O_FDCE(injectionVector[274]),
.p_ZFF_X2_14_rep1_Z_p_O_FDCE(injectionVector[275]),
.p_desc375_p_O_FDCE(injectionVector[276]),
.p_ZFF_X0_14_rep1_Z_p_O_FDCE(injectionVector[277]),
.p_desc376_p_O_FDCE(injectionVector[278]),
.p_ZFF_X0_15_rep1_Z_p_O_FDCE(injectionVector[279]),
.p_desc377_p_O_FDCE(injectionVector[280]),
.p_ZFF_X2_15_rep1_Z_p_O_FDCE(injectionVector[281]),
.p_desc378_p_O_FDCE(injectionVector[282]),
.p_ZFF_Y1_6_rep1_Z_p_O_FDCE(injectionVector[283]),
.p_desc379_p_O_FDCE(injectionVector[284]),
.p_ZFF_Y1_13_rep1_Z_p_O_FDCE(injectionVector[285]),
.p_desc380_p_O_FDCE(injectionVector[286]),
.p_ZFF_Y1_7_rep1_Z_p_O_FDCE(injectionVector[287]),
.p_desc381_p_O_FDCE(injectionVector[288]),
.p_ZFF_Y1_14_rep1_Z_p_O_FDCE(injectionVector[289]),
.p_desc382_p_O_FDCE(injectionVector[290]),
.p_ZFF_X1_3_rep1_Z_p_O_FDCE(injectionVector[291]),
.p_desc383_p_O_FDCE(injectionVector[292]),
.p_ZFF_X1_0_rep1_Z_p_O_FDCE(injectionVector[293]),
.p_desc384_p_O_FDCE(injectionVector[294]),
.p_ZFF_Y1_9_rep1_Z_p_O_FDCE(injectionVector[295]),
.p_desc385_p_O_FDCE(injectionVector[296]),
.p_ZFF_X1_7_rep1_Z_p_O_FDCE(injectionVector[297]),
.p_desc386_p_O_FDCE(injectionVector[298]),
.p_ZFF_X1_4_rep1_Z_p_O_FDCE(injectionVector[299]),
.p_desc387_p_O_FDCE(injectionVector[300]),
.p_ZFF_X1_1_rep1_Z_p_O_FDCE(injectionVector[301]),
.p_desc388_p_O_FDCE(injectionVector[302]),
.p_ZFF_Y1_10_rep1_Z_p_O_FDCE(injectionVector[303]),
.p_desc389_p_O_FDCE(injectionVector[304]),
.p_ZFF_X1_8_rep1_Z_p_O_FDCE(injectionVector[305]),
.p_desc390_p_O_FDCE(injectionVector[306]),
.p_ZFF_X1_9_rep1_Z_p_O_FDCE(injectionVector[307]),
.p_desc391_p_O_FDCE(injectionVector[308]),
.p_ZFF_X1_11_rep1_Z_p_O_FDCE(injectionVector[309]),
.p_desc392_p_O_FDCE(injectionVector[310]),
.p_ZFF_X1_15_rep1_Z_p_O_FDCE(injectionVector[311]),
.p_desc393_p_O_FDCE(injectionVector[312]),
.p_ZFF_X1_2_rep1_Z_p_O_FDCE(injectionVector[313]),
.p_desc394_p_O_FDCE(injectionVector[314]),
.p_ZFF_Y1_12_rep1_Z_p_O_FDCE(injectionVector[315]),
.p_desc395_p_O_FDCE(injectionVector[316]),
.p_ZFF_X0_16_rep1_Z_p_O_FDCE(injectionVector[317]),
.p_desc396_p_O_FDCE(injectionVector[318]),
.p_desc397_p_O_FDCE(injectionVector[319]),
.p_ZFF_Y1_17_rep1_Z_p_O_FDCE(injectionVector[320]),
.p_desc398_p_O_FDCE(injectionVector[321]),
.p_ZFF_X1_5_rep1_Z_p_O_FDCE(injectionVector[322]),
.p_desc399_p_O_FDCE(injectionVector[323]),
.p_ZFF_Y1_8_rep1_Z_p_O_FDCE(injectionVector[324]),
.p_desc400_p_O_FDCE(injectionVector[325]),
.p_desc401_p_O_FDCE(injectionVector[326]),
.p_desc402_p_O_FDCE(injectionVector[327]),
.p_ZFF_X1_6_rep1_Z_p_O_FDCE(injectionVector[328]),
.p_desc403_p_O_FDCE(injectionVector[329]),
.p_ZFF_X1_12_rep1_Z_p_O_FDCE(injectionVector[330]),
.p_desc404_p_O_FDCE(injectionVector[331]),
.p_ZFF_X1_10_rep1_Z_p_O_FDCE(injectionVector[332]),
.p_desc405_p_O_FDCE(injectionVector[333]),
.p_ZFF_X1_13_rep1_Z_p_O_FDCE(injectionVector[334]),
.p_desc406_p_O_FDCE(injectionVector[335]),
.p_ZFF_Y1_11_rep1_Z_p_O_FDCE(injectionVector[336]),
.p_desc407_p_O_FDCE(injectionVector[337]),
.p_ZFF_Y2_8_rep1_Z_p_O_FDCE(injectionVector[338]),
.p_desc408_p_O_FDCE(injectionVector[339]),
.p_desc409_p_O_FDCE(injectionVector[340]),
.p_ZFF_Y2_6_rep1_Z_p_O_FDCE(injectionVector[341]),
.p_desc410_p_O_FDCE(injectionVector[342]),
.p_ZFF_Y2_7_rep1_Z_p_O_FDCE(injectionVector[343]),
.p_desc411_p_O_FDCE(injectionVector[344]),
.p_ZFF_Y2_14_rep1_Z_p_O_FDCE(injectionVector[345]));
endmodule