module pre_norm_addsub_inj (pre_norm_sqrt_fracta_o_0,pre_norm_sqrt_fracta_o_18,s_exp_10_o_0,s_exp_10_o,prenorm_addsub_exp_o,v_count_56_0_2,v_count_1_0_1,v_count_1_0_2,s_opa_i,s_opb_i,v_count,v_count_i,pre_norm_div_dvdnd_8,pre_norm_div_dvdnd_9,pre_norm_div_dvdnd_0,pre_norm_div_dvdnd_4,prenorm_addsub_fractb_28_o,prenorm_addsub_fracta_28_o,s_expa_lt_expb,N_1084_i,N_41,N_43,N_1628,N_1630,N_1264,N_46,N_1236,N_70,N_1624,N_53,N_1242,N_1257_i,N_1077,N_1083,un2_s_snan_o_20,N_1051,N_1050,N_987,un4_s_expb_in_2_i_0_e,N_378_i,N_2103,m46_0_e,clk_i,un4_s_expb_in_2_i_o2_2_lut6_2_O5,N_1232_i,N_2220,un4_s_expb_in_2_i_o2_2,un4_s_expb_in_2_i_o2_0,un4_s_expb_in_2_i_o2_1,result_1_i_o3,result_i_o3_lut6_2_O6,N_2240,N_399,N_396,N_1227,N_48_0,N_59,un1_s_infb,result_2_10,un2_s_snan_o_22,un2_s_snan_o_8,un4_s_infa_1,un4_s_infa,N_1041,N_1170,un3_s_snan_o_0,N_1241,N_30_0,N_38_0,N_1617,N_1238,N_27_0,N_1245,N_143_mux,N_1140);
output pre_norm_sqrt_fracta_o_0 ;
output pre_norm_sqrt_fracta_o_18 ;
input s_exp_10_o_0 ;
output s_exp_10_o ;
output [7:0] prenorm_addsub_exp_o ;
input [4:4] v_count_56_0_2 ;
input v_count_1_0_1 ;
input v_count_1_0_2 ;
input [30:0] s_opa_i ;
input [30:0] s_opb_i ;
input [4:0] v_count ;
input v_count_i ;
output pre_norm_div_dvdnd_8 ;
output pre_norm_div_dvdnd_9 ;
output pre_norm_div_dvdnd_0 ;
output pre_norm_div_dvdnd_4 ;
output [26:0] prenorm_addsub_fractb_28_o ;
output [26:0] prenorm_addsub_fracta_28_o ;
output s_expa_lt_expb ;
input N_1084_i ;
input N_41 ;
input N_43 ;
input N_1628 ;
input N_1630 ;
output N_1264 ;
input N_46 ;
output N_1236 ;
output N_70 ;
input N_1624 ;
input N_53 ;
output N_1242 ;
output N_1257_i ;
input N_1077 ;
input N_1083 ;
output un2_s_snan_o_20 ;
output N_1051 ;
output N_1050 ;
output N_987 ;
output un4_s_expb_in_2_i_0_e ;
output N_378_i ;
input N_2103 ;
output m46_0_e ;
input clk_i ;
input un4_s_expb_in_2_i_o2_2_lut6_2_O5 ;
input N_1232_i ;
input N_2220 ;
input un4_s_expb_in_2_i_o2_2 ;
input un4_s_expb_in_2_i_o2_0 ;
input un4_s_expb_in_2_i_o2_1 ;
input result_1_i_o3 ;
input result_i_o3_lut6_2_O6 ;
output N_2240 ;
input N_399 ;
input N_396 ;
input N_1227 ;
output N_48_0 ;
input N_59 ;
output un1_s_infb ;
input result_2_10 ;
input un2_s_snan_o_22 ;
input un2_s_snan_o_8 ;
input un4_s_infa_1 ;
output un4_s_infa ;
input N_1041 ;
input N_1170 ;
output un3_s_snan_o_0 ;
output N_1241 ;
output N_30_0 ;
output N_38_0 ;
input N_1617 ;
output N_1238 ;
output N_27_0 ;
output N_1245 ;
output N_143_mux ;
input N_1140 ;
wire pre_norm_sqrt_fracta_o_0 ;
wire pre_norm_sqrt_fracta_o_18 ;
wire pre_norm_div_dvdnd_8 ;
wire pre_norm_div_dvdnd_9 ;
wire pre_norm_div_dvdnd_0 ;
wire pre_norm_div_dvdnd_4 ;
wire s_expa_lt_expb ;
wire N_1084_i ;
wire N_41 ;
wire N_43 ;
wire N_1628 ;
wire N_1630 ;
wire N_1264 ;
wire N_46 ;
wire N_1236 ;
wire N_70 ;
wire N_1624 ;
wire N_53 ;
wire N_1242 ;
wire N_1257_i ;
wire N_1077 ;
wire N_1083 ;
wire un2_s_snan_o_20 ;
wire N_1051 ;
wire N_1050 ;
wire N_987 ;
wire un4_s_expb_in_2_i_0_e ;
wire N_378_i ;
wire N_2103 ;
wire m46_0_e ;
wire clk_i ;
wire un4_s_expb_in_2_i_o2_2_lut6_2_O5 ;
wire N_1232_i ;
wire N_2220 ;
wire un4_s_expb_in_2_i_o2_2 ;
wire un4_s_expb_in_2_i_o2_0 ;
wire un4_s_expb_in_2_i_o2_1 ;
wire result_1_i_o3 ;
wire result_i_o3_lut6_2_O6 ;
wire N_2240 ;
wire N_399 ;
wire N_396 ;
wire N_1227 ;
wire N_48_0 ;
wire N_59 ;
wire un1_s_infb ;
wire result_2_10 ;
wire un2_s_snan_o_22 ;
wire un2_s_snan_o_8 ;
wire un4_s_infa_1 ;
wire un4_s_infa ;
wire N_1041 ;
wire N_1170 ;
wire un3_s_snan_o_0 ;
wire N_1241 ;
wire N_30_0 ;
wire N_38_0 ;
wire N_1617 ;
wire N_1238 ;
wire N_27_0 ;
wire N_1245 ;
wire N_143_mux ;
wire N_1140 ;
wire [7:0] s_exp_diff ;
wire [4:0] v_count_56_0 ;
wire [4:0] v_count_56_1 ;
wire [4:4] s_fractb_28_o_i_o4_RNIN0MT_O5 ;
wire v_count_56_1_0_2 ;
wire [7:5] un27_0_i_m3_lut6_2_O6 ;
wire [7:5] un27_0_i_m3_lut6_2_O5 ;
wire [7:7] un1_opa_i_i_m3_lut6_2_O6 ;
wire [7:0] s_exp_o ;
wire un27_0_i_m3 ;
wire [26:3] s_fractb_28_o ;
wire [25:11] s_fractb_28_o_i_m3 ;
wire [19:8] s_fractb_28_o_i_m2 ;
wire [19:8] s_fracta_28_o_i_m2 ;
wire [21:3] s_fracta_28_o ;
wire [25:11] s_fracta_28_o_i_m3 ;
wire [5:5] s_fracta_28_o_i_m4 ;
wire [4:0] un5_s_sticky_0_cry ;
wire [4:0] un5_s_sticky_1_cry ;
wire [4:0] s_expa_lt_expb_cry ;
wire s_mux_diff ;
wire v_count_56_1_3_tz ;
wire v_count_0_0_0 ;
wire v_count_0_0_0_1 ;
wire [7:7] un27 ;
wire [7:0] un1_opa_i_3_5 ;
wire [7:7] un1_opa_i_2_i ;
wire v_count_56_1_5_tz ;
wire [7:0] un1_opa_i_3_4 ;
wire v_count_56_1_0_3 ;
wire v_count_56_1_1 ;
wire [1:1] s_fract_shr_28 ;
wire GND ;
wire VCC ;
wire un5_s_sticky_0_df0 ;
wire un5_s_sticky_0_lt0 ;
wire N_194_i ;
wire un5_s_sticky_0_df2 ;
wire un5_s_sticky_0_lt2 ;
wire un5_s_sticky_0_df4 ;
wire un5_s_sticky_0_lt4 ;
wire un5_s_sticky_0_df6 ;
wire un5_s_sticky_0_lt6 ;
wire un5_s_sticky_1_df0 ;
wire un5_s_sticky_1_lt0 ;
wire N_64_mux ;
wire un5_s_sticky_1_df2 ;
wire un5_s_sticky_1_lt2 ;
wire un5_s_sticky_1_df4 ;
wire un5_s_sticky_1_lt4 ;
wire un5_s_sticky_1_df6 ;
wire un5_s_sticky_1_lt6 ;
wire s_expa_lt_expb_df0 ;
wire s_expa_lt_expb_lt0 ;
wire s_expa_lt_expb_df2 ;
wire s_expa_lt_expb_lt2 ;
wire s_expa_lt_expb_df4 ;
wire s_expa_lt_expb_lt4 ;
wire s_expa_lt_expb_df6 ;
wire s_expa_lt_expb_lt6 ;
wire N_2107 ;
wire N_1139 ;
wire N_2129_i ;
wire N_67 ;
wire N_33_0 ;
wire N_26_0 ;
wire N_1249 ;
wire N_1217 ;
wire N_2118 ;
wire N_70_0 ;
wire N_78 ;
wire OUT13_1 ;
wire N_2119 ;
wire N_22 ;
wire N_24 ;
wire N_26 ;
wire N_106 ;
wire N_45 ;
wire N_49 ;
wire N_53_0 ;
wire N_17 ;
wire N_1043 ;
wire N_23 ;
wire N_25 ;
wire N_1057 ;
wire N_989 ;
wire N_51 ;
wire N_11 ;
wire N_13 ;
wire N_995 ;
wire N_39 ;
wire N_1137 ;
wire N_168_2 ;
wire N_5 ;
wire N_7 ;
wire N_9 ;
wire N_2095 ;
wire N_33 ;
wire N_21 ;
wire N_15 ;
wire N_17_0 ;
wire N_43_0 ;
wire N_19 ;
wire N_8 ;
wire N_10 ;
wire N_47 ;
wire N_36 ;
wire N_4 ;
wire N_6 ;
wire N_35 ;
wire N_32 ;
wire N_138 ;
wire N_2180 ;
wire N_2254 ;
wire un3_s_fracta_28_o_0_o4_3_0 ;
wire N_1159 ;
wire N_255 ;
wire N_1286 ;
wire N_2197 ;
wire N_1294 ;
wire N_2242 ;
wire N_227 ;
wire N_1230 ;
wire OVER ;
wire N_163 ;
wire N_164 ;
wire N_254 ;
wire N_1596 ;
wire N_267 ;
wire N_1604 ;
wire N_757 ;
wire N_761 ;
wire N_244 ;
wire N_2234 ;
wire N_1053 ;
wire N_60_mux ;
wire N_1138 ;
wire un1_opa_i_3_4_axb_1 ;
wire s_expa_lt_expb_i ;
wire un1_opa_i_3_s_6 ;
wire un1_opa_i_3_s_7 ;
wire un1_opa_i_3_axb_0 ;
wire un1_opa_i_3_s_1 ;
wire un1_opa_i_3_s_2 ;
wire un1_opa_i_3_s_3 ;
wire un1_opa_i_3_s_4 ;
wire un1_opa_i_3_s_5 ;
wire N_2223_i ;
wire N_2225_i ;
wire N_2229_i ;
wire N_2122_i ;
wire N_1231_i ;
wire un5_s_sticky0 ;
wire un5_s_sticky1 ;
wire un1_opa_i_3_5_axb_1 ;
wire N_2253 ;
wire N_119 ;
wire N_103 ;
wire N_87 ;
wire fractb_28_oc ;
wire N_1666 ;
wire N_1633_1 ;
wire N_1636 ;
wire N_1023 ;
wire N_1195 ;
wire N_243 ;
wire un1_opa_i_3_5_axb_7 ;
wire N_1054 ;
wire un1_opa_i_3_5_axb_5 ;
wire un1_opa_i_3_5_axb_3 ;
wire un1_opa_i_3_5_axb_4 ;
wire un1_opa_i_3_5_axb_2 ;
wire un1_opa_i_3_5_axb_6 ;
wire N_74 ;
wire N_992 ;
wire N_72 ;
wire N_66 ;
wire un1_opa_i_3_4_axb_5 ;
wire un1_opa_i_3_4_axb_3 ;
wire un1_opa_i_3_4_axb_4 ;
wire un1_opa_i_3_4_axb_2 ;
wire N_1277 ;
wire N_168_5 ;
wire un1_opa_i_3_axb_7 ;
wire un1_opa_i_3_axb_6 ;
wire un1_opa_i_3_axb_5 ;
wire un1_opa_i_3_axb_4 ;
wire un1_opa_i_3_axb_3 ;
wire un1_opa_i_3_axb_2 ;
wire un1_opa_i_3_axb_1 ;
wire N_168_2_0_1 ;
wire un3_s_fracta_28_o_0_o4_2_2 ;
wire un3_s_fracta_28_o_0_o4_2_1 ;
wire un3_s_fracta_28_o_0_o4_1_1 ;
wire un3_s_fracta_28_o_0_o4_0_1 ;
wire N_1107_i ;
wire N_251_2 ;
wire N_2173 ;
wire N_1665 ;
wire N_2210 ;
wire N_12 ;
wire N_14 ;
wire N_16 ;
wire N_18 ;
wire N_20 ;
wire un3_s_fracta_28_o_0_o4_2_3 ;
wire un3_s_fracta_28_o_0_o4_1_3 ;
wire un3_s_fracta_28_o_0_o4_0_3 ;
wire un3_s_fracta_28_o_0_o4_3 ;
wire N_168_1_0 ;
wire N_168_2_0 ;
wire N_169_0_2 ;
wire N_169_1 ;
wire un3_s_fracta_28_o_0_o4_1 ;
wire N_31 ;
wire N_229 ;
wire N_2212 ;
wire N_247 ;
wire un3_s_fracta_28_o_0_o4_2_4 ;
wire un3_s_fracta_28_o_0_o4_1_4 ;
wire N_1022 ;
wire N_169_0 ;
wire N_154_1 ;
wire N_115 ;
wire N_988 ;
wire N_68 ;
wire N_69 ;
wire N_2096 ;
wire N_194_1 ;
wire N_1224 ;
wire N_88 ;
wire N_116 ;
wire N_131_mux ;
wire N_169_2 ;
wire un1_opa_i_3_4_axb_7 ;
wire N_2125 ;
wire N_2243 ;
wire N_1024 ;
wire N_168_0 ;
wire N_2217 ;
wire N_52 ;
wire N_2141 ;
wire N_1177 ;
wire N_77 ;
wire N_76 ;
wire N_2224 ;
wire N_104 ;
wire N_2199_1 ;
wire N_1239 ;
wire N_129_mux ;
wire un3_s_fracta_28_o ;
wire N_1240 ;
wire N_1267 ;
wire N_1292 ;
wire N_1108_i ;
wire N_1109_i ;
wire N_1110_i ;
wire N_1111_i ;
wire N_1112_i ;
wire N_1113_i ;
wire un1_opa_i_3_4_axb_6 ;
wire un1_opa_i_3_cry_6 ;
wire un1_opa_i_3_cry_5 ;
wire un1_opa_i_3_cry_4 ;
wire un1_opa_i_3_cry_3 ;
wire un1_opa_i_3_cry_2 ;
wire un1_opa_i_3_cry_1 ;
wire un1_opa_i_3_cry_0 ;
wire un1_opa_i_3_4_cry_6 ;
wire un1_opa_i_3_4_cry_5 ;
wire un1_opa_i_3_4_cry_4 ;
wire un1_opa_i_3_4_cry_3 ;
wire un1_opa_i_3_4_cry_2 ;
wire un1_opa_i_3_4_cry_1 ;
wire un1_opa_i_3_4_cry_0 ;
wire un1_opa_i_3_5_cry_6 ;
wire un1_opa_i_3_5_cry_5 ;
wire un1_opa_i_3_5_cry_4 ;
wire un1_opa_i_3_5_cry_3 ;
wire un1_opa_i_3_5_cry_2 ;
wire un1_opa_i_3_5_cry_1 ;
wire un1_opa_i_3_5_cry_0 ;
wire N_3393 ;
// instances
  LUT6_2 desc0(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_22),.I3(N_24),.I4(N_26),.I5(s_exp_diff[3:3]),.O6(N_106),.O5(N_78));
defparam desc0.INIT=64'h0000000076325410;
  LUT6_2 desc1(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(N_23),.I3(N_25),.I4(N_1057),.I5(s_exp_diff[2:2]),.O6(N_989),.O5(N_51));
defparam desc1.INIT=64'h00001111FC30FC30;
  LUT6_2 desc2(.I0(s_exp_diff[1:1]),.I1(N_5),.I2(N_7),.I3(N_9),.I4(N_11),.I5(s_exp_diff[2:2]),.O6(N_2095),.O5(N_33));
defparam desc2.INIT=64'hFFAA5500E4E4E4E4;
  LUT5 m46_0_e_c(.I0(N_2103),.I1(v_count[1:1]),.I2(v_count[2:2]),.I3(v_count[3:3]),.I4(v_count[4:4]),.O(m46_0_e));
defparam m46_0_e_c.INIT=32'h00000002;
  LUT4 un1_opa_i_3_4_axb_1_cZ(.I0(N_1137),.I1(N_1138),.I2(s_expa_lt_expb),.I3(s_opb_i[24:24]),.O(un1_opa_i_3_4_axb_1));
defparam un1_opa_i_3_4_axb_1_cZ.INIT=16'hE0AE;
  INV desc3(.I(s_expa_lt_expb),.O(s_expa_lt_expb_i));
  FD desc4(.Q(s_exp_diff[6:6]),.D(un1_opa_i_3_s_6),.C(clk_i));
  FD desc5(.Q(s_exp_diff[7:7]),.D(un1_opa_i_3_s_7),.C(clk_i));
  FD desc6(.Q(s_exp_o[7:7]),.D(un27_0_i_m3),.C(clk_i));
  FD desc7(.Q(prenorm_addsub_exp_o[0:0]),.D(s_exp_o[0:0]),.C(clk_i));
  FD desc8(.Q(prenorm_addsub_exp_o[1:1]),.D(s_exp_o[1:1]),.C(clk_i));
  FD desc9(.Q(prenorm_addsub_exp_o[2:2]),.D(s_exp_o[2:2]),.C(clk_i));
  FD desc10(.Q(prenorm_addsub_exp_o[3:3]),.D(s_exp_o[3:3]),.C(clk_i));
  FD desc11(.Q(prenorm_addsub_exp_o[4:4]),.D(s_exp_o[4:4]),.C(clk_i));
  FD desc12(.Q(prenorm_addsub_exp_o[5:5]),.D(s_exp_o[5:5]),.C(clk_i));
  FD desc13(.Q(prenorm_addsub_exp_o[6:6]),.D(s_exp_o[6:6]),.C(clk_i));
  FD desc14(.Q(prenorm_addsub_exp_o[7:7]),.D(s_exp_o[7:7]),.C(clk_i));
  FD desc15(.Q(s_exp_diff[0:0]),.D(un1_opa_i_3_axb_0),.C(clk_i));
  FD desc16(.Q(s_exp_diff[1:1]),.D(un1_opa_i_3_s_1),.C(clk_i));
  FD desc17(.Q(s_exp_diff[2:2]),.D(un1_opa_i_3_s_2),.C(clk_i));
  FD desc18(.Q(s_exp_diff[3:3]),.D(un1_opa_i_3_s_3),.C(clk_i));
  FD desc19(.Q(s_exp_diff[4:4]),.D(un1_opa_i_3_s_4),.C(clk_i));
  FD desc20(.Q(s_exp_diff[5:5]),.D(un1_opa_i_3_s_5),.C(clk_i));
  FD desc21(.Q(s_exp_o[0:0]),.D(un27_0_i_m3_lut6_2_O6[7:7]),.C(clk_i));
  FD desc22(.Q(s_exp_o[1:1]),.D(un27_0_i_m3_lut6_2_O5[7:7]),.C(clk_i));
  FD desc23(.Q(s_exp_o[2:2]),.D(un27_0_i_m3_lut6_2_O6[5:5]),.C(clk_i));
  FD desc24(.Q(s_exp_o[3:3]),.D(un27_0_i_m3_lut6_2_O5[5:5]),.C(clk_i));
  FD desc25(.Q(s_exp_o[4:4]),.D(un4_s_expb_in_2_i_o2_2_lut6_2_O5),.C(clk_i));
  FD desc26(.Q(s_exp_o[5:5]),.D(N_163),.C(clk_i));
  FD desc27(.Q(s_exp_o[6:6]),.D(N_164),.C(clk_i));
  FD desc28(.Q(prenorm_addsub_fractb_28_o[21:21]),.D(s_fractb_28_o[21:21]),.C(clk_i));
  FD desc29(.Q(prenorm_addsub_fractb_28_o[22:22]),.D(s_fractb_28_o[22:22]),.C(clk_i));
  FD desc30(.Q(prenorm_addsub_fractb_28_o[23:23]),.D(s_fractb_28_o[23:23]),.C(clk_i));
  FD desc31(.Q(prenorm_addsub_fractb_28_o[24:24]),.D(s_fractb_28_o_i_m3[24:24]),.C(clk_i));
  FD desc32(.Q(prenorm_addsub_fractb_28_o[25:25]),.D(s_fractb_28_o_i_m3[25:25]),.C(clk_i));
  FD desc33(.Q(prenorm_addsub_fractb_28_o[26:26]),.D(s_fractb_28_o[26:26]),.C(clk_i));
  FD desc34(.Q(prenorm_addsub_fractb_28_o[6:6]),.D(s_fractb_28_o[6:6]),.C(clk_i));
  FD desc35(.Q(prenorm_addsub_fractb_28_o[7:7]),.D(s_fractb_28_o[7:7]),.C(clk_i));
  FD desc36(.Q(prenorm_addsub_fractb_28_o[8:8]),.D(s_fractb_28_o_i_m2[8:8]),.C(clk_i));
  FD desc37(.Q(prenorm_addsub_fractb_28_o[9:9]),.D(s_fractb_28_o_i_m2[9:9]),.C(clk_i));
  FD desc38(.Q(prenorm_addsub_fractb_28_o[10:10]),.D(s_fractb_28_o[10:10]),.C(clk_i));
  FD desc39(.Q(prenorm_addsub_fractb_28_o[11:11]),.D(s_fractb_28_o_i_m3[11:11]),.C(clk_i));
  FD desc40(.Q(prenorm_addsub_fractb_28_o[12:12]),.D(s_fractb_28_o[12:12]),.C(clk_i));
  FD desc41(.Q(prenorm_addsub_fractb_28_o[13:13]),.D(s_fractb_28_o[13:13]),.C(clk_i));
  FD desc42(.Q(prenorm_addsub_fractb_28_o[14:14]),.D(s_fractb_28_o[14:14]),.C(clk_i));
  FD desc43(.Q(prenorm_addsub_fractb_28_o[15:15]),.D(N_1232_i),.C(clk_i));
  FD desc44(.Q(prenorm_addsub_fractb_28_o[16:16]),.D(s_fractb_28_o[16:16]),.C(clk_i));
  FD desc45(.Q(prenorm_addsub_fractb_28_o[17:17]),.D(s_fractb_28_o[17:17]),.C(clk_i));
  FD desc46(.Q(prenorm_addsub_fractb_28_o[18:18]),.D(s_fractb_28_o[18:18]),.C(clk_i));
  FD desc47(.Q(prenorm_addsub_fractb_28_o[19:19]),.D(s_fractb_28_o_i_m2[19:19]),.C(clk_i));
  FD desc48(.Q(prenorm_addsub_fractb_28_o[20:20]),.D(s_fractb_28_o[20:20]),.C(clk_i));
  FD desc49(.Q(prenorm_addsub_fracta_28_o[19:19]),.D(s_fracta_28_o_i_m2[19:19]),.C(clk_i));
  FD desc50(.Q(prenorm_addsub_fracta_28_o[20:20]),.D(N_2223_i),.C(clk_i));
  FD desc51(.Q(prenorm_addsub_fracta_28_o[21:21]),.D(s_fracta_28_o[21:21]),.C(clk_i));
  FD desc52(.Q(prenorm_addsub_fracta_28_o[22:22]),.D(N_2225_i),.C(clk_i));
  FD desc53(.Q(prenorm_addsub_fracta_28_o[23:23]),.D(N_2229_i),.C(clk_i));
  FD desc54(.Q(prenorm_addsub_fracta_28_o[24:24]),.D(s_fracta_28_o_i_m3[24:24]),.C(clk_i));
  FD desc55(.Q(prenorm_addsub_fracta_28_o[25:25]),.D(s_fracta_28_o_i_m3[25:25]),.C(clk_i));
  FD desc56(.Q(prenorm_addsub_fractb_28_o[3:3]),.D(s_fractb_28_o[3:3]),.C(clk_i));
  FD desc57(.Q(prenorm_addsub_fractb_28_o[4:4]),.D(N_2129_i),.C(clk_i));
  FD desc58(.Q(prenorm_addsub_fractb_28_o[5:5]),.D(N_2122_i),.C(clk_i));
  FD desc59(.Q(prenorm_addsub_fracta_28_o[4:4]),.D(s_fractb_28_o_i_o4_RNIN0MT_O5[4:4]),.C(clk_i));
  FD desc60(.Q(prenorm_addsub_fracta_28_o[5:5]),.D(s_fracta_28_o_i_m4[5:5]),.C(clk_i));
  FD desc61(.Q(prenorm_addsub_fracta_28_o[6:6]),.D(s_fracta_28_o[6:6]),.C(clk_i));
  FD desc62(.Q(prenorm_addsub_fracta_28_o[7:7]),.D(s_fracta_28_o[7:7]),.C(clk_i));
  FD desc63(.Q(prenorm_addsub_fracta_28_o[8:8]),.D(s_fracta_28_o_i_m2[8:8]),.C(clk_i));
  FD desc64(.Q(prenorm_addsub_fracta_28_o[9:9]),.D(s_fracta_28_o_i_m2[9:9]),.C(clk_i));
  FD desc65(.Q(prenorm_addsub_fracta_28_o[10:10]),.D(s_fracta_28_o[10:10]),.C(clk_i));
  FD desc66(.Q(prenorm_addsub_fracta_28_o[11:11]),.D(s_fracta_28_o_i_m3[11:11]),.C(clk_i));
  FD desc67(.Q(prenorm_addsub_fracta_28_o[12:12]),.D(s_fracta_28_o[12:12]),.C(clk_i));
  FD desc68(.Q(prenorm_addsub_fracta_28_o[13:13]),.D(s_fracta_28_o[13:13]),.C(clk_i));
  FD desc69(.Q(prenorm_addsub_fracta_28_o[14:14]),.D(s_fracta_28_o[14:14]),.C(clk_i));
  FD desc70(.Q(prenorm_addsub_fracta_28_o[15:15]),.D(N_1231_i),.C(clk_i));
  FD desc71(.Q(prenorm_addsub_fracta_28_o[16:16]),.D(s_fracta_28_o[16:16]),.C(clk_i));
  FD desc72(.Q(prenorm_addsub_fracta_28_o[17:17]),.D(s_fracta_28_o[17:17]),.C(clk_i));
  FD desc73(.Q(prenorm_addsub_fracta_28_o[18:18]),.D(s_fracta_28_o[18:18]),.C(clk_i));
  FD desc74(.Q(prenorm_addsub_fracta_28_o[3:3]),.D(s_fracta_28_o[3:3]),.C(clk_i));
  MUXCY desc75(.DI(un5_s_sticky_0_lt6),.CI(un5_s_sticky_0_cry[4:4]),.S(un5_s_sticky_0_df6),.O(un5_s_sticky0));
  MUXCY desc76(.DI(un5_s_sticky_1_lt6),.CI(un5_s_sticky_1_cry[4:4]),.S(un5_s_sticky_1_df6),.O(un5_s_sticky1));
  MUXCY desc77(.DI(s_expa_lt_expb_lt6),.CI(s_expa_lt_expb_cry[4:4]),.S(s_expa_lt_expb_df6),.O(s_expa_lt_expb));
  LUT5 desc78(.I0(s_opb_i[24:24]),.I1(s_opa_i[24:24]),.I2(N_1077),.I3(s_expa_lt_expb),.I4(N_1084_i),.O(un1_opa_i_3_5_axb_1));
defparam desc78.INIT=32'hA9CF9A98;
  LUT3 desc79(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(N_1084_i),.O(s_mux_diff));
defparam desc79.INIT=8'hE1;
  LUT6_L un5_s_sticky_1_df0_lut6_2_RNO_4(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[12:12]),.I3(s_opb_i[3:3]),.I4(s_opb_i[1:1]),.I5(s_opb_i[7:7]),.LO(v_count_56_1_3_tz));
defparam un5_s_sticky_1_df0_lut6_2_RNO_4.INIT=64'h00000000000000BA;
  LUT6 m48_e(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[12:12]),.I3(s_opb_i[8:8]),.I4(s_opb_i[9:9]),.I5(N_2220),.O(N_2253));
defparam m48_e.INIT=64'h0000000100000000;
  LUT6_L desc80(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_opb_i[4:4]),.I4(s_expa_lt_expb),.I5(N_119),.LO(s_fractb_28_o[7:7]));
defparam desc80.INIT=64'h0101FF000000FF00;
  LUT6_L desc81(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_opa_i[10:10]),.I4(s_expa_lt_expb),.I5(OUT13_1),.LO(s_fracta_28_o[13:13]));
defparam desc81.INIT=64'hFF000101FF000000;
  LUT6_L desc82(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_opa_i[4:4]),.I4(s_expa_lt_expb),.I5(N_119),.LO(s_fracta_28_o[7:7]));
defparam desc82.INIT=64'hFF000101FF000000;
  LUT6 fracta_28_oc(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_exp_diff[4:4]),.I4(N_103),.I5(N_87),.O(fractb_28_oc));
defparam fracta_28_oc.INIT=64'h0101000101000000;
  LUT6_L desc83(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_opb_i[10:10]),.I4(s_expa_lt_expb),.I5(OUT13_1),.LO(s_fractb_28_o[13:13]));
defparam desc83.INIT=64'h0101FF000000FF00;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_2(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[1:1]),.I3(s_opa_i[4:4]),.I4(s_opa_i[0:0]),.I5(v_count_0_0_0),.LO(v_count_0_0_0_1));
defparam un5_s_sticky_0_df0_lut6_2_RNO_2.INIT=64'hFFFFFFFFFFFF0B0A;
  LUT6 un5_s_sticky_0_df4_lut6_2_RNO(.I0(s_opa_i[12:12]),.I1(s_opa_i[10:10]),.I2(s_opa_i[11:11]),.I3(s_opa_i[0:0]),.I4(v_count_56_0_2[4:4]),.I5(N_254),.O(v_count_56_0[4:4]));
defparam un5_s_sticky_0_df4_lut6_2_RNO.INIT=64'h0001000000000000;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_6(.I0(s_opa_i[12:12]),.I1(s_opa_i[7:7]),.I2(s_opa_i[10:10]),.I3(s_opa_i[11:11]),.I4(s_opa_i[9:9]),.I5(N_1666),.LO(N_1633_1));
defparam un5_s_sticky_0_df0_lut6_2_RNO_6.INIT=64'hCCCCCFCFCCCCCFCE;
  LUT6 un5_s_sticky_0_df0_lut6_2_RNO_0(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[1:1]),.I3(s_opa_i[4:4]),.I4(s_opa_i[0:0]),.I5(N_1636),.O(v_count_56_0[1:1]));
defparam un5_s_sticky_0_df0_lut6_2_RNO_0.INIT=64'hFFFFFFFFFFFF0504;
  LUT6_L desc84(.I0(s_opa_i[21:21]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_53_0),.LO(s_fracta_28_o_i_m3[24:24]));
defparam desc84.INIT=64'hAAAA0003AAAA0000;
  LUT6_L desc85(.I0(s_opb_i[21:21]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_53_0),.LO(s_fractb_28_o_i_m3[24:24]));
defparam desc85.INIT=64'h0003AAAA0000AAAA;
  LUT5 desc86(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(N_4),.O(N_1023));
defparam desc86.INIT=32'h00040000;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_7(.I0(s_opa_i[3:3]),.I1(s_opa_i[7:7]),.I2(s_opa_i[1:1]),.I3(s_opa_i[10:10]),.I4(s_opa_i[9:9]),.I5(s_opa_i[5:5]),.LO(N_1195));
defparam un5_s_sticky_0_df0_lut6_2_RNO_7.INIT=64'h0000000000000100;
  LUT6 desc87(.I0(s_opb_i[24:24]),.I1(s_opb_i[23:23]),.I2(s_opa_i[24:24]),.I3(un4_s_expb_in_2_i_o2_2),.I4(un4_s_expb_in_2_i_o2_0),.I5(un4_s_expb_in_2_i_o2_1),.O(N_1138));
defparam desc87.INIT=64'h0000000000000010;
  LUT6 desc88(.I0(s_opb_i[24:24]),.I1(s_opb_i[23:23]),.I2(un4_s_expb_in_2_i_o2_2),.I3(un4_s_expb_in_2_i_o2_0),.I4(un4_s_expb_in_2_i_o2_1),.I5(s_expa_lt_expb),.O(N_243));
defparam desc88.INIT=64'h0000000100000000;
  LUT6 un1_opa_i_3_4_cry_0_RNO(.I0(s_opb_i[23:23]),.I1(s_opa_i[24:24]),.I2(s_opa_i[23:23]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(un27[7:7]));
defparam un1_opa_i_3_4_cry_0_RNO.INIT=64'hF0F0002200000022;
  LUT6 desc89(.I0(s_opb_i[23:23]),.I1(s_opa_i[24:24]),.I2(s_opa_i[23:23]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(un1_opa_i_3_5[0:0]));
defparam desc89.INIT=64'h55550F0FA595A587;
  LUT6 un1_opa_i_3_5_axb_7_cZ(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(s_opa_i[24:24]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(un1_opa_i_3_5_axb_7));
defparam un1_opa_i_3_5_axb_7_cZ.INIT=64'h5555333399959993;
  LUT6 desc90(.I0(s_opb_i[23:23]),.I1(s_opa_i[24:24]),.I2(s_opa_i[23:23]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(un1_opa_i_2_i[7:7]));
defparam desc90.INIT=64'hFFFFFFFF0F3F5577;
  LUT6 desc91(.I0(s_exp_diff[0:0]),.I1(s_opa_i[24:24]),.I2(s_exp_diff[1:1]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(N_1054));
defparam desc91.INIT=64'h0000050405050504;
  LUT6 desc92(.I0(s_opa_i[28:28]),.I1(s_opb_i[28:28]),.I2(s_opa_i[24:24]),.I3(N_1077),.I4(s_expa_lt_expb),.I5(N_1084_i),.O(un1_opa_i_3_5_axb_5));
defparam desc92.INIT=64'h3333555599939995;
  LUT6 desc93(.I0(s_opa_i[26:26]),.I1(s_opb_i[26:26]),.I2(s_opa_i[24:24]),.I3(result_1_i_o3),.I4(N_1077),.I5(s_expa_lt_expb),.O(un1_opa_i_3_5_axb_3));
defparam desc93.INIT=64'h9933933399559555;
  LUT6 desc94(.I0(s_opa_i[27:27]),.I1(s_opb_i[27:27]),.I2(s_opa_i[24:24]),.I3(result_1_i_o3),.I4(N_1077),.I5(s_expa_lt_expb),.O(un1_opa_i_3_5_axb_4));
defparam desc94.INIT=64'h9933933399559555;
  LUT6 desc95(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(s_opa_i[24:24]),.I3(result_1_i_o3),.I4(N_1077),.I5(s_expa_lt_expb),.O(un1_opa_i_3_5_axb_2));
defparam desc95.INIT=64'h9955955599339333;
  LUT6 desc96(.I0(s_opa_i[29:29]),.I1(s_opb_i[29:29]),.I2(s_opa_i[24:24]),.I3(result_1_i_o3),.I4(N_1077),.I5(s_expa_lt_expb),.O(un1_opa_i_3_5_axb_6));
defparam desc96.INIT=64'h9933933399559555;
  LUT6_L un5_s_sticky_1_df0_lut6_2_RNO_6(.I0(s_opb_i[11:11]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[7:7]),.I4(s_opb_i[16:16]),.I5(N_757),.LO(v_count_56_1_5_tz));
defparam un5_s_sticky_1_df0_lut6_2_RNO_6.INIT=64'h0045004400000000;
  LUT6_L desc97(.I0(s_opa_i[6:6]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_74),.I5(N_992),.LO(s_fracta_28_o_i_m2[9:9]));
defparam desc97.INIT=64'hAA3FAA33AA0CAA00;
  LUT6_L desc98(.I0(s_opb_i[6:6]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_74),.I5(N_992),.LO(s_fractb_28_o_i_m2[9:9]));
defparam desc98.INIT=64'h3FAA33AA0CAA00AA;
  LUT6 desc99(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(s_expa_lt_expb),.I3(N_1084_i),.I4(N_25),.I5(result_i_o3_lut6_2_O6),.O(N_53_0));
defparam desc99.INIT=64'h3777044433730040;
  LUT4_L desc100(.I0(N_987),.I1(result_1_i_o3),.I2(s_expa_lt_expb),.I3(N_2234),.LO(s_fractb_28_o[26:26]));
defparam desc100.INIT=16'h5C0C;
  LUT6 desc101(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(s_exp_diff[3:3]),.I3(N_24),.I4(N_26),.I5(N_72),.O(N_2240));
defparam desc101.INIT=64'h5F4F1F0F50401000;
  LUT6 desc102(.I0(s_exp_diff[4:4]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[1:1]),.I3(OVER),.I4(N_66),.I5(N_26),.O(N_992));
defparam desc102.INIT=64'h0057000200550000;
  LUT5 un1_opa_i_3_4_axb_5_cZ(.I0(s_opa_i[28:28]),.I1(s_opb_i[28:28]),.I2(N_1138),.I3(s_expa_lt_expb),.I4(N_1137),.O(un1_opa_i_3_4_axb_5));
defparam un1_opa_i_3_4_axb_5_cZ.INIT=32'hDD33D030;
  LUT5 un1_opa_i_3_4_axb_3_cZ(.I0(s_opa_i[26:26]),.I1(s_opb_i[26:26]),.I2(N_1138),.I3(s_expa_lt_expb),.I4(N_1137),.O(un1_opa_i_3_4_axb_3));
defparam un1_opa_i_3_4_axb_3_cZ.INIT=32'hDD33D030;
  LUT5 un1_opa_i_3_4_axb_4_cZ(.I0(s_opa_i[27:27]),.I1(s_opb_i[27:27]),.I2(N_1138),.I3(s_expa_lt_expb),.I4(N_1137),.O(un1_opa_i_3_4_axb_4));
defparam un1_opa_i_3_4_axb_4_cZ.INIT=32'hDD33D030;
  LUT5 un1_opa_i_3_4_axb_2_cZ(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(N_1138),.I3(s_expa_lt_expb),.I4(N_1137),.O(un1_opa_i_3_4_axb_2));
defparam un1_opa_i_3_4_axb_2_cZ.INIT=32'hBB55B050;
  LUT6 m117(.I0(s_opa_i[10:10]),.I1(s_opa_i[11:11]),.I2(N_399),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(N_1277));
defparam m117.INIT=64'h5555555555555553;
  LUT5 m83(.I0(N_1227),.I1(v_count[3:3]),.I2(N_48_0),.I3(N_67),.I4(N_59),.O(pre_norm_div_dvdnd_9));
defparam m83.INIT=32'hFDA87520;
  LUT6 un5_s_sticky_1_df2_lut6_2_RNO(.I0(s_opb_i[8:8]),.I1(s_opb_i[0:0]),.I2(N_2220),.I3(N_2254),.I4(N_2242),.I5(N_2253),.O(N_64_mux));
defparam un5_s_sticky_1_df2_lut6_2_RNO.INIT=64'hFF33003350335033;
  LUT6 un1_s_infb_c(.I0(s_opb_i[26:26]),.I1(s_opb_i[29:29]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.I4(N_168_5),.I5(N_168_2),.O(un1_s_infb));
defparam un1_s_infb_c.INIT=64'h8000000000000000;
  LUT2 un1_s_infb_2(.I0(s_opb_i[25:25]),.I1(s_opb_i[24:24]),.O(N_168_5));
defparam un1_s_infb_2.INIT=4'h8;
  LUT2_L un1_opa_i_3_axb_7_cZ(.I0(un1_opa_i_3_5[7:7]),.I1(un1_opa_i_3_4[7:7]),.LO(un1_opa_i_3_axb_7));
defparam un1_opa_i_3_axb_7_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_6_cZ(.I0(un1_opa_i_3_5[6:6]),.I1(un1_opa_i_3_4[6:6]),.LO(un1_opa_i_3_axb_6));
defparam un1_opa_i_3_axb_6_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_5_cZ(.I0(un1_opa_i_3_5[5:5]),.I1(un1_opa_i_3_4[5:5]),.LO(un1_opa_i_3_axb_5));
defparam un1_opa_i_3_axb_5_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_4_cZ(.I0(un1_opa_i_3_5[4:4]),.I1(un1_opa_i_3_4[4:4]),.LO(un1_opa_i_3_axb_4));
defparam un1_opa_i_3_axb_4_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_3_cZ(.I0(un1_opa_i_3_5[3:3]),.I1(un1_opa_i_3_4[3:3]),.LO(un1_opa_i_3_axb_3));
defparam un1_opa_i_3_axb_3_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_2_cZ(.I0(un1_opa_i_3_5[2:2]),.I1(un1_opa_i_3_4[2:2]),.LO(un1_opa_i_3_axb_2));
defparam un1_opa_i_3_axb_2_cZ.INIT=4'h6;
  LUT2_L un1_opa_i_3_axb_1_cZ(.I0(un1_opa_i_3_5[1:1]),.I1(un1_opa_i_3_4[1:1]),.LO(un1_opa_i_3_axb_1));
defparam un1_opa_i_3_axb_1_cZ.INIT=4'h6;
  LUT3_L desc103(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(s_expa_lt_expb),.LO(un27_0_i_m3));
defparam desc103.INIT=8'hCA;
  LUT3 un3_s_snan_o_0_a2_2_1(.I0(s_opb_i[21:21]),.I1(s_opb_i[14:14]),.I2(s_opb_i[22:22]),.O(N_168_2_0_1));
defparam un3_s_snan_o_0_a2_2_1.INIT=8'h01;
  LUT5 un3_s_fracta_28_o_0_o4_2_2_cZ(.I0(s_opb_i[21:21]),.I1(s_opb_i[2:2]),.I2(s_opa_i[2:2]),.I3(s_opa_i[21:21]),.I4(s_expa_lt_expb),.O(un3_s_fracta_28_o_0_o4_2_2));
defparam un3_s_fracta_28_o_0_o4_2_2_cZ.INIT=32'hEEEEFFF0;
  LUT5_L un3_s_fracta_28_o_0_o4_2_1_cZ(.I0(s_opb_i[3:3]),.I1(s_opa_i[3:3]),.I2(s_opb_i[1:1]),.I3(s_opa_i[1:1]),.I4(s_expa_lt_expb),.LO(un3_s_fracta_28_o_0_o4_2_1));
defparam un3_s_fracta_28_o_0_o4_2_1_cZ.INIT=32'hFAFAFFCC;
  LUT5_L un3_s_fracta_28_o_0_o4_1_1_cZ(.I0(s_opa_i[6:6]),.I1(s_opb_i[6:6]),.I2(s_opb_i[9:9]),.I3(s_opa_i[9:9]),.I4(s_expa_lt_expb),.LO(un3_s_fracta_28_o_0_o4_1_1));
defparam un3_s_fracta_28_o_0_o4_1_1_cZ.INIT=32'hFCFCFFAA;
  LUT5_L un3_s_fracta_28_o_0_o4_0_1_cZ(.I0(s_opb_i[13:13]),.I1(s_opb_i[4:4]),.I2(s_opa_i[13:13]),.I3(s_opa_i[4:4]),.I4(s_expa_lt_expb),.LO(un3_s_fracta_28_o_0_o4_0_1));
defparam un3_s_fracta_28_o_0_o4_0_1_cZ.INIT=32'hEEEEFFF0;
  LUT3 un1_opa_i_3_5_cry_0_RNO(.I0(s_opb_i[23:23]),.I1(s_opa_i[23:23]),.I2(s_expa_lt_expb),.O(N_1107_i));
defparam un1_opa_i_3_5_cry_0_RNO.INIT=8'h53;
  LUT6 un5_s_sticky_0_df2_lut6_2_RNO_2(.I0(s_opa_i[16:16]),.I1(s_opa_i[14:14]),.I2(s_opa_i[13:13]),.I3(s_opa_i[19:19]),.I4(s_opa_i[15:15]),.I5(s_opa_i[20:20]),.O(N_251_2));
defparam un5_s_sticky_0_df2_lut6_2_RNO_2.INIT=64'h0000000000000001;
  LUT6 un3_s_fracta_28_o_0_a3(.I0(s_opb_i[0:0]),.I1(s_opa_i[0:0]),.I2(s_exp_diff[0:0]),.I3(s_exp_diff[2:2]),.I4(s_exp_diff[1:1]),.I5(s_expa_lt_expb),.O(N_2173));
defparam un3_s_fracta_28_o_0_a3.INIT=64'h00A0000000C00000;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_9(.I0(s_opa_i[17:17]),.I1(s_opa_i[18:18]),.I2(s_opa_i[19:19]),.I3(s_opa_i[21:21]),.I4(s_opa_i[22:22]),.I5(s_opa_i[20:20]),.LO(N_1665));
defparam un5_s_sticky_0_df0_lut6_2_RNO_9.INIT=64'h1111111110101011;
  LUT6_L un5_s_sticky_1_df0_lut6_2_RNO_8(.I0(s_opb_i[21:21]),.I1(s_opb_i[17:17]),.I2(s_opb_i[19:19]),.I3(s_opb_i[20:20]),.I4(s_opb_i[18:18]),.I5(s_opb_i[22:22]),.LO(N_2210));
defparam un5_s_sticky_1_df0_lut6_2_RNO_8.INIT=64'h0000333000003331;
  LUT6 desc104(.I0(s_opb_i[1:1]),.I1(s_opb_i[0:0]),.I2(s_opa_i[1:1]),.I3(s_opa_i[0:0]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_4));
defparam desc104.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc105(.I0(s_opb_i[2:2]),.I1(s_opa_i[2:2]),.I2(s_opb_i[1:1]),.I3(s_opa_i[1:1]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_5));
defparam desc105.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc106(.I0(s_opb_i[2:2]),.I1(s_opa_i[2:2]),.I2(s_opb_i[3:3]),.I3(s_opa_i[3:3]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_6));
defparam desc106.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6 desc107(.I0(s_opb_i[3:3]),.I1(s_opb_i[4:4]),.I2(s_opa_i[3:3]),.I3(s_opa_i[4:4]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_7));
defparam desc107.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc108(.I0(s_opb_i[4:4]),.I1(s_opb_i[5:5]),.I2(s_opa_i[4:4]),.I3(s_opa_i[5:5]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_8));
defparam desc108.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc109(.I0(s_opa_i[6:6]),.I1(s_opb_i[6:6]),.I2(s_opb_i[5:5]),.I3(s_opa_i[5:5]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_9));
defparam desc109.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6 desc110(.I0(s_opa_i[6:6]),.I1(s_opb_i[6:6]),.I2(s_opb_i[7:7]),.I3(s_opa_i[7:7]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_10));
defparam desc110.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc111(.I0(s_opb_i[8:8]),.I1(s_opb_i[7:7]),.I2(s_opa_i[7:7]),.I3(s_opa_i[8:8]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_11));
defparam desc111.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc112(.I0(s_opb_i[8:8]),.I1(s_opb_i[9:9]),.I2(s_opa_i[8:8]),.I3(s_opa_i[9:9]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_12));
defparam desc112.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc113(.I0(s_opb_i[10:10]),.I1(s_opb_i[9:9]),.I2(s_opa_i[10:10]),.I3(s_opa_i[9:9]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_13));
defparam desc113.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc114(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opa_i[10:10]),.I3(s_opa_i[11:11]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_14));
defparam desc114.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc115(.I0(s_opb_i[11:11]),.I1(s_opb_i[12:12]),.I2(s_opa_i[12:12]),.I3(s_opa_i[11:11]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_15));
defparam desc115.INIT=64'hCCCCAAAAF0F0FF00;
  LUT6 desc116(.I0(s_opb_i[13:13]),.I1(s_opb_i[12:12]),.I2(s_opa_i[12:12]),.I3(s_opa_i[13:13]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_16));
defparam desc116.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc117(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opa_i[14:14]),.I3(s_opa_i[13:13]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_17_0));
defparam desc117.INIT=64'hCCCCAAAAF0F0FF00;
  LUT6 desc118(.I0(s_opb_i[14:14]),.I1(s_opb_i[15:15]),.I2(s_opa_i[14:14]),.I3(s_opa_i[15:15]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_18));
defparam desc118.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc119(.I0(s_opa_i[16:16]),.I1(s_opb_i[15:15]),.I2(s_opa_i[15:15]),.I3(s_opb_i[16:16]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_19));
defparam desc119.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc120(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opb_i[17:17]),.I3(s_opb_i[16:16]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_20));
defparam desc120.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc121(.I0(s_opa_i[17:17]),.I1(s_opb_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opb_i[18:18]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_21));
defparam desc121.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc122(.I0(s_opb_i[19:19]),.I1(s_opa_i[18:18]),.I2(s_opa_i[19:19]),.I3(s_opb_i[18:18]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_22));
defparam desc122.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc123(.I0(s_opb_i[19:19]),.I1(s_opb_i[20:20]),.I2(s_opa_i[19:19]),.I3(s_opa_i[20:20]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_23));
defparam desc123.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc124(.I0(s_opb_i[21:21]),.I1(s_opb_i[20:20]),.I2(s_opa_i[21:21]),.I3(s_opa_i[20:20]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_24));
defparam desc124.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc125(.I0(s_opb_i[21:21]),.I1(s_opa_i[21:21]),.I2(s_opa_i[22:22]),.I3(s_opb_i[22:22]),.I4(s_exp_diff[0:0]),.I5(s_expa_lt_expb),.O(N_25));
defparam desc125.INIT=64'hFF00AAAAF0F0CCCC;
  LUT6 un3_s_fracta_28_o_0_o4_2_3_cZ(.I0(s_opa_i[16:16]),.I1(s_opa_i[18:18]),.I2(s_opb_i[16:16]),.I3(s_opb_i[18:18]),.I4(s_expa_lt_expb),.I5(un3_s_fracta_28_o_0_o4_2_1),.O(un3_s_fracta_28_o_0_o4_2_3));
defparam un3_s_fracta_28_o_0_o4_2_3_cZ.INIT=64'hFFFFFFFFFFF0EEEE;
  LUT6_L un3_s_fracta_28_o_0_o4_1_3_cZ(.I0(s_opb_i[5:5]),.I1(s_opa_i[22:22]),.I2(s_opa_i[5:5]),.I3(s_opb_i[22:22]),.I4(s_expa_lt_expb),.I5(un3_s_fracta_28_o_0_o4_1_1),.LO(un3_s_fracta_28_o_0_o4_1_3));
defparam un3_s_fracta_28_o_0_o4_1_3_cZ.INIT=64'hFFFFFFFFFFAAFCFC;
  LUT6 un3_s_fracta_28_o_0_o4_0_3_cZ(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opa_i[10:10]),.I3(s_opa_i[11:11]),.I4(s_expa_lt_expb),.I5(un3_s_fracta_28_o_0_o4_0_1),.O(un3_s_fracta_28_o_0_o4_0_3));
defparam un3_s_fracta_28_o_0_o4_0_3_cZ.INIT=64'hFFFFFFFFEEEEFFF0;
  LUT6 un3_s_fracta_28_o_0_o4_3_cZ(.I0(s_opb_i[19:19]),.I1(s_opb_i[20:20]),.I2(s_opa_i[19:19]),.I3(s_opa_i[20:20]),.I4(s_expa_lt_expb),.I5(un3_s_fracta_28_o_0_o4_3_0),.O(un3_s_fracta_28_o_0_o4_3));
defparam un3_s_fracta_28_o_0_o4_3_cZ.INIT=64'hFFFFFFFFEEEEFFF0;
  LUT6 un3_s_snan_o_0_a2_1_1(.I0(s_opb_i[10:10]),.I1(s_opb_i[6:6]),.I2(s_opb_i[12:12]),.I3(s_opb_i[8:8]),.I4(s_opb_i[0:0]),.I5(N_168_5),.O(N_168_1_0));
defparam un3_s_snan_o_0_a2_1_1.INIT=64'h0001000000000000;
  LUT6 un3_s_snan_o_0_a2_2(.I0(s_opb_i[2:2]),.I1(s_opb_i[4:4]),.I2(s_opb_i[20:20]),.I3(s_opb_i[16:16]),.I4(N_168_2_0_1),.I5(result_2_10),.O(N_168_2_0));
defparam un3_s_snan_o_0_a2_2.INIT=64'h0000000000010000;
  LUT5_L un3_s_snan_o_0_a2_0_0_2(.I0(s_opa_i[21:21]),.I1(s_opa_i[22:22]),.I2(s_opa_i[20:20]),.I3(un2_s_snan_o_20),.I4(un2_s_snan_o_22),.LO(N_169_0_2));
defparam un3_s_snan_o_0_a2_0_0_2.INIT=32'h01000000;
  LUT6 un3_s_snan_o_0_a2_0_1(.I0(s_opa_i[25:25]),.I1(s_opa_i[27:27]),.I2(s_opa_i[24:24]),.I3(N_1159),.I4(pre_norm_sqrt_fracta_o_0),.I5(un2_s_snan_o_8),.O(N_169_1));
defparam un3_s_snan_o_0_a2_0_1.INIT=64'h0080000000000000;
  LUT6 un4_s_infa_c(.I0(s_opa_i[28:28]),.I1(s_opa_i[29:29]),.I2(s_opa_i[25:25]),.I3(s_opa_i[27:27]),.I4(s_opa_i[23:23]),.I5(un4_s_infa_1),.O(un4_s_infa));
defparam un4_s_infa_c.INIT=64'h8000000000000000;
  LUT6_L un3_s_fracta_28_o_0_o4_1_cZ(.I0(s_opb_i[8:8]),.I1(s_opb_i[7:7]),.I2(s_opa_i[7:7]),.I3(s_opa_i[8:8]),.I4(s_expa_lt_expb),.I5(un3_s_fracta_28_o_0_o4_1_3),.LO(un3_s_fracta_28_o_0_o4_1));
defparam un3_s_fracta_28_o_0_o4_1_cZ.INIT=64'hFFFFFFFFEEEEFFF0;
  LUT3 desc126(.I0(s_exp_diff[1:1]),.I1(N_17_0),.I2(N_19),.O(N_45));
defparam desc126.INIT=8'hE4;
  LUT6 desc127(.I0(s_opb_i[0:0]),.I1(s_opa_i[0:0]),.I2(s_exp_diff[0:0]),.I3(s_exp_diff[1:1]),.I4(s_expa_lt_expb),.I5(N_5),.O(N_31));
defparam desc127.INIT=64'hFFA0FFC000A000C0;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_5(.I0(s_opa_i[6:6]),.I1(s_opa_i[7:7]),.I2(s_opa_i[8:8]),.I3(s_opa_i[5:5]),.I4(N_1217),.I5(N_1195),.LO(v_count_0_0_0));
defparam un5_s_sticky_0_df0_lut6_2_RNO_5.INIT=64'hFFFFFFFF00BA0000;
  LUT6 un5_s_sticky_1_df4_lut6_2_RNO(.I0(s_opb_i[12:12]),.I1(s_opb_i[8:8]),.I2(s_opb_i[9:9]),.I3(N_1041),.I4(N_2220),.I5(N_2254),.O(v_count_56_1[4:4]));
defparam un5_s_sticky_1_df4_lut6_2_RNO.INIT=64'h0100000000000000;
  LUT6_L un5_s_sticky_0_df2_lut6_2_RNO_4(.I0(s_opa_i[8:8]),.I1(s_opa_i[10:10]),.I2(s_opa_i[9:9]),.I3(s_opa_i[5:5]),.I4(N_1596),.I5(un2_s_snan_o_8),.LO(N_229));
defparam un5_s_sticky_0_df2_lut6_2_RNO_4.INIT=64'hFFFFFFFEFFFFFFFF;
  LUT5_L un5_s_sticky_0_df0_lut6_2_RNO_8(.I0(s_opa_i[16:16]),.I1(s_opa_i[14:14]),.I2(s_opa_i[13:13]),.I3(s_opa_i[15:15]),.I4(N_1665),.LO(N_1666));
defparam un5_s_sticky_0_df0_lut6_2_RNO_8.INIT=32'h03030302;
  LUT5_L un5_s_sticky_1_df0_lut6_2_RNO_7(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[16:16]),.I4(N_2210),.LO(N_2212));
defparam un5_s_sticky_1_df0_lut6_2_RNO_7.INIT=32'h11111110;
  LUT5 un5_s_sticky_0_df2_lut6_2_RNO_3(.I0(s_opa_i[16:16]),.I1(s_opa_i[14:14]),.I2(s_opa_i[13:13]),.I3(s_opa_i[15:15]),.I4(N_267),.O(N_247));
defparam un5_s_sticky_0_df2_lut6_2_RNO_3.INIT=32'hFFFE0000;
  LUT6 un3_s_fracta_28_o_0_o4_2_4_cZ(.I0(s_opb_i[0:0]),.I1(s_opa_i[0:0]),.I2(s_expa_lt_expb),.I3(un3_s_fracta_28_o_0_o4_2_2),.I4(un3_s_fracta_28_o_0_o4_2_3),.I5(un3_s_fracta_28_o_0_o4_3),.O(un3_s_fracta_28_o_0_o4_2_4));
defparam un3_s_fracta_28_o_0_o4_2_4_cZ.INIT=64'hFFFFFFFFFFFFFFAC;
  LUT6 un3_s_fracta_28_o_0_o4_1_4_cZ(.I0(s_opa_i[17:17]),.I1(s_opb_i[17:17]),.I2(s_expa_lt_expb),.I3(N_1230),.I4(un3_s_fracta_28_o_0_o4_0_3),.I5(un3_s_fracta_28_o_0_o4_1),.O(un3_s_fracta_28_o_0_o4_1_4));
defparam un3_s_fracta_28_o_0_o4_1_4_cZ.INIT=64'hFFFFFFFFFFFFCAFF;
  LUT6 desc128(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(N_6),.I5(N_8),.O(N_1022));
defparam desc128.INIT=64'h000A000800020000;
  LUT6_L un3_s_snan_o_0_a2_0_0(.I0(s_opa_i[28:28]),.I1(s_opa_i[29:29]),.I2(s_opa_i[26:26]),.I3(s_opa_i[13:13]),.I4(N_1604),.I5(N_169_0_2),.LO(N_169_0));
defparam un3_s_snan_o_0_a2_0_0.INIT=64'h0000008000000000;
  LUT6 un3_s_snan_o_0_a2_1_0(.I0(s_opb_i[13:13]),.I1(s_opb_i[15:15]),.I2(s_opb_i[17:17]),.I3(s_opb_i[9:9]),.I4(s_opb_i[5:5]),.I5(N_761),.O(N_154_1));
defparam un3_s_snan_o_0_a2_1_0.INIT=64'h0000000100000000;
  LUT6 desc129(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_8),.I3(N_10),.I4(N_12),.I5(N_14),.O(N_115));
defparam desc129.INIT=64'hFEBADC9876325410;
  LUT6 desc130(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_21),.I3(N_15),.I4(N_17_0),.I5(N_19),.O(N_988));
defparam desc130.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc131(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_10),.I3(N_12),.I4(N_14),.I5(N_16),.O(N_66));
defparam desc131.INIT=64'hFEBADC9876325410;
  LUT6 desc132(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_12),.I3(N_14),.I4(N_16),.I5(N_18),.O(N_68));
defparam desc132.INIT=64'hFEBADC9876325410;
  LUT6 desc133(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_13),.I3(N_15),.I4(N_17_0),.I5(N_19),.O(N_69));
defparam desc133.INIT=64'hFEBADC9876325410;
  LUT6 desc134(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_14),.I3(N_16),.I4(N_18),.I5(N_20),.O(N_70_0));
defparam desc134.INIT=64'hFEBADC9876325410;
  LUT6 desc135(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_16),.I3(N_18),.I4(N_20),.I5(N_22),.O(N_72));
defparam desc135.INIT=64'hFEBADC9876325410;
  LUT6 desc136(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_18),.I3(N_20),.I4(N_22),.I5(N_24),.O(N_74));
defparam desc136.INIT=64'hFEBADC9876325410;
  LUT6 desc137(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_9),.I3(N_11),.I4(N_13),.I5(N_15),.O(N_2096));
defparam desc137.INIT=64'hFEBADC9876325410;
  LUT6 desc138(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_6),.I3(N_8),.I4(N_10),.I5(N_12),.O(N_2118));
defparam desc138.INIT=64'hFEBADC9876325410;
  LUT6 un5_s_sticky_1_df0_lut6_2_RNO_1(.I0(s_opb_i[8:8]),.I1(s_opb_i[9:9]),.I2(s_opb_i[5:5]),.I3(s_opb_i[7:7]),.I4(N_757),.I5(v_count_56_1_3_tz),.O(v_count_56_1_0_3));
defparam un5_s_sticky_1_df0_lut6_2_RNO_1.INIT=64'h030B0303000A0000;
  LUT6 un5_s_sticky_0_df2_lut6_2_RNO_1(.I0(s_opa_i[17:17]),.I1(s_opa_i[18:18]),.I2(s_opa_i[19:19]),.I3(s_opa_i[20:20]),.I4(s_opa_i[0:0]),.I5(N_267),.O(N_194_1));
defparam un5_s_sticky_0_df2_lut6_2_RNO_1.INIT=64'hFFFF0001FFFF0000;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_4(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opa_i[19:19]),.I4(s_opa_i[15:15]),.I5(N_1170),.LO(N_1224));
defparam un5_s_sticky_0_df0_lut6_2_RNO_4.INIT=64'h0000BABB0000BABA;
  LUT6 un5_s_sticky_1_df2_lut6_2_RNO_0(.I0(s_opb_i[17:17]),.I1(s_opb_i[18:18]),.I2(N_2180),.I3(N_2197),.I4(N_2254),.I5(N_2253),.O(v_count_56_1[3:3]));
defparam un5_s_sticky_1_df2_lut6_2_RNO_0.INIT=64'h01000000FFFF0000;
  LUT6 un5_s_sticky_0_df2_lut6_2_RNO(.I0(s_opa_i[17:17]),.I1(s_opa_i[18:18]),.I2(s_opa_i[0:0]),.I3(N_254),.I4(N_251_2),.I5(N_229),.O(v_count_56_0[3:3]));
defparam un5_s_sticky_0_df2_lut6_2_RNO.INIT=64'h0F000F0001000000;
  LUT5 desc139(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_32),.I3(N_36),.I4(N_68),.O(N_88));
defparam desc139.INIT=32'hFEDC3210;
  LUT6 desc140(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_35),.I3(N_39),.I4(N_47),.I5(N_43_0),.O(N_116));
defparam desc140.INIT=64'hFEDC7654BA983210;
  LUT6 desc141(.I0(s_opa_i[22:22]),.I1(s_opb_i[22:22]),.I2(s_exp_diff[0:0]),.I3(s_expa_lt_expb),.I4(N_1084_i),.I5(result_i_o3_lut6_2_O6),.O(N_26));
defparam desc141.INIT=64'h0CFAFCFA0C0AFC0A;
  LUT6_L m109(.I0(s_opb_i[2:2]),.I1(s_opb_i[6:6]),.I2(s_opb_i[3:3]),.I3(s_opb_i[4:4]),.I4(s_opb_i[5:5]),.I5(N_1286),.LO(N_131_mux));
defparam m109.INIT=64'h3333003033330031;
  LUT6 desc142(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_31),.I3(N_35),.I4(N_39),.I5(N_43_0),.O(N_87));
defparam desc142.INIT=64'hFEDCBA9876543210;
  LUT6_L un5_s_sticky_1_df0_lut6_2_RNO_3(.I0(s_opb_i[13:13]),.I1(s_opb_i[6:6]),.I2(s_opb_i[9:9]),.I3(s_opb_i[5:5]),.I4(N_757),.I5(v_count_56_1_5_tz),.LO(v_count_56_1_1));
defparam un5_s_sticky_1_df0_lut6_2_RNO_3.INIT=64'h00CD000500CC0000;
  LUT6_L un3_s_snan_o_0_a2_0_2(.I0(s_opa_i[30:30]),.I1(s_opa_i[2:2]),.I2(s_opa_i[12:12]),.I3(s_opa_i[1:1]),.I4(s_opa_i[5:5]),.I5(N_169_0),.LO(N_169_2));
defparam un3_s_snan_o_0_a2_0_2.INIT=64'h0000000200000000;
  LUT5 un1_opa_i_3_4_axb_7_cZ(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(N_243),.I3(N_244),.I4(s_mux_diff),.O(un1_opa_i_3_4_axb_7));
defparam un1_opa_i_3_4_axb_7_cZ.INIT=32'h153FEAC0;
  LUT5 un3_s_fracta_28_o_0_m3(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_2173),.I3(N_33),.I4(N_2096),.O(N_2125));
defparam un3_s_fracta_28_o_0_m3.INIT=32'hFEFC3230;
  LUT6 desc143(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_39),.I3(N_51),.I4(N_47),.I5(N_43_0),.O(N_2243));
defparam desc143.INIT=64'h018945CD23AB67EF;
  LUT6 desc144(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(N_45),.I4(N_49),.I5(N_2096),.O(N_1024));
defparam desc144.INIT=64'h0F0B07030C080400;
  LUT6 un3_s_snan_o_0_a2_0(.I0(s_opb_i[26:26]),.I1(s_opb_i[29:29]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.I4(N_168_2),.I5(N_154_1),.O(N_168_0));
defparam un3_s_snan_o_0_a2_0.INIT=64'h8000000000000000;
  LUT5_L un5_s_sticky_1_df0_lut6_2_RNO_5(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[12:12]),.I3(s_opb_i[9:9]),.I4(N_2212),.LO(N_2217));
defparam un5_s_sticky_1_df0_lut6_2_RNO_5.INIT=32'h00550054;
  LUT3 desc145(.I0(s_exp_diff[1:1]),.I1(N_24),.I2(N_26),.O(N_52));
defparam desc145.INIT=8'hE4;
  LUT6 desc146(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(N_1043),.I3(s_expa_lt_expb),.I4(N_1084_i),.I5(result_i_o3_lut6_2_O6),.O(N_2234));
defparam desc146.INIT=64'h0010101000001000;
  LUT6_L un3_s_fracta_28_o_0_a2(.I0(s_expa_lt_expb),.I1(N_1057),.I2(un3_s_fracta_28_o_0_o4_2_4),.I3(un3_s_fracta_28_o_0_o4_1_4),.I4(un5_s_sticky0),.I5(un5_s_sticky1),.LO(N_2141));
defparam un3_s_fracta_28_o_0_a2.INIT=64'hFFF3AAA255510000;
  LUT6 un5_s_sticky_0_df2_lut6_2_RNO_0(.I0(s_opa_i[8:8]),.I1(s_opa_i[5:5]),.I2(un2_s_snan_o_8),.I3(N_254),.I4(N_194_1),.I5(N_247),.O(N_194_i));
defparam un5_s_sticky_0_df2_lut6_2_RNO_0.INIT=64'h00000000000010FF;
  LUT4 un5_s_sticky_0_df0_lut6_2_RNO_1(.I0(s_opa_i[14:14]),.I1(s_opa_i[12:12]),.I2(s_opa_i[13:13]),.I3(N_1224),.O(N_1177));
defparam un5_s_sticky_0_df0_lut6_2_RNO_1.INIT=16'hCFCE;
  LUT6 desc147(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[1:1]),.I3(N_25),.I4(N_1057),.I5(N_49),.O(N_77));
defparam desc147.INIT=64'h3F337F730C004C40;
  LUT5 desc148(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_1054),.I3(N_51),.I4(N_47),.O(N_103));
defparam desc148.INIT=32'h73516240;
  LUT6 desc149(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_20),.I3(N_22),.I4(N_24),.I5(N_26),.O(N_76));
defparam desc149.INIT=64'hFEBADC9876325410;
  LUT6_L un5_s_sticky_0_df0_lut6_2_RNO_3(.I0(s_opa_i[6:6]),.I1(s_opa_i[2:2]),.I2(s_opa_i[8:8]),.I3(s_opa_i[1:1]),.I4(s_opa_i[5:5]),.I5(N_1633_1),.LO(N_1636));
defparam un5_s_sticky_0_df0_lut6_2_RNO_3.INIT=64'h0000001100000010;
  LUT6 un5_s_sticky_1_df0_lut6_2_RNO(.I0(s_opb_i[0:0]),.I1(v_count_56_1_0_2),.I2(N_138),.I3(v_count_56_1_0_3),.I4(N_154_1),.I5(v_count_56_1_1),.O(v_count_56_1[0:0]));
defparam un5_s_sticky_1_df0_lut6_2_RNO.INIT=64'hFFFFFFFFFFFEFFEE;
  LUT6_L desc150(.I0(s_opa_i[22:22]),.I1(s_exp_diff[1:1]),.I2(N_1043),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_26),.LO(s_fracta_28_o_i_m3[25:25]));
defparam desc150.INIT=64'hAAAA0030AAAA0000;
  LUT6_L desc151(.I0(s_opb_i[22:22]),.I1(s_exp_diff[1:1]),.I2(N_1043),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_26),.LO(s_fractb_28_o_i_m3[25:25]));
defparam desc151.INIT=64'h0030AAAA0000AAAA;
  LUT6 desc152(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(s_exp_diff[3:3]),.I3(N_23),.I4(N_25),.I5(N_1054),.O(N_2224));
defparam desc152.INIT=64'h0F0E0B0A05040100;
  LUT6 desc153(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(s_exp_diff[3:3]),.I3(N_20),.I4(N_22),.I5(N_52),.O(N_104));
defparam desc153.INIT=64'h0F0E0B0A05040100;
  LUT5_L un5_s_sticky_1_df0_lut6_2_RNO_2(.I0(s_opb_i[6:6]),.I1(s_opb_i[8:8]),.I2(s_opb_i[5:5]),.I3(s_opb_i[7:7]),.I4(N_2217),.LO(N_2199_1));
defparam un5_s_sticky_1_df0_lut6_2_RNO_2.INIT=32'h05050504;
  LUT6 un5_s_sticky_0_df0_lut6_2_RNO(.I0(s_opa_i[7:7]),.I1(s_opa_i[11:11]),.I2(N_255),.I3(N_1217),.I4(N_1177),.I5(v_count_0_0_0_1),.O(v_count_56_0[0:0]));
defparam un5_s_sticky_0_df0_lut6_2_RNO.INIT=64'hFFFFFFFF10000000;
  LUT6_L desc154(.I0(s_opa_i[5:5]),.I1(N_1043),.I2(N_1053),.I3(s_expa_lt_expb),.I4(N_53_0),.I5(N_1024),.LO(s_fracta_28_o_i_m2[8:8]));
defparam desc154.INIT=64'hAAFFAAFFAAC0AA00;
  LUT6_L desc155(.I0(s_opb_i[5:5]),.I1(N_1043),.I2(N_1053),.I3(s_expa_lt_expb),.I4(N_53_0),.I5(N_1024),.LO(s_fractb_28_o_i_m2[8:8]));
defparam desc155.INIT=64'hFFAAFFAAC0AA00AA;
  LUT5 un3_s_snan_o_0_c(.I0(N_168_1_0),.I1(N_168_2_0),.I2(N_169_1),.I3(N_168_0),.I4(N_169_2),.O(un3_s_snan_o_0));
defparam un3_s_snan_o_0_c.INIT=32'hF8F08800;
  LUT6 desc156(.I0(s_exp_diff[4:4]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[3:3]),.I3(N_115),.I4(N_72),.I5(N_52),.O(N_119));
defparam desc156.INIT=64'h5752070255500500;
  LUT5_L desc157(.I0(s_opa_i[13:13]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_17),.LO(s_fracta_28_o[16:16]));
defparam desc157.INIT=32'hAA00AA03;
  LUT6 m20(.I0(s_opa_i[12:12]),.I1(s_opa_i[13:13]),.I2(N_399),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(N_1239));
defparam m20.INIT=64'h5555555555555553;
  LUT5_L desc158(.I0(s_opb_i[15:15]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_103),.LO(s_fractb_28_o[18:18]));
defparam desc158.INIT=32'h03AA00AA;
  LUT5_L desc159(.I0(s_opa_i[15:15]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_103),.LO(s_fracta_28_o[18:18]));
defparam desc159.INIT=32'hAA03AA00;
  LUT6_L m105_e(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[8:8]),.I3(s_opb_i[9:9]),.I4(s_opb_i[7:7]),.I5(N_131_mux),.LO(N_129_mux));
defparam m105_e.INIT=64'h2232223222322233;
  LUT5_L desc160(.I0(s_opb_i[13:13]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_17),.LO(s_fractb_28_o[16:16]));
defparam desc160.INIT=32'h00AA03AA;
  LUT6_L desc161(.I0(s_opa_i[7:7]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_2234),.I5(N_2243),.LO(s_fracta_28_o[10:10]));
defparam desc161.INIT=64'hAA0CAA00AA0FAA03;
  LUT6_L desc162(.I0(s_opb_i[7:7]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_2234),.I5(N_2243),.LO(s_fractb_28_o[10:10]));
defparam desc162.INIT=64'h0CAA00AA0FAA03AA;
  LUT6 desc163(.I0(s_exp_diff[3:3]),.I1(N_1053),.I2(N_1023),.I3(N_1022),.I4(N_74),.I5(N_992),.O(s_fract_shr_28[1:1]));
defparam desc163.INIT=64'hFFFEFFFAFFF4FFF0;
  LUT6_L desc164(.I0(s_opa_i[18:18]),.I1(s_exp_diff[4:4]),.I2(s_exp_diff[3:3]),.I3(OVER),.I4(s_expa_lt_expb),.I5(N_78),.LO(s_fracta_28_o[21:21]));
defparam desc164.INIT=64'hAAAA0003AAAA0000;
  LUT6_L desc165(.I0(s_opb_i[18:18]),.I1(s_exp_diff[4:4]),.I2(s_exp_diff[3:3]),.I3(OVER),.I4(s_expa_lt_expb),.I5(N_78),.LO(s_fractb_28_o[21:21]));
defparam desc165.INIT=64'h0003AAAA0000AAAA;
  LUT6_L desc166(.I0(s_opa_i[14:14]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_74),.I5(N_995),.LO(s_fracta_28_o[17:17]));
defparam desc166.INIT=64'hAA03AA00AA0FAA0C;
  LUT6_L desc167(.I0(s_opb_i[14:14]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_74),.I5(N_995),.LO(s_fractb_28_o[17:17]));
defparam desc167.INIT=64'h03AA00AA0FAA0CAA;
  LUT5_L desc168(.I0(s_opb_i[17:17]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_77),.LO(s_fractb_28_o[20:20]));
defparam desc168.INIT=32'h03AA00AA;
  LUT5_L desc169(.I0(s_opb_i[19:19]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_989),.LO(s_fractb_28_o[22:22]));
defparam desc169.INIT=32'h03AA00AA;
  LUT6_L desc170(.I0(s_opb_i[20:20]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_52),.LO(s_fractb_28_o[23:23]));
defparam desc170.INIT=64'h0003AAAA0000AAAA;
  LUT6 desc171(.I0(s_exp_diff[4:4]),.I1(s_exp_diff[3:3]),.I2(OVER),.I3(N_2095),.I4(N_69),.I5(N_77),.O(N_2107));
defparam desc171.INIT=64'hF8F9FCFDFAFBFEFF;
  LUT6_L desc172(.I0(s_opa_i[16:16]),.I1(s_exp_diff[4:4]),.I2(s_exp_diff[3:3]),.I3(OVER),.I4(s_expa_lt_expb),.I5(N_76),.LO(s_fracta_28_o_i_m2[19:19]));
defparam desc172.INIT=64'hAAAA0003AAAA0000;
  LUT6_L desc173(.I0(s_opb_i[16:16]),.I1(s_exp_diff[4:4]),.I2(s_exp_diff[3:3]),.I3(OVER),.I4(s_expa_lt_expb),.I5(N_76),.LO(s_fractb_28_o_i_m2[19:19]));
defparam desc173.INIT=64'h0003AAAA0000AAAA;
  LUT5 un3_s_fracta_28_o_0(.I0(s_exp_diff[4:4]),.I1(OVER),.I2(N_2125),.I3(N_17),.I4(N_2141),.O(un3_s_fracta_28_o));
defparam un3_s_fracta_28_o_0.INIT=32'hFFFF1032;
  LUT6 m17(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[4:4]),.I3(s_opa_i[5:5]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_1236));
defparam m17.INIT=64'h55550F0F333300FF;
  LUT5 m22(.I0(s_opa_i[10:10]),.I1(s_opa_i[11:11]),.I2(v_count[1:1]),.I3(N_1239),.I4(v_count_i),.O(N_1240));
defparam m22.INIT=32'h3F305F50;
  LUT6 m25(.I0(s_opa_i[6:6]),.I1(s_opa_i[7:7]),.I2(s_opa_i[8:8]),.I3(s_opa_i[9:9]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_26_0));
defparam m25.INIT=64'h55550F0F333300FF;
  LUT6 m28(.I0(s_opa_i[14:14]),.I1(s_opa_i[12:12]),.I2(s_opa_i[13:13]),.I3(s_opa_i[15:15]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_1241));
defparam m28.INIT=64'h333355550F0F00FF;
  LUT5 m29(.I0(s_opa_i[8:8]),.I1(s_opa_i[9:9]),.I2(v_count[1:1]),.I3(N_1277),.I4(v_count[0:0]),.O(N_30_0));
defparam m29.INIT=32'h5F503F30;
  LUT6 m32(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[14:14]),.I3(s_opa_i[15:15]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_33_0));
defparam m32.INIT=64'h0F0F555500FF3333;
  LUT6 m37(.I0(s_opa_i[6:6]),.I1(s_opa_i[7:7]),.I2(s_opa_i[4:4]),.I3(s_opa_i[5:5]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_38_0));
defparam m37.INIT=64'h0F0F555500FF3333;
  LUT6_L desc174(.I0(s_opa_i[3:3]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_2224),.I5(N_116),.LO(s_fracta_28_o[6:6]));
defparam desc174.INIT=64'hAA0FAA03AA0CAA00;
  LUT6_L desc175(.I0(s_opa_i[8:8]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_68),.I5(N_76),.LO(s_fracta_28_o_i_m3[11:11]));
defparam desc175.INIT=64'hAA0FAA0CAA03AA00;
  LUT6_L desc176(.I0(s_opb_i[8:8]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_68),.I5(N_76),.LO(s_fractb_28_o_i_m3[11:11]));
defparam desc176.INIT=64'h0FAA0CAA03AA00AA;
  LUT6_L desc177(.I0(s_opb_i[11:11]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_988),.I5(N_989),.LO(s_fractb_28_o[14:14]));
defparam desc177.INIT=64'h0FAA0CAA03AA00AA;
  LUT6_L desc178(.I0(s_opa_i[11:11]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_988),.I5(N_989),.LO(s_fracta_28_o[14:14]));
defparam desc178.INIT=64'hAA0FAA0CAA03AA00;
  LUT6_L desc179(.I0(s_opb_i[3:3]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_2224),.I5(N_116),.LO(s_fractb_28_o[6:6]));
defparam desc179.INIT=64'h0FAA03AA0CAA00AA;
  LUT6_L desc180(.I0(s_opb_i[9:9]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_69),.I5(N_77),.LO(s_fractb_28_o[12:12]));
defparam desc180.INIT=64'h0FAA0CAA03AA00AA;
  LUT6_L desc181(.I0(s_opa_i[9:9]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_69),.I5(N_77),.LO(s_fracta_28_o[12:12]));
defparam desc181.INIT=64'hAA0FAA0CAA03AA00;
  LUT6_L desc182(.I0(s_opa_i[20:20]),.I1(s_exp_diff[2:2]),.I2(s_exp_diff[3:3]),.I3(N_987),.I4(s_expa_lt_expb),.I5(N_52),.LO(N_2229_i));
defparam desc182.INIT=64'hAAAA0003AAAA0000;
  LUT5_L desc183(.I0(s_opa_i[19:19]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_989),.LO(N_2225_i));
defparam desc183.INIT=32'hAA03AA00;
  LUT5_L desc184(.I0(s_opa_i[17:17]),.I1(s_exp_diff[3:3]),.I2(N_987),.I3(s_expa_lt_expb),.I4(N_77),.LO(N_2223_i));
defparam desc184.INIT=32'hAA03AA00;
  LUT6 un5_s_sticky_1_df0_lut6_2_RNO_0(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[1:1]),.I4(s_opb_i[0:0]),.I5(N_2199_1),.O(v_count_56_1[1:1]));
defparam un5_s_sticky_1_df0_lut6_2_RNO_0.INIT=64'hFFFF0055FFFF0054;
  LUT6_L desc185(.I0(s_opa_i[2:2]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_106),.I5(N_2119),.LO(s_fracta_28_o_i_m4[5:5]));
defparam desc185.INIT=64'hAA0FAA03AA0CAA00;
  LUT6_L desc186(.I0(s_opa_i[0:0]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_88),.I5(N_104),.LO(s_fracta_28_o[3:3]));
defparam desc186.INIT=64'hAA0FAA0CAA03AA00;
  LUT5 m47(.I0(s_opa_i[0:0]),.I1(v_count[1:1]),.I2(v_count[2:2]),.I3(N_1617),.I4(v_count_i),.O(N_48_0));
defparam m47.INIT=32'h0B080300;
  LUT6_L desc187(.I0(s_opb_i[0:0]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_88),.I5(N_104),.LO(s_fractb_28_o[3:3]));
defparam desc187.INIT=64'h0FAA0CAA03AA00AA;
  LUT4_L desc188(.I0(s_opa_i[12:12]),.I1(N_987),.I2(s_expa_lt_expb),.I3(N_2240),.LO(N_1231_i));
defparam desc188.INIT=16'hA3A0;
  LUT4 m19(.I0(v_count[1:1]),.I1(v_count[2:2]),.I2(N_2103),.I3(N_1236),.O(N_1238));
defparam m19.INIT=16'h4073;
  LUT5 m26(.I0(v_count[1:1]),.I1(v_count[2:2]),.I2(N_1239),.I3(N_1277),.I4(N_26_0),.O(N_27_0));
defparam m26.INIT=32'hFEDC3210;
  LUT6 m45(.I0(s_opa_i[1:1]),.I1(s_opa_i[0:0]),.I2(v_count[1:1]),.I3(v_count[3:3]),.I4(v_count[2:2]),.I5(v_count[0:0]),.O(N_1245));
defparam m45.INIT=64'h0000000C0000000A;
  LUT5 m78(.I0(v_count[1:1]),.I1(v_count[2:2]),.I2(N_1239),.I3(N_1277),.I4(N_33_0),.O(N_1267));
defparam m78.INIT=32'hFB73C840;
  LUT6_L desc189(.I0(s_opb_i[2:2]),.I1(s_exp_diff[4:4]),.I2(OVER),.I3(s_expa_lt_expb),.I4(N_106),.I5(N_2119),.LO(N_2122_i));
defparam desc189.INIT=64'h0FAA03AA0CAA00AA;
  LUT6 m58(.I0(v_count[1:1]),.I1(v_count[3:3]),.I2(v_count[2:2]),.I3(N_2103),.I4(N_26_0),.I5(N_1236),.O(pre_norm_div_dvdnd_0));
defparam m58.INIT=64'h0400070334303733;
  LUT5_L m69(.I0(v_count[3:3]),.I1(v_count[2:2]),.I2(N_1240),.I3(N_26_0),.I4(N_1238),.LO(pre_norm_div_dvdnd_4));
defparam m69.INIT=32'hABEF0145;
  LUT6_L m93_e(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[12:12]),.I4(s_opb_i[16:16]),.I5(N_129_mux),.LO(N_1292));
defparam m93_e.INIT=64'h0000F2F20000F2F3;
  LUT5 m80(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(N_1245),.I3(N_1267),.I4(N_1249),.O(pre_norm_div_dvdnd_8));
defparam m80.INIT=32'hC0D1E2F3;
  LUT6 m96(.I0(s_opb_i[21:21]),.I1(s_opb_i[17:17]),.I2(s_opb_i[19:19]),.I3(N_1294),.I4(N_1084_i),.I5(N_1292),.O(N_143_mux));
defparam m96.INIT=64'h0055000001550000;
  LUT3 un1_opa_i_3_5_cry_1_RNO(.I0(s_opb_i[24:24]),.I1(s_opa_i[24:24]),.I2(s_expa_lt_expb),.O(N_1108_i));
defparam un1_opa_i_3_5_cry_1_RNO.INIT=8'h53;
  LUT3 un1_opa_i_3_5_cry_2_RNO(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(s_expa_lt_expb),.O(N_1109_i));
defparam un1_opa_i_3_5_cry_2_RNO.INIT=8'h53;
  LUT3 un1_opa_i_3_5_cry_3_RNO(.I0(s_opa_i[26:26]),.I1(s_opb_i[26:26]),.I2(s_expa_lt_expb),.O(N_1110_i));
defparam un1_opa_i_3_5_cry_3_RNO.INIT=8'h35;
  LUT3 un1_opa_i_3_5_cry_4_RNO(.I0(s_opa_i[27:27]),.I1(s_opb_i[27:27]),.I2(s_expa_lt_expb),.O(N_1111_i));
defparam un1_opa_i_3_5_cry_4_RNO.INIT=8'h35;
  LUT3 un1_opa_i_3_5_cry_5_RNO(.I0(s_opa_i[28:28]),.I1(s_opb_i[28:28]),.I2(s_expa_lt_expb),.O(N_1112_i));
defparam un1_opa_i_3_5_cry_5_RNO.INIT=8'h35;
  LUT3 un1_opa_i_3_5_cry_6_RNO(.I0(s_opa_i[29:29]),.I1(s_opb_i[29:29]),.I2(s_expa_lt_expb),.O(N_1113_i));
defparam un1_opa_i_3_5_cry_6_RNO.INIT=8'h35;
  LUT5 un1_opa_i_3_4_cry_0_RNO_0(.I0(s_opb_i[23:23]),.I1(s_opa_i[23:23]),.I2(N_243),.I3(N_244),.I4(s_mux_diff),.O(un1_opa_i_3_4[0:0]));
defparam un1_opa_i_3_4_cry_0_RNO_0.INIT=32'hEAC0153F;
  LUT5 desc190(.I0(s_opb_i[29:29]),.I1(N_1138),.I2(N_227),.I3(N_244),.I4(N_1137),.O(un1_opa_i_3_4_axb_6));
defparam desc190.INIT=32'h050F363C;
  LUT5 desc191(.I0(un1_opa_i_i_m3_lut6_2_O6[7:7]),.I1(N_1140),.I2(N_1139),.I3(un1_opa_i_2_i[7:7]),.I4(s_mux_diff),.O(un1_opa_i_3_axb_0));
defparam desc191.INIT=32'hA95656A9;
  FDR desc192(.Q(prenorm_addsub_fractb_28_o[0:0]),.D(un3_s_fracta_28_o),.C(clk_i),.R(s_expa_lt_expb_i));
  FDR desc193(.Q(prenorm_addsub_fractb_28_o[1:1]),.D(s_fract_shr_28[1:1]),.C(clk_i),.R(s_expa_lt_expb_i));
  FDR desc194(.Q(prenorm_addsub_fractb_28_o[2:2]),.D(fractb_28_oc),.C(clk_i),.R(s_expa_lt_expb_i));
  FDS desc195(.Q(prenorm_addsub_fracta_28_o[26:26]),.D(N_60_mux),.C(clk_i),.S(s_expa_lt_expb));
  FDR desc196(.Q(prenorm_addsub_fracta_28_o[0:0]),.D(un3_s_fracta_28_o),.C(clk_i),.R(s_expa_lt_expb));
  FDR desc197(.Q(prenorm_addsub_fracta_28_o[1:1]),.D(s_fract_shr_28[1:1]),.C(clk_i),.R(s_expa_lt_expb));
  FDR desc198(.Q(prenorm_addsub_fracta_28_o[2:2]),.D(fractb_28_oc),.C(clk_i),.R(s_expa_lt_expb));
  XORCY un1_opa_i_3_s_7_cZ(.LI(un1_opa_i_3_axb_7),.CI(un1_opa_i_3_cry_6),.O(un1_opa_i_3_s_7));
  XORCY un1_opa_i_3_s_6_cZ(.LI(un1_opa_i_3_axb_6),.CI(un1_opa_i_3_cry_5),.O(un1_opa_i_3_s_6));
  MUXCY_L un1_opa_i_3_cry_6_cZ(.DI(un1_opa_i_3_4[6:6]),.CI(un1_opa_i_3_cry_5),.S(un1_opa_i_3_axb_6),.LO(un1_opa_i_3_cry_6));
  XORCY un1_opa_i_3_s_5_cZ(.LI(un1_opa_i_3_axb_5),.CI(un1_opa_i_3_cry_4),.O(un1_opa_i_3_s_5));
  MUXCY_L un1_opa_i_3_cry_5_cZ(.DI(un1_opa_i_3_4[5:5]),.CI(un1_opa_i_3_cry_4),.S(un1_opa_i_3_axb_5),.LO(un1_opa_i_3_cry_5));
  XORCY un1_opa_i_3_s_4_cZ(.LI(un1_opa_i_3_axb_4),.CI(un1_opa_i_3_cry_3),.O(un1_opa_i_3_s_4));
  MUXCY_L un1_opa_i_3_cry_4_cZ(.DI(un1_opa_i_3_4[4:4]),.CI(un1_opa_i_3_cry_3),.S(un1_opa_i_3_axb_4),.LO(un1_opa_i_3_cry_4));
  XORCY un1_opa_i_3_s_3_cZ(.LI(un1_opa_i_3_axb_3),.CI(un1_opa_i_3_cry_2),.O(un1_opa_i_3_s_3));
  MUXCY_L un1_opa_i_3_cry_3_cZ(.DI(un1_opa_i_3_4[3:3]),.CI(un1_opa_i_3_cry_2),.S(un1_opa_i_3_axb_3),.LO(un1_opa_i_3_cry_3));
  XORCY un1_opa_i_3_s_2_cZ(.LI(un1_opa_i_3_axb_2),.CI(un1_opa_i_3_cry_1),.O(un1_opa_i_3_s_2));
  MUXCY_L un1_opa_i_3_cry_2_cZ(.DI(un1_opa_i_3_4[2:2]),.CI(un1_opa_i_3_cry_1),.S(un1_opa_i_3_axb_2),.LO(un1_opa_i_3_cry_2));
  XORCY un1_opa_i_3_s_1_cZ(.LI(un1_opa_i_3_axb_1),.CI(un1_opa_i_3_cry_0),.O(un1_opa_i_3_s_1));
  MUXCY_L un1_opa_i_3_cry_1_cZ(.DI(un1_opa_i_3_4[1:1]),.CI(un1_opa_i_3_cry_0),.S(un1_opa_i_3_axb_1),.LO(un1_opa_i_3_cry_1));
  MUXCY_L un1_opa_i_3_cry_0_cZ(.DI(un1_opa_i_3_5[0:0]),.CI(GND),.S(un1_opa_i_3_axb_0),.LO(un1_opa_i_3_cry_0));
  XORCY un1_opa_i_3_4_s_7(.LI(un1_opa_i_3_4_axb_7),.CI(un1_opa_i_3_4_cry_6),.O(un1_opa_i_3_4[7:7]));
  XORCY un1_opa_i_3_4_s_6(.LI(un1_opa_i_3_4_axb_6),.CI(un1_opa_i_3_4_cry_5),.O(un1_opa_i_3_4[6:6]));
  MUXCY_L un1_opa_i_3_4_cry_6_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_5),.S(un1_opa_i_3_4_axb_6),.LO(un1_opa_i_3_4_cry_6));
  XORCY un1_opa_i_3_4_s_5(.LI(un1_opa_i_3_4_axb_5),.CI(un1_opa_i_3_4_cry_4),.O(un1_opa_i_3_4[5:5]));
  MUXCY_L un1_opa_i_3_4_cry_5_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_4),.S(un1_opa_i_3_4_axb_5),.LO(un1_opa_i_3_4_cry_5));
  XORCY un1_opa_i_3_4_s_4(.LI(un1_opa_i_3_4_axb_4),.CI(un1_opa_i_3_4_cry_3),.O(un1_opa_i_3_4[4:4]));
  MUXCY_L un1_opa_i_3_4_cry_4_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_3),.S(un1_opa_i_3_4_axb_4),.LO(un1_opa_i_3_4_cry_4));
  XORCY un1_opa_i_3_4_s_3(.LI(un1_opa_i_3_4_axb_3),.CI(un1_opa_i_3_4_cry_2),.O(un1_opa_i_3_4[3:3]));
  MUXCY_L un1_opa_i_3_4_cry_3_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_2),.S(un1_opa_i_3_4_axb_3),.LO(un1_opa_i_3_4_cry_3));
  XORCY un1_opa_i_3_4_s_2(.LI(un1_opa_i_3_4_axb_2),.CI(un1_opa_i_3_4_cry_1),.O(un1_opa_i_3_4[2:2]));
  MUXCY_L un1_opa_i_3_4_cry_2_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_1),.S(un1_opa_i_3_4_axb_2),.LO(un1_opa_i_3_4_cry_2));
  XORCY un1_opa_i_3_4_s_1(.LI(un1_opa_i_3_4_axb_1),.CI(un1_opa_i_3_4_cry_0),.O(un1_opa_i_3_4[1:1]));
  MUXCY_L un1_opa_i_3_4_cry_1_cZ(.DI(s_mux_diff),.CI(un1_opa_i_3_4_cry_0),.S(un1_opa_i_3_4_axb_1),.LO(un1_opa_i_3_4_cry_1));
  MUXCY_L un1_opa_i_3_4_cry_0_cZ(.DI(un27[7:7]),.CI(GND),.S(un1_opa_i_3_4[0:0]),.LO(un1_opa_i_3_4_cry_0));
  XORCY un1_opa_i_3_5_s_7(.LI(un1_opa_i_3_5_axb_7),.CI(un1_opa_i_3_5_cry_6),.O(un1_opa_i_3_5[7:7]));
  XORCY un1_opa_i_3_5_s_6(.LI(un1_opa_i_3_5_axb_6),.CI(un1_opa_i_3_5_cry_5),.O(un1_opa_i_3_5[6:6]));
  MUXCY_L un1_opa_i_3_5_cry_6_cZ(.DI(N_1113_i),.CI(un1_opa_i_3_5_cry_5),.S(un1_opa_i_3_5_axb_6),.LO(un1_opa_i_3_5_cry_6));
  XORCY un1_opa_i_3_5_s_5(.LI(un1_opa_i_3_5_axb_5),.CI(un1_opa_i_3_5_cry_4),.O(un1_opa_i_3_5[5:5]));
  MUXCY_L un1_opa_i_3_5_cry_5_cZ(.DI(N_1112_i),.CI(un1_opa_i_3_5_cry_4),.S(un1_opa_i_3_5_axb_5),.LO(un1_opa_i_3_5_cry_5));
  XORCY un1_opa_i_3_5_s_4(.LI(un1_opa_i_3_5_axb_4),.CI(un1_opa_i_3_5_cry_3),.O(un1_opa_i_3_5[4:4]));
  MUXCY_L un1_opa_i_3_5_cry_4_cZ(.DI(N_1111_i),.CI(un1_opa_i_3_5_cry_3),.S(un1_opa_i_3_5_axb_4),.LO(un1_opa_i_3_5_cry_4));
  XORCY un1_opa_i_3_5_s_3(.LI(un1_opa_i_3_5_axb_3),.CI(un1_opa_i_3_5_cry_2),.O(un1_opa_i_3_5[3:3]));
  MUXCY_L un1_opa_i_3_5_cry_3_cZ(.DI(N_1110_i),.CI(un1_opa_i_3_5_cry_2),.S(un1_opa_i_3_5_axb_3),.LO(un1_opa_i_3_5_cry_3));
  XORCY un1_opa_i_3_5_s_2(.LI(un1_opa_i_3_5_axb_2),.CI(un1_opa_i_3_5_cry_1),.O(un1_opa_i_3_5[2:2]));
  MUXCY_L un1_opa_i_3_5_cry_2_cZ(.DI(N_1109_i),.CI(un1_opa_i_3_5_cry_1),.S(un1_opa_i_3_5_axb_2),.LO(un1_opa_i_3_5_cry_2));
  XORCY un1_opa_i_3_5_s_1(.LI(un1_opa_i_3_5_axb_1),.CI(un1_opa_i_3_5_cry_0),.O(un1_opa_i_3_5[1:1]));
  MUXCY_L un1_opa_i_3_5_cry_1_cZ(.DI(N_1108_i),.CI(un1_opa_i_3_5_cry_0),.S(un1_opa_i_3_5_axb_1),.LO(un1_opa_i_3_5_cry_1));
  MUXCY_L un1_opa_i_3_5_cry_0_cZ(.DI(N_1107_i),.CI(GND),.S(un1_opa_i_3_5[0:0]),.LO(un1_opa_i_3_5_cry_0));
  MUXCY_L desc199(.DI(s_expa_lt_expb_lt4),.CI(s_expa_lt_expb_cry[2:2]),.S(s_expa_lt_expb_df4),.LO(s_expa_lt_expb_cry[4:4]));
  MUXCY_L desc200(.DI(s_expa_lt_expb_lt2),.CI(s_expa_lt_expb_cry[0:0]),.S(s_expa_lt_expb_df2),.LO(s_expa_lt_expb_cry[2:2]));
  MUXCY_L desc201(.DI(s_expa_lt_expb_lt0),.CI(GND),.S(s_expa_lt_expb_df0),.LO(s_expa_lt_expb_cry[0:0]));
  MUXCY_L desc202(.DI(un5_s_sticky_1_lt4),.CI(un5_s_sticky_1_cry[2:2]),.S(un5_s_sticky_1_df4),.LO(un5_s_sticky_1_cry[4:4]));
  MUXCY_L desc203(.DI(un5_s_sticky_1_lt2),.CI(un5_s_sticky_1_cry[0:0]),.S(un5_s_sticky_1_df2),.LO(un5_s_sticky_1_cry[2:2]));
  MUXCY_L desc204(.DI(un5_s_sticky_1_lt0),.CI(GND),.S(un5_s_sticky_1_df0),.LO(un5_s_sticky_1_cry[0:0]));
  MUXCY_L desc205(.DI(un5_s_sticky_0_lt4),.CI(un5_s_sticky_0_cry[2:2]),.S(un5_s_sticky_0_df4),.LO(un5_s_sticky_0_cry[4:4]));
  MUXCY_L desc206(.DI(un5_s_sticky_0_lt2),.CI(un5_s_sticky_0_cry[0:0]),.S(un5_s_sticky_0_df2),.LO(un5_s_sticky_0_cry[2:2]));
  MUXCY_L desc207(.DI(un5_s_sticky_0_lt0),.CI(GND),.S(un5_s_sticky_0_df0),.LO(un5_s_sticky_0_cry[0:0]));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT4 desc208(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_exp_diff[4:4]),.O(N_1053));
defparam desc208.INIT=16'h0100;
  LUT5 desc209(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_exp_diff[4:4]),.I4(N_2234),.O(N_60_mux));
defparam desc209.INIT=32'h00010000;
  LUT4 desc210(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_expa_lt_expb),.I3(N_1084_i),.O(N_1057));
defparam desc210.INIT=16'hF101;
  LUT3 desc211(.I0(s_opa_i[24:24]),.I1(s_opa_i[23:23]),.I2(N_1077),.O(N_378_i));
defparam desc211.INIT=8'hC9;
  LUT3 desc212(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_expa_lt_expb),.O(N_244));
defparam desc212.INIT=8'h01;
  LUT3 desc213(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_exp_10_o_0),.O(s_exp_10_o));
defparam desc213.INIT=8'hE1;
  LUT2 desc214(.I0(s_opb_i[3:3]),.I1(s_opb_i[1:1]),.O(N_757));
defparam desc214.INIT=4'h1;
  LUT4 desc215(.I0(s_opb_i[11:11]),.I1(s_opb_i[3:3]),.I2(s_opb_i[1:1]),.I3(s_opb_i[7:7]),.O(N_761));
defparam desc215.INIT=16'h0001;
  LUT2 desc216(.I0(s_opa_i[3:3]),.I1(s_opa_i[4:4]),.O(N_1604));
defparam desc216.INIT=4'hE;
  LUT4 desc217(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[4:4]),.I3(s_opa_i[1:1]),.O(N_254));
defparam desc217.INIT=16'h0001;
  LUT2 desc218(.I0(s_opa_i[12:12]),.I1(s_opa_i[11:11]),.O(N_1596));
defparam desc218.INIT=4'hE;
  LUT5 desc219(.I0(s_opa_i[12:12]),.I1(s_opa_i[11:11]),.I2(s_opa_i[10:10]),.I3(s_opa_i[9:9]),.I4(N_254),.O(N_267));
defparam desc219.INIT=32'h00010000;
  LUT3 desc220(.I0(s_opb_i[23:23]),.I1(s_opa_i[23:23]),.I2(s_expa_lt_expb),.O(un1_opa_i_i_m3_lut6_2_O6[7:7]));
defparam desc220.INIT=8'hAC;
  LUT2 desc221(.I0(N_1083),.I1(s_opb_i[23:23]),.O(un4_s_expb_in_2_i_0_e));
defparam desc221.INIT=4'hD;
  LUT3 desc222(.I0(s_opb_i[23:23]),.I1(s_opa_i[23:23]),.I2(s_expa_lt_expb),.O(un27_0_i_m3_lut6_2_O6[7:7]));
defparam desc222.INIT=8'hCA;
  LUT3 desc223(.I0(s_opb_i[24:24]),.I1(s_opa_i[24:24]),.I2(s_expa_lt_expb),.O(un27_0_i_m3_lut6_2_O5[7:7]));
defparam desc223.INIT=8'hCA;
  LUT3 desc224(.I0(s_opa_i[28:28]),.I1(s_opb_i[28:28]),.I2(s_expa_lt_expb),.O(N_163));
defparam desc224.INIT=8'hAC;
  LUT3 desc225(.I0(s_opa_i[29:29]),.I1(s_opb_i[29:29]),.I2(s_expa_lt_expb),.O(N_164));
defparam desc225.INIT=8'hAC;
  LUT3 desc226(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(s_expa_lt_expb),.O(un27_0_i_m3_lut6_2_O6[5:5]));
defparam desc226.INIT=8'hCA;
  LUT3 desc227(.I0(s_opa_i[26:26]),.I1(s_opb_i[26:26]),.I2(s_expa_lt_expb),.O(un27_0_i_m3_lut6_2_O5[5:5]));
defparam desc227.INIT=8'hAC;
  LUT3 desc228(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.O(OVER));
defparam desc228.INIT=8'hFE;
  LUT4 desc229(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[6:6]),.I2(s_exp_diff[7:7]),.I3(s_exp_diff[4:4]),.O(N_987));
defparam desc229.INIT=16'hFFFE;
  LUT4 desc230(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[16:16]),.O(N_2197));
defparam desc230.INIT=16'h0001;
  LUT4 desc231(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[12:12]),.O(N_1050));
defparam desc231.INIT=16'h0001;
  LUT3 desc232(.I0(s_opa_i[29:29]),.I1(s_expa_lt_expb),.I2(N_1084_i),.O(N_227));
defparam desc232.INIT=8'h80;
  LUT3 desc233(.I0(s_opb_i[12:12]),.I1(s_opa_i[12:12]),.I2(s_expa_lt_expb),.O(N_1230));
defparam desc233.INIT=8'h53;
  LUT3 m96_e_lut6_2_o6(.I0(s_opb_i[19:19]),.I1(s_opb_i[20:20]),.I2(s_opb_i[18:18]),.O(N_1294));
defparam m96_e_lut6_2_o6.INIT=8'h23;
  LUT5 m96_e_lut6_2_o5(.I0(s_opb_i[17:17]),.I1(s_opb_i[19:19]),.I2(s_opb_i[20:20]),.I3(s_opb_i[18:18]),.I4(N_2197),.O(N_2242));
defparam m96_e_lut6_2_o5.INIT=32'hFFFE0000;
  LUT3 m123_e_lut6_2_o6(.I0(s_opb_i[2:2]),.I1(s_opb_i[1:1]),.I2(s_opb_i[0:0]),.O(N_1286));
defparam m123_e_lut6_2_o6.INIT=8'h10;
  LUT4 m123_e_lut6_2_o5(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[1:1]),.I3(s_opb_i[0:0]),.O(N_1051));
defparam m123_e_lut6_2_o5.INIT=16'h0001;
  LUT4 desc234(.I0(s_opa_i[8:8]),.I1(s_opa_i[10:10]),.I2(s_opa_i[11:11]),.I3(s_opa_i[9:9]),.O(un2_s_snan_o_20));
defparam desc234.INIT=16'h0001;
  LUT2 desc235(.I0(s_opa_i[9:9]),.I1(s_opa_i[5:5]),.O(N_255));
defparam desc235.INIT=4'h1;
  LUT5 un3_s_fracta_28_o_0_o4_3_0_lut6_2_o6(.I0(s_opb_i[14:14]),.I1(s_opb_i[15:15]),.I2(s_opa_i[14:14]),.I3(s_opa_i[15:15]),.I4(s_expa_lt_expb),.O(un3_s_fracta_28_o_0_o4_3_0));
defparam un3_s_fracta_28_o_0_o4_3_0_lut6_2_o6.INIT=32'hEEEEFFF0;
  LUT2 un3_s_fracta_28_o_0_o4_3_0_lut6_2_o5(.I0(s_opa_i[14:14]),.I1(s_opa_i[15:15]),.O(N_1159));
defparam un3_s_fracta_28_o_0_o4_3_0_lut6_2_o5.INIT=4'hE;
  LUT4 desc236(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[1:1]),.O(v_count_56_1_0_2));
defparam desc236.INIT=16'h00BA;
  LUT5 desc237(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[1:1]),.I4(s_opb_i[0:0]),.O(N_2254));
defparam desc237.INIT=32'h00000001;
  LUT5 desc238(.I0(s_opb_i[21:21]),.I1(s_opb_i[19:19]),.I2(s_opb_i[20:20]),.I3(s_opb_i[18:18]),.I4(s_opb_i[22:22]),.O(N_138));
defparam desc238.INIT=32'hFF31FF30;
  LUT2 desc239(.I0(s_opb_i[19:19]),.I1(s_opb_i[20:20]),.O(N_2180));
defparam desc239.INIT=4'hE;
  LUT3 desc240(.I0(s_exp_diff[1:1]),.I1(N_7),.I2(N_9),.O(N_35));
defparam desc240.INIT=8'hE4;
  LUT3 desc241(.I0(s_exp_diff[1:1]),.I1(N_4),.I2(N_6),.O(N_32));
defparam desc241.INIT=8'hE4;
  LUT3 desc242(.I0(s_exp_diff[1:1]),.I1(N_21),.I2(N_19),.O(N_47));
defparam desc242.INIT=8'hD8;
  LUT3 desc243(.I0(s_exp_diff[1:1]),.I1(N_8),.I2(N_10),.O(N_36));
defparam desc243.INIT=8'hE4;
  LUT3 desc244(.I0(s_exp_diff[1:1]),.I1(N_21),.I2(N_23),.O(N_49));
defparam desc244.INIT=8'hE4;
  LUT3 desc245(.I0(s_exp_diff[1:1]),.I1(N_15),.I2(N_17_0),.O(N_43_0));
defparam desc245.INIT=8'hE4;
  LUT4 desc246(.I0(s_opb_i[23:23]),.I1(s_opa_i[24:24]),.I2(N_1077),.I3(N_1083),.O(N_1137));
defparam desc246.INIT=16'h0312;
  LUT2 desc247(.I0(s_opb_i[30:30]),.I1(s_opb_i[23:23]),.O(N_168_2));
defparam desc247.INIT=4'h8;
  LUT3 desc248(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[1:1]),.I2(N_26),.O(N_995));
defparam desc248.INIT=8'hEF;
  LUT3 desc249(.I0(s_exp_diff[1:1]),.I1(N_11),.I2(N_13),.O(N_39));
defparam desc249.INIT=8'hE4;
  LUT5 desc250(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_45),.I3(N_49),.I4(N_53_0),.O(N_17));
defparam desc250.INIT=32'h89ABCDEF;
  LUT2 desc251(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.O(N_1043));
defparam desc251.INIT=4'h1;
  LUT4 desc252(.I0(s_exp_diff[4:4]),.I1(s_exp_diff[3:3]),.I2(N_70_0),.I3(N_78),.O(OUT13_1));
defparam desc252.INIT=16'h5410;
  LUT3 desc253(.I0(s_exp_diff[3:3]),.I1(N_2118),.I2(N_70_0),.O(N_2119));
defparam desc253.INIT=8'hE4;
  LUT2 desc254(.I0(s_opa_i[3:3]),.I1(s_opa_i[1:1]),.O(N_1217));
defparam desc254.INIT=4'h1;
  LUT3 desc255(.I0(s_opa_i[1:1]),.I1(s_expa_lt_expb),.I2(N_2107),.O(s_fractb_28_o_i_o4_RNIN0MT_O5[4:4]));
defparam desc255.INIT=8'h8B;
  LUT3 m36_lut6_2_o6(.I0(v_count[2:2]),.I1(N_1624),.I2(N_1628),.O(N_1242));
defparam m36_lut6_2_o6.INIT=8'h27;
  LUT5 m36_lut6_2_o5(.I0(v_count[3:3]),.I1(v_count[2:2]),.I2(N_1624),.I3(N_1628),.I4(N_53),.O(N_1257_i));
defparam m36_lut6_2_o5.INIT=32'hFBEA5140;
  LUT3 m57_lut6_2_o6(.I0(v_count[2:2]),.I1(N_26_0),.I2(N_1236),.O(N_1249));
defparam m57_lut6_2_o6.INIT=8'hE4;
  LUT3 m57_lut6_2_o5(.I0(v_count[2:2]),.I1(N_46),.I2(N_33_0),.O(N_70));
defparam m57_lut6_2_o5.INIT=8'h4E;
  LUT3 m75_lut6_2_o6(.I0(v_count[2:2]),.I1(N_41),.I2(N_1628),.O(N_1264));
defparam m75_lut6_2_o6.INIT=8'h1B;
  LUT3 m75_lut6_2_o5(.I0(v_count[2:2]),.I1(N_43),.I2(N_1630),.O(N_67));
defparam m75_lut6_2_o5.INIT=8'hE4;
  LUT3 desc256(.I0(s_opa_i[23:23]),.I1(s_expa_lt_expb),.I2(N_1084_i),.O(N_1139));
defparam desc256.INIT=8'h80;
  LUT3 desc257(.I0(s_opb_i[1:1]),.I1(s_expa_lt_expb),.I2(N_2107),.O(N_2129_i));
defparam desc257.INIT=8'h2E;
  LUT2 desc258(.I0(s_opa_i[0:0]),.I1(s_opa_i[23:23]),.O(pre_norm_sqrt_fracta_o_0));
defparam desc258.INIT=4'h8;
  LUT3 desc259(.I0(s_opa_i[23:23]),.I1(pre_norm_div_dvdnd_8),.I2(pre_norm_div_dvdnd_9),.O(pre_norm_sqrt_fracta_o_18));
defparam desc259.INIT=8'hE4;
  LUT4 s_expa_lt_expb_df6_lut6_2_o6(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(s_opa_i[29:29]),.I3(s_opb_i[29:29]),.O(s_expa_lt_expb_df6));
defparam s_expa_lt_expb_df6_lut6_2_o6.INIT=16'h9009;
  LUT4 s_expa_lt_expb_df6_lut6_2_o5(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(s_opa_i[29:29]),.I3(s_opb_i[29:29]),.O(s_expa_lt_expb_lt6));
defparam s_expa_lt_expb_df6_lut6_2_o5.INIT=16'h44D4;
  LUT4 s_expa_lt_expb_df4_lut6_2_o6(.I0(s_opa_i[28:28]),.I1(s_opa_i[27:27]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.O(s_expa_lt_expb_df4));
defparam s_expa_lt_expb_df4_lut6_2_o6.INIT=16'h8421;
  LUT4 s_expa_lt_expb_df4_lut6_2_o5(.I0(s_opa_i[28:28]),.I1(s_opa_i[27:27]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.O(s_expa_lt_expb_lt4));
defparam s_expa_lt_expb_df4_lut6_2_o5.INIT=16'h0A8E;
  LUT4 s_expa_lt_expb_df2_lut6_2_o6(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(s_opa_i[26:26]),.I3(s_opb_i[26:26]),.O(s_expa_lt_expb_df2));
defparam s_expa_lt_expb_df2_lut6_2_o6.INIT=16'h9009;
  LUT4 s_expa_lt_expb_df2_lut6_2_o5(.I0(s_opb_i[25:25]),.I1(s_opa_i[25:25]),.I2(s_opa_i[26:26]),.I3(s_opb_i[26:26]),.O(s_expa_lt_expb_lt2));
defparam s_expa_lt_expb_df2_lut6_2_o5.INIT=16'h40F4;
  LUT4 s_expa_lt_expb_df0_lut6_2_o6(.I0(s_opb_i[24:24]),.I1(s_opb_i[23:23]),.I2(s_opa_i[24:24]),.I3(s_opa_i[23:23]),.O(s_expa_lt_expb_df0));
defparam s_expa_lt_expb_df0_lut6_2_o6.INIT=16'h8421;
  LUT4 s_expa_lt_expb_df0_lut6_2_o5(.I0(s_opb_i[24:24]),.I1(s_opb_i[23:23]),.I2(s_opa_i[24:24]),.I3(s_opa_i[23:23]),.O(s_expa_lt_expb_lt0));
defparam s_expa_lt_expb_df0_lut6_2_o5.INIT=16'h7150;
  LUT2 un5_s_sticky_1_df6_lut6_2_o6(.I0(s_exp_diff[6:6]),.I1(s_exp_diff[7:7]),.O(un5_s_sticky_1_df6));
defparam un5_s_sticky_1_df6_lut6_2_o6.INIT=4'h1;
  LUT2 un5_s_sticky_1_df6_lut6_2_o5(.I0(s_exp_diff[6:6]),.I1(s_exp_diff[7:7]),.O(un5_s_sticky_1_lt6));
defparam un5_s_sticky_1_df6_lut6_2_o5.INIT=4'hE;
  LUT3 un5_s_sticky_1_df4_lut6_2_o6(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[4:4]),.I2(v_count_56_1[4:4]),.O(un5_s_sticky_1_df4));
defparam un5_s_sticky_1_df4_lut6_2_o6.INIT=8'h41;
  LUT3 un5_s_sticky_1_df4_lut6_2_o5(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[4:4]),.I2(v_count_56_1[4:4]),.O(un5_s_sticky_1_lt4));
defparam un5_s_sticky_1_df4_lut6_2_o5.INIT=8'hAE;
  LUT4 un5_s_sticky_1_df2_lut6_2_o6(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_64_mux),.I3(v_count_56_1[3:3]),.O(un5_s_sticky_1_df2));
defparam un5_s_sticky_1_df2_lut6_2_o6.INIT=16'h8421;
  LUT4 un5_s_sticky_1_df2_lut6_2_o5(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(N_64_mux),.I3(v_count_56_1[3:3]),.O(un5_s_sticky_1_lt2));
defparam un5_s_sticky_1_df2_lut6_2_o5.INIT=16'h08CE;
  LUT4 un5_s_sticky_1_df0_lut6_2_o6(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(v_count_56_1[0:0]),.I3(v_count_56_1[1:1]),.O(un5_s_sticky_1_df0));
defparam un5_s_sticky_1_df0_lut6_2_o6.INIT=16'h8421;
  LUT4 un5_s_sticky_1_df0_lut6_2_o5(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(v_count_56_1[0:0]),.I3(v_count_56_1[1:1]),.O(un5_s_sticky_1_lt0));
defparam un5_s_sticky_1_df0_lut6_2_o5.INIT=16'h08CE;
  LUT2 un5_s_sticky_0_df6_lut6_2_o6(.I0(s_exp_diff[6:6]),.I1(s_exp_diff[7:7]),.O(un5_s_sticky_0_df6));
defparam un5_s_sticky_0_df6_lut6_2_o6.INIT=4'h1;
  LUT2 un5_s_sticky_0_df6_lut6_2_o5(.I0(s_exp_diff[6:6]),.I1(s_exp_diff[7:7]),.O(un5_s_sticky_0_lt6));
defparam un5_s_sticky_0_df6_lut6_2_o5.INIT=4'hE;
  LUT3 un5_s_sticky_0_df4_lut6_2_o6(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[4:4]),.I2(v_count_56_0[4:4]),.O(un5_s_sticky_0_df4));
defparam un5_s_sticky_0_df4_lut6_2_o6.INIT=8'h41;
  LUT3 un5_s_sticky_0_df4_lut6_2_o5(.I0(s_exp_diff[5:5]),.I1(s_exp_diff[4:4]),.I2(v_count_56_0[4:4]),.O(un5_s_sticky_0_lt4));
defparam un5_s_sticky_0_df4_lut6_2_o5.INIT=8'hAE;
  LUT4 un5_s_sticky_0_df2_lut6_2_o6(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(v_count_56_0[3:3]),.I3(N_194_i),.O(un5_s_sticky_0_df2));
defparam un5_s_sticky_0_df2_lut6_2_o6.INIT=16'h8241;
  LUT4 un5_s_sticky_0_df2_lut6_2_o5(.I0(s_exp_diff[2:2]),.I1(s_exp_diff[3:3]),.I2(v_count_56_0[3:3]),.I3(N_194_i),.O(un5_s_sticky_0_lt2));
defparam un5_s_sticky_0_df2_lut6_2_o5.INIT=16'h0C8E;
  LUT4 un5_s_sticky_0_df0_lut6_2_o6(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(v_count_56_0[0:0]),.I3(v_count_56_0[1:1]),.O(un5_s_sticky_0_df0));
defparam un5_s_sticky_0_df0_lut6_2_o6.INIT=16'h8421;
  LUT4 un5_s_sticky_0_df0_lut6_2_o5(.I0(s_exp_diff[0:0]),.I1(s_exp_diff[1:1]),.I2(v_count_56_0[0:0]),.I3(v_count_56_0[1:1]),.O(un5_s_sticky_0_lt0));
defparam un5_s_sticky_0_df0_lut6_2_o5.INIT=16'h08CE;
endmodule
module addsub_28_inj (prenorm_addsub_fracta_28_o,prenorm_addsub_fractb_28_o,s_fpu_op_i,addsub_fract_o,s_opb_i_26,s_opb_i_1,s_opb_i_0,s_opb_i_2,s_opa_i_27,s_opa_i_0,s_opa_i_1,N_1941,N_1942_i,clk_i,result_2_2,N_1055,un1_s_infb,N_1979,addsub_sign_o,un2_s_snan_o_8,N_1166,un4_s_infa,result_3_0_0_i,N_36_0,result_2,N_1948);
input [26:0] prenorm_addsub_fracta_28_o ;
input [26:0] prenorm_addsub_fractb_28_o ;
input s_fpu_op_i ;
output [27:0] addsub_fract_o ;
input s_opb_i_26 ;
input s_opb_i_1 ;
input s_opb_i_0 ;
input s_opb_i_2 ;
input s_opa_i_27 ;
input s_opa_i_0 ;
input s_opa_i_1 ;
output N_1941 ;
output N_1942_i ;
input clk_i ;
input result_2_2 ;
input N_1055 ;
input un1_s_infb ;
output N_1979 ;
output addsub_sign_o ;
input un2_s_snan_o_8 ;
input N_1166 ;
input un4_s_infa ;
input result_3_0_0_i ;
output N_36_0 ;
input result_2 ;
output N_1948 ;
wire s_opb_i_26 ;
wire s_opb_i_1 ;
wire s_opb_i_0 ;
wire s_opb_i_2 ;
wire s_opa_i_27 ;
wire s_opa_i_0 ;
wire s_opa_i_1 ;
wire N_1941 ;
wire N_1942_i ;
wire clk_i ;
wire result_2_2 ;
wire N_1055 ;
wire un1_s_infb ;
wire N_1979 ;
wire addsub_sign_o ;
wire un2_s_snan_o_8 ;
wire N_1166 ;
wire un4_s_infa ;
wire result_3_0_0_i ;
wire N_36_0 ;
wire result_2 ;
wire N_1948 ;
wire [27:0] un1_fracta_i_10 ;
wire [27:0] un1_fracta_i_11 ;
wire [24:0] fracta_lt_fractb_cry ;
wire GND ;
wire VCC ;
wire fracta_lt_fractb_df0 ;
wire fracta_lt_fractb_lt0 ;
wire fracta_lt_fractb_df2 ;
wire fracta_lt_fractb_lt2 ;
wire fracta_lt_fractb_df4 ;
wire fracta_lt_fractb_lt4 ;
wire fracta_lt_fractb_df6 ;
wire fracta_lt_fractb_lt6 ;
wire fracta_lt_fractb_df8 ;
wire fracta_lt_fractb_lt8 ;
wire fracta_lt_fractb_df10 ;
wire fracta_lt_fractb_lt10 ;
wire fracta_lt_fractb_df12 ;
wire fracta_lt_fractb_lt12 ;
wire fracta_lt_fractb_df14 ;
wire fracta_lt_fractb_lt14 ;
wire fracta_lt_fractb_df16 ;
wire fracta_lt_fractb_lt16 ;
wire fracta_lt_fractb_df18 ;
wire fracta_lt_fractb_lt18 ;
wire fracta_lt_fractb_df20 ;
wire fracta_lt_fractb_lt20 ;
wire fracta_lt_fractb_df22 ;
wire fracta_lt_fractb_lt22 ;
wire fracta_lt_fractb_df24 ;
wire fracta_lt_fractb_lt24 ;
wire fracta_lt_fractb_df26 ;
wire fracta_lt_fractb_lt26 ;
wire fracta_lt_fractb ;
wire un1_fracta_i_s0_s_14_RNID77E1_O6 ;
wire N_2604_i ;
wire m33_2_1 ;
wire N_2605_i ;
wire N_2606_i ;
wire N_59_0_i ;
wire N_2607_i ;
wire N_2609_i ;
wire m33_3_1 ;
wire N_2610_i ;
wire N_2611_i ;
wire N_2613_i ;
wire N_2612_i ;
wire N_2614_i ;
wire m33_4_1 ;
wire N_2615_i ;
wire N_2616_i ;
wire N_2590_i ;
wire N_2617_i ;
wire N_2591_i ;
wire m33_0_1 ;
wire N_62_0_i ;
wire un1_fracta_i_s0_s_24_RNI55IC1_O6 ;
wire N_65_0_i ;
wire N_2595_i ;
wire N_2600_i ;
wire N_2596_i ;
wire N_2601_i ;
wire N_2597_i ;
wire N_2602_i ;
wire m33_1_1 ;
wire N_2598_i ;
wire N_2599_i ;
wire N_2603_i ;
wire un1_fracta_i_s0_cry_0_cy_RNO ;
wire un1_fracta_i_0_cry_0_cy_RNO ;
wire N_2608_i ;
wire un1_fracta_i_0_s_27_RNO ;
wire m33_1_4 ;
wire sign_o ;
wire un1_fracta_i_0_cry_0_cy ;
wire un1_fracta_i_s0_cry_0_cy ;
wire s_addop_1_1 ;
wire m33_3_3 ;
wire m33_2_3 ;
wire m33_1_3 ;
wire m33_0_3 ;
wire un1_fracta_i_s0_axb_26 ;
wire un1_fracta_i_s0_axb_25 ;
wire un1_fracta_i_s0_axb_24 ;
wire un1_fracta_i_s0_axb_23 ;
wire un1_fracta_i_s0_axb_22 ;
wire un1_fracta_i_s0_axb_21 ;
wire un1_fracta_i_s0_axb_20 ;
wire un1_fracta_i_s0_axb_19 ;
wire un1_fracta_i_s0_axb_18 ;
wire un1_fracta_i_s0_axb_17 ;
wire un1_fracta_i_s0_axb_16 ;
wire un1_fracta_i_s0_axb_15 ;
wire un1_fracta_i_s0_axb_14 ;
wire un1_fracta_i_s0_axb_13 ;
wire un1_fracta_i_s0_axb_12 ;
wire un1_fracta_i_s0_axb_11 ;
wire un1_fracta_i_s0_axb_10 ;
wire un1_fracta_i_s0_axb_9 ;
wire un1_fracta_i_s0_axb_8 ;
wire un1_fracta_i_s0_axb_7 ;
wire un1_fracta_i_s0_axb_6 ;
wire un1_fracta_i_s0_axb_5 ;
wire un1_fracta_i_s0_axb_4 ;
wire un1_fracta_i_s0_axb_3 ;
wire un1_fracta_i_s0_axb_2 ;
wire un1_fracta_i_s0_axb_1 ;
wire un1_fracta_i_s0_axb_0 ;
wire un1_fracta_i_0_axb_26 ;
wire un1_fracta_i_0_axb_25 ;
wire un1_fracta_i_0_axb_24 ;
wire un1_fracta_i_0_axb_23 ;
wire un1_fracta_i_0_axb_22 ;
wire un1_fracta_i_0_axb_21 ;
wire un1_fracta_i_0_axb_20 ;
wire un1_fracta_i_0_axb_19 ;
wire un1_fracta_i_0_axb_18 ;
wire un1_fracta_i_0_axb_17 ;
wire un1_fracta_i_0_axb_16 ;
wire un1_fracta_i_0_axb_15 ;
wire un1_fracta_i_0_axb_14 ;
wire un1_fracta_i_0_axb_13 ;
wire un1_fracta_i_0_axb_12 ;
wire un1_fracta_i_0_axb_11 ;
wire un1_fracta_i_0_axb_10 ;
wire un1_fracta_i_0_axb_9 ;
wire un1_fracta_i_0_axb_8 ;
wire un1_fracta_i_0_axb_7 ;
wire un1_fracta_i_0_axb_6 ;
wire un1_fracta_i_0_axb_5 ;
wire un1_fracta_i_0_axb_4 ;
wire un1_fracta_i_0_axb_3 ;
wire un1_fracta_i_0_axb_2 ;
wire un1_fracta_i_0_axb_1 ;
wire un1_fracta_i_0_axb_0 ;
wire m33_3 ;
wire m33_2 ;
wire m33_1 ;
wire m33_0 ;
wire un1_fracta_i_s0_cry_26 ;
wire un1_fracta_i_s0_cry_25 ;
wire un1_fracta_i_s0_cry_24 ;
wire un1_fracta_i_s0_cry_23 ;
wire un1_fracta_i_s0_cry_22 ;
wire un1_fracta_i_s0_cry_21 ;
wire un1_fracta_i_s0_cry_20 ;
wire un1_fracta_i_s0_cry_19 ;
wire un1_fracta_i_s0_cry_18 ;
wire un1_fracta_i_s0_cry_17 ;
wire un1_fracta_i_s0_cry_16 ;
wire un1_fracta_i_s0_cry_15 ;
wire un1_fracta_i_s0_cry_14 ;
wire un1_fracta_i_s0_cry_13 ;
wire un1_fracta_i_s0_cry_12 ;
wire un1_fracta_i_s0_cry_11 ;
wire un1_fracta_i_s0_cry_10 ;
wire un1_fracta_i_s0_cry_9 ;
wire un1_fracta_i_s0_cry_8 ;
wire un1_fracta_i_s0_cry_7 ;
wire un1_fracta_i_s0_cry_6 ;
wire un1_fracta_i_s0_cry_5 ;
wire un1_fracta_i_s0_cry_4 ;
wire un1_fracta_i_s0_cry_3 ;
wire un1_fracta_i_s0_cry_2 ;
wire un1_fracta_i_s0_cry_1 ;
wire un1_fracta_i_s0_cry_0 ;
wire un1_fracta_i_0_cry_26 ;
wire un1_fracta_i_0_cry_25 ;
wire un1_fracta_i_0_cry_24 ;
wire un1_fracta_i_0_cry_23 ;
wire un1_fracta_i_0_cry_22 ;
wire un1_fracta_i_0_cry_21 ;
wire un1_fracta_i_0_cry_20 ;
wire un1_fracta_i_0_cry_19 ;
wire un1_fracta_i_0_cry_18 ;
wire un1_fracta_i_0_cry_17 ;
wire un1_fracta_i_0_cry_16 ;
wire un1_fracta_i_0_cry_15 ;
wire un1_fracta_i_0_cry_14 ;
wire un1_fracta_i_0_cry_13 ;
wire un1_fracta_i_0_cry_12 ;
wire un1_fracta_i_0_cry_11 ;
wire un1_fracta_i_0_cry_10 ;
wire un1_fracta_i_0_cry_9 ;
wire un1_fracta_i_0_cry_8 ;
wire un1_fracta_i_0_cry_7 ;
wire un1_fracta_i_0_cry_6 ;
wire un1_fracta_i_0_cry_5 ;
wire un1_fracta_i_0_cry_4 ;
wire un1_fracta_i_0_cry_3 ;
wire un1_fracta_i_0_cry_2 ;
wire un1_fracta_i_0_cry_1 ;
wire un1_fracta_i_0_cry_0 ;
// instances
  LUT3 un1_fracta_i_s0_cry_0_cy_RNO_cZ(.I0(s_fpu_op_i),.I1(s_opa_i_27),.I2(s_opb_i_26),.O(un1_fracta_i_s0_cry_0_cy_RNO));
defparam un1_fracta_i_s0_cry_0_cy_RNO_cZ.INIT=8'h96;
  LUT3 un1_fracta_i_0_cry_0_cy_RNO_cZ(.I0(s_fpu_op_i),.I1(s_opa_i_27),.I2(s_opb_i_26),.O(un1_fracta_i_0_cry_0_cy_RNO));
defparam un1_fracta_i_0_cry_0_cy_RNO_cZ.INIT=8'h96;
  FD desc260(.Q(addsub_fract_o[14:14]),.D(N_2604_i),.C(clk_i));
  FD desc261(.Q(addsub_fract_o[15:15]),.D(N_2605_i),.C(clk_i));
  FD desc262(.Q(addsub_fract_o[16:16]),.D(N_2606_i),.C(clk_i));
  FD desc263(.Q(addsub_fract_o[17:17]),.D(N_2607_i),.C(clk_i));
  FD desc264(.Q(addsub_fract_o[18:18]),.D(N_2608_i),.C(clk_i));
  FD desc265(.Q(addsub_fract_o[19:19]),.D(N_2609_i),.C(clk_i));
  FD desc266(.Q(addsub_fract_o[20:20]),.D(N_2610_i),.C(clk_i));
  FD desc267(.Q(addsub_fract_o[21:21]),.D(N_2611_i),.C(clk_i));
  FD desc268(.Q(addsub_fract_o[22:22]),.D(N_2612_i),.C(clk_i));
  FD desc269(.Q(addsub_fract_o[23:23]),.D(N_2613_i),.C(clk_i));
  FD desc270(.Q(addsub_fract_o[24:24]),.D(N_2614_i),.C(clk_i));
  FD desc271(.Q(addsub_fract_o[25:25]),.D(N_2615_i),.C(clk_i));
  FD desc272(.Q(addsub_fract_o[26:26]),.D(N_2616_i),.C(clk_i));
  FD desc273(.Q(addsub_fract_o[27:27]),.D(N_2617_i),.C(clk_i));
  FD desc274(.Q(addsub_fract_o[0:0]),.D(N_2590_i),.C(clk_i));
  FD desc275(.Q(addsub_fract_o[1:1]),.D(N_2591_i),.C(clk_i));
  FD desc276(.Q(addsub_fract_o[2:2]),.D(N_59_0_i),.C(clk_i));
  FD desc277(.Q(addsub_fract_o[3:3]),.D(N_62_0_i),.C(clk_i));
  FD desc278(.Q(addsub_fract_o[4:4]),.D(N_65_0_i),.C(clk_i));
  FD desc279(.Q(addsub_fract_o[5:5]),.D(N_2595_i),.C(clk_i));
  FD desc280(.Q(addsub_fract_o[6:6]),.D(N_2596_i),.C(clk_i));
  FD desc281(.Q(addsub_fract_o[7:7]),.D(N_2597_i),.C(clk_i));
  FD desc282(.Q(addsub_fract_o[8:8]),.D(N_2598_i),.C(clk_i));
  FD desc283(.Q(addsub_fract_o[9:9]),.D(N_2599_i),.C(clk_i));
  FD desc284(.Q(addsub_fract_o[10:10]),.D(N_2600_i),.C(clk_i));
  FD desc285(.Q(addsub_fract_o[11:11]),.D(N_2601_i),.C(clk_i));
  FD desc286(.Q(addsub_fract_o[12:12]),.D(N_2602_i),.C(clk_i));
  FD desc287(.Q(addsub_fract_o[13:13]),.D(N_2603_i),.C(clk_i));
  MUXCY desc288(.DI(fracta_lt_fractb_lt26),.CI(fracta_lt_fractb_cry[24:24]),.S(fracta_lt_fractb_df26),.O(fracta_lt_fractb));
  LUT3 un1_fracta_i_0_s_27_RNO_cZ(.I0(s_fpu_op_i),.I1(s_opa_i_27),.I2(s_opb_i_26),.O(un1_fracta_i_0_s_27_RNO));
defparam un1_fracta_i_0_s_27_RNO_cZ.INIT=8'h96;
  LUT6_L sign_o_r(.I0(s_fpu_op_i),.I1(s_opa_i_27),.I2(s_opb_i_26),.I3(fracta_lt_fractb),.I4(un1_fracta_i_s0_s_14_RNID77E1_O6),.I5(m33_1_4),.LO(sign_o));
defparam sign_o_r.INIT=64'hC040CC5ACC5ACC5A;
  LUT6 m41_e(.I0(s_opb_i_1),.I1(s_opb_i_0),.I2(s_opb_i_2),.I3(result_2_2),.I4(N_1055),.I5(un1_s_infb),.O(N_1979));
defparam m41_e.INIT=64'hFFFEFFFF00000000;
  MUXCY_L un1_fracta_i_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_fracta_i_0_cry_0_cy_RNO),.LO(un1_fracta_i_0_cry_0_cy));
  MUXCY_L un1_fracta_i_s0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_fracta_i_s0_cry_0_cy_RNO),.LO(un1_fracta_i_s0_cry_0_cy));
  FD sign_o_Z(.Q(addsub_sign_o),.D(sign_o),.C(clk_i));
  LUT3 m49(.I0(s_fpu_op_i),.I1(s_opa_i_27),.I2(s_opb_i_26),.O(s_addop_1_1));
defparam m49.INIT=8'h96;
  LUT3_L desc289(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[18:18]),.I2(un1_fracta_i_11[18:18]),.LO(N_2608_i));
defparam desc289.INIT=8'hE4;
  LUT6_L sign_o_r_RNO_7(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[22:22]),.I2(un1_fracta_i_11[22:22]),.I3(un1_fracta_i_10[23:23]),.I4(un1_fracta_i_11[23:23]),.I5(m33_3_1),.LO(m33_3_3));
defparam sign_o_r_RNO_7.INIT=64'h00110A1B00000000;
  LUT6_L sign_o_r_RNO_6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[16:16]),.I2(un1_fracta_i_11[16:16]),.I3(un1_fracta_i_10[17:17]),.I4(un1_fracta_i_11[17:17]),.I5(m33_2_1),.LO(m33_2_3));
defparam sign_o_r_RNO_6.INIT=64'h00110A1B00000000;
  LUT6_L sign_o_r_RNO_5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[10:10]),.I2(un1_fracta_i_11[10:10]),.I3(un1_fracta_i_10[11:11]),.I4(un1_fracta_i_11[11:11]),.I5(m33_1_1),.LO(m33_1_3));
defparam sign_o_r_RNO_5.INIT=64'h00110A1B00000000;
  LUT6_L sign_o_r_RNO_4(.I0(un1_fracta_i_10[4:4]),.I1(un1_fracta_i_11[4:4]),.I2(un1_fracta_i_10[5:5]),.I3(un1_fracta_i_11[5:5]),.I4(fracta_lt_fractb),.I5(m33_0_1),.LO(m33_0_3));
defparam sign_o_r_RNO_4.INIT=64'h0033050500000000;
  LUT5 un1_fracta_i_s0_axb_26_cZ(.I0(prenorm_addsub_fracta_28_o[26:26]),.I1(prenorm_addsub_fractb_28_o[26:26]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_26));
defparam un1_fracta_i_s0_axb_26_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_25_cZ(.I0(prenorm_addsub_fracta_28_o[25:25]),.I1(prenorm_addsub_fractb_28_o[25:25]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_25));
defparam un1_fracta_i_s0_axb_25_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_24_cZ(.I0(prenorm_addsub_fracta_28_o[24:24]),.I1(prenorm_addsub_fractb_28_o[24:24]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_24));
defparam un1_fracta_i_s0_axb_24_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_23_cZ(.I0(prenorm_addsub_fracta_28_o[23:23]),.I1(prenorm_addsub_fractb_28_o[23:23]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_23));
defparam un1_fracta_i_s0_axb_23_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_22_cZ(.I0(prenorm_addsub_fracta_28_o[22:22]),.I1(prenorm_addsub_fractb_28_o[22:22]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_22));
defparam un1_fracta_i_s0_axb_22_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_21_cZ(.I0(prenorm_addsub_fracta_28_o[21:21]),.I1(prenorm_addsub_fractb_28_o[21:21]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_21));
defparam un1_fracta_i_s0_axb_21_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_20_cZ(.I0(prenorm_addsub_fracta_28_o[20:20]),.I1(prenorm_addsub_fractb_28_o[20:20]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_20));
defparam un1_fracta_i_s0_axb_20_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_19_cZ(.I0(prenorm_addsub_fracta_28_o[19:19]),.I1(prenorm_addsub_fractb_28_o[19:19]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_19));
defparam un1_fracta_i_s0_axb_19_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_18_cZ(.I0(prenorm_addsub_fracta_28_o[18:18]),.I1(prenorm_addsub_fractb_28_o[18:18]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_18));
defparam un1_fracta_i_s0_axb_18_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_17_cZ(.I0(prenorm_addsub_fracta_28_o[17:17]),.I1(prenorm_addsub_fractb_28_o[17:17]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_17));
defparam un1_fracta_i_s0_axb_17_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_16_cZ(.I0(prenorm_addsub_fracta_28_o[16:16]),.I1(prenorm_addsub_fractb_28_o[16:16]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_16));
defparam un1_fracta_i_s0_axb_16_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_15_cZ(.I0(prenorm_addsub_fracta_28_o[15:15]),.I1(prenorm_addsub_fractb_28_o[15:15]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_15));
defparam un1_fracta_i_s0_axb_15_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_14_cZ(.I0(prenorm_addsub_fracta_28_o[14:14]),.I1(prenorm_addsub_fractb_28_o[14:14]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_14));
defparam un1_fracta_i_s0_axb_14_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_13_cZ(.I0(prenorm_addsub_fracta_28_o[13:13]),.I1(prenorm_addsub_fractb_28_o[13:13]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_13));
defparam un1_fracta_i_s0_axb_13_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_12_cZ(.I0(prenorm_addsub_fracta_28_o[12:12]),.I1(prenorm_addsub_fractb_28_o[12:12]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_12));
defparam un1_fracta_i_s0_axb_12_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_11_cZ(.I0(prenorm_addsub_fracta_28_o[11:11]),.I1(prenorm_addsub_fractb_28_o[11:11]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_11));
defparam un1_fracta_i_s0_axb_11_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_10_cZ(.I0(prenorm_addsub_fracta_28_o[10:10]),.I1(prenorm_addsub_fractb_28_o[10:10]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_10));
defparam un1_fracta_i_s0_axb_10_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_9_cZ(.I0(prenorm_addsub_fracta_28_o[9:9]),.I1(prenorm_addsub_fractb_28_o[9:9]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_9));
defparam un1_fracta_i_s0_axb_9_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_8_cZ(.I0(prenorm_addsub_fracta_28_o[8:8]),.I1(prenorm_addsub_fractb_28_o[8:8]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_8));
defparam un1_fracta_i_s0_axb_8_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_7_cZ(.I0(prenorm_addsub_fracta_28_o[7:7]),.I1(prenorm_addsub_fractb_28_o[7:7]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_7));
defparam un1_fracta_i_s0_axb_7_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_6_cZ(.I0(prenorm_addsub_fracta_28_o[6:6]),.I1(prenorm_addsub_fractb_28_o[6:6]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_6));
defparam un1_fracta_i_s0_axb_6_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_5_cZ(.I0(prenorm_addsub_fracta_28_o[5:5]),.I1(prenorm_addsub_fractb_28_o[5:5]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_5));
defparam un1_fracta_i_s0_axb_5_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_4_cZ(.I0(prenorm_addsub_fracta_28_o[4:4]),.I1(prenorm_addsub_fractb_28_o[4:4]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_4));
defparam un1_fracta_i_s0_axb_4_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_3_cZ(.I0(prenorm_addsub_fracta_28_o[3:3]),.I1(prenorm_addsub_fractb_28_o[3:3]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_3));
defparam un1_fracta_i_s0_axb_3_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_2_cZ(.I0(prenorm_addsub_fracta_28_o[2:2]),.I1(prenorm_addsub_fractb_28_o[2:2]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_2));
defparam un1_fracta_i_s0_axb_2_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_1_cZ(.I0(prenorm_addsub_fracta_28_o[1:1]),.I1(prenorm_addsub_fractb_28_o[1:1]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_1));
defparam un1_fracta_i_s0_axb_1_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_s0_axb_0_cZ(.I0(prenorm_addsub_fracta_28_o[0:0]),.I1(prenorm_addsub_fractb_28_o[0:0]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_s0_axb_0));
defparam un1_fracta_i_s0_axb_0_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_26_cZ(.I0(prenorm_addsub_fracta_28_o[26:26]),.I1(prenorm_addsub_fractb_28_o[26:26]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_26));
defparam un1_fracta_i_0_axb_26_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_25_cZ(.I0(prenorm_addsub_fracta_28_o[25:25]),.I1(prenorm_addsub_fractb_28_o[25:25]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_25));
defparam un1_fracta_i_0_axb_25_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_24_cZ(.I0(prenorm_addsub_fracta_28_o[24:24]),.I1(prenorm_addsub_fractb_28_o[24:24]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_24));
defparam un1_fracta_i_0_axb_24_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_23_cZ(.I0(prenorm_addsub_fracta_28_o[23:23]),.I1(prenorm_addsub_fractb_28_o[23:23]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_23));
defparam un1_fracta_i_0_axb_23_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_22_cZ(.I0(prenorm_addsub_fracta_28_o[22:22]),.I1(prenorm_addsub_fractb_28_o[22:22]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_22));
defparam un1_fracta_i_0_axb_22_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_21_cZ(.I0(prenorm_addsub_fracta_28_o[21:21]),.I1(prenorm_addsub_fractb_28_o[21:21]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_21));
defparam un1_fracta_i_0_axb_21_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_20_cZ(.I0(prenorm_addsub_fracta_28_o[20:20]),.I1(prenorm_addsub_fractb_28_o[20:20]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_20));
defparam un1_fracta_i_0_axb_20_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_19_cZ(.I0(prenorm_addsub_fracta_28_o[19:19]),.I1(prenorm_addsub_fractb_28_o[19:19]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_19));
defparam un1_fracta_i_0_axb_19_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_18_cZ(.I0(prenorm_addsub_fracta_28_o[18:18]),.I1(prenorm_addsub_fractb_28_o[18:18]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_18));
defparam un1_fracta_i_0_axb_18_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_17_cZ(.I0(prenorm_addsub_fracta_28_o[17:17]),.I1(prenorm_addsub_fractb_28_o[17:17]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_17));
defparam un1_fracta_i_0_axb_17_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_16_cZ(.I0(prenorm_addsub_fracta_28_o[16:16]),.I1(prenorm_addsub_fractb_28_o[16:16]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_16));
defparam un1_fracta_i_0_axb_16_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_15_cZ(.I0(prenorm_addsub_fracta_28_o[15:15]),.I1(prenorm_addsub_fractb_28_o[15:15]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_15));
defparam un1_fracta_i_0_axb_15_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_14_cZ(.I0(prenorm_addsub_fracta_28_o[14:14]),.I1(prenorm_addsub_fractb_28_o[14:14]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_14));
defparam un1_fracta_i_0_axb_14_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_13_cZ(.I0(prenorm_addsub_fracta_28_o[13:13]),.I1(prenorm_addsub_fractb_28_o[13:13]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_13));
defparam un1_fracta_i_0_axb_13_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_12_cZ(.I0(prenorm_addsub_fracta_28_o[12:12]),.I1(prenorm_addsub_fractb_28_o[12:12]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_12));
defparam un1_fracta_i_0_axb_12_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_11_cZ(.I0(prenorm_addsub_fracta_28_o[11:11]),.I1(prenorm_addsub_fractb_28_o[11:11]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_11));
defparam un1_fracta_i_0_axb_11_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_10_cZ(.I0(prenorm_addsub_fracta_28_o[10:10]),.I1(prenorm_addsub_fractb_28_o[10:10]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_10));
defparam un1_fracta_i_0_axb_10_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_9_cZ(.I0(prenorm_addsub_fracta_28_o[9:9]),.I1(prenorm_addsub_fractb_28_o[9:9]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_9));
defparam un1_fracta_i_0_axb_9_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_8_cZ(.I0(prenorm_addsub_fracta_28_o[8:8]),.I1(prenorm_addsub_fractb_28_o[8:8]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_8));
defparam un1_fracta_i_0_axb_8_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_7_cZ(.I0(prenorm_addsub_fracta_28_o[7:7]),.I1(prenorm_addsub_fractb_28_o[7:7]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_7));
defparam un1_fracta_i_0_axb_7_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_6_cZ(.I0(prenorm_addsub_fracta_28_o[6:6]),.I1(prenorm_addsub_fractb_28_o[6:6]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_6));
defparam un1_fracta_i_0_axb_6_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_5_cZ(.I0(prenorm_addsub_fracta_28_o[5:5]),.I1(prenorm_addsub_fractb_28_o[5:5]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_5));
defparam un1_fracta_i_0_axb_5_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_4_cZ(.I0(prenorm_addsub_fracta_28_o[4:4]),.I1(prenorm_addsub_fractb_28_o[4:4]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_4));
defparam un1_fracta_i_0_axb_4_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_3_cZ(.I0(prenorm_addsub_fracta_28_o[3:3]),.I1(prenorm_addsub_fractb_28_o[3:3]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_3));
defparam un1_fracta_i_0_axb_3_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_2_cZ(.I0(prenorm_addsub_fracta_28_o[2:2]),.I1(prenorm_addsub_fractb_28_o[2:2]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_2));
defparam un1_fracta_i_0_axb_2_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_1_cZ(.I0(prenorm_addsub_fracta_28_o[1:1]),.I1(prenorm_addsub_fractb_28_o[1:1]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_1));
defparam un1_fracta_i_0_axb_1_cZ.INIT=32'h96696996;
  LUT5 un1_fracta_i_0_axb_0_cZ(.I0(prenorm_addsub_fracta_28_o[0:0]),.I1(prenorm_addsub_fractb_28_o[0:0]),.I2(s_fpu_op_i),.I3(s_opa_i_27),.I4(s_opb_i_26),.O(un1_fracta_i_0_axb_0));
defparam un1_fracta_i_0_axb_0_cZ.INIT=32'h96696996;
  LUT6_L sign_o_r_RNO_3(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[18:18]),.I2(un1_fracta_i_11[18:18]),.I3(un1_fracta_i_10[19:19]),.I4(un1_fracta_i_11[19:19]),.I5(m33_3_3),.LO(m33_3));
defparam sign_o_r_RNO_3.INIT=64'h00110A1B00000000;
  LUT6 sign_o_r_RNO_2(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[12:12]),.I2(un1_fracta_i_11[12:12]),.I3(un1_fracta_i_10[13:13]),.I4(un1_fracta_i_11[13:13]),.I5(m33_2_3),.O(m33_2));
defparam sign_o_r_RNO_2.INIT=64'h00110A1B00000000;
  LUT6 sign_o_r_RNO_1(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[6:6]),.I2(un1_fracta_i_11[6:6]),.I3(un1_fracta_i_10[7:7]),.I4(un1_fracta_i_11[7:7]),.I5(m33_1_3),.O(m33_1));
defparam sign_o_r_RNO_1.INIT=64'h00110A1B00000000;
  LUT6 sign_o_r_RNO_0(.I0(un1_fracta_i_10[0:0]),.I1(un1_fracta_i_11[0:0]),.I2(un1_fracta_i_10[1:1]),.I3(un1_fracta_i_11[1:1]),.I4(fracta_lt_fractb),.I5(m33_0_3),.O(m33_0));
defparam sign_o_r_RNO_0.INIT=64'h0033050500000000;
  LUT6 m35(.I0(s_opa_i_0),.I1(s_opa_i_1),.I2(un2_s_snan_o_8),.I3(N_1166),.I4(un4_s_infa),.I5(result_3_0_0_i),.O(N_36_0));
defparam m35.INIT=64'hFFEF0000FFFF0000;
  LUT6_L sign_o_r_RNO(.I0(un1_fracta_i_s0_s_24_RNI55IC1_O6),.I1(m33_4_1),.I2(m33_0),.I3(m33_1),.I4(m33_2),.I5(m33_3),.LO(m33_1_4));
defparam sign_o_r_RNO.INIT=64'h8000000000000000;
  LUT5 m48(.I0(s_addop_1_1),.I1(un4_s_infa),.I2(un1_s_infb),.I3(result_2),.I4(N_36_0),.O(N_1948));
defparam m48.INIT=32'h00200F7F;
  XORCY un1_fracta_i_s0_s_27(.LI(s_addop_1_1),.CI(un1_fracta_i_s0_cry_26),.O(un1_fracta_i_10[27:27]));
  XORCY un1_fracta_i_s0_s_26(.LI(un1_fracta_i_s0_axb_26),.CI(un1_fracta_i_s0_cry_25),.O(un1_fracta_i_10[26:26]));
  MUXCY_L un1_fracta_i_s0_cry_26_cZ(.DI(prenorm_addsub_fractb_28_o[26:26]),.CI(un1_fracta_i_s0_cry_25),.S(un1_fracta_i_s0_axb_26),.LO(un1_fracta_i_s0_cry_26));
  XORCY un1_fracta_i_s0_s_25(.LI(un1_fracta_i_s0_axb_25),.CI(un1_fracta_i_s0_cry_24),.O(un1_fracta_i_10[25:25]));
  MUXCY_L un1_fracta_i_s0_cry_25_cZ(.DI(prenorm_addsub_fractb_28_o[25:25]),.CI(un1_fracta_i_s0_cry_24),.S(un1_fracta_i_s0_axb_25),.LO(un1_fracta_i_s0_cry_25));
  XORCY un1_fracta_i_s0_s_24(.LI(un1_fracta_i_s0_axb_24),.CI(un1_fracta_i_s0_cry_23),.O(un1_fracta_i_10[24:24]));
  MUXCY_L un1_fracta_i_s0_cry_24_cZ(.DI(prenorm_addsub_fractb_28_o[24:24]),.CI(un1_fracta_i_s0_cry_23),.S(un1_fracta_i_s0_axb_24),.LO(un1_fracta_i_s0_cry_24));
  XORCY un1_fracta_i_s0_s_23(.LI(un1_fracta_i_s0_axb_23),.CI(un1_fracta_i_s0_cry_22),.O(un1_fracta_i_10[23:23]));
  MUXCY_L un1_fracta_i_s0_cry_23_cZ(.DI(prenorm_addsub_fractb_28_o[23:23]),.CI(un1_fracta_i_s0_cry_22),.S(un1_fracta_i_s0_axb_23),.LO(un1_fracta_i_s0_cry_23));
  XORCY un1_fracta_i_s0_s_22(.LI(un1_fracta_i_s0_axb_22),.CI(un1_fracta_i_s0_cry_21),.O(un1_fracta_i_10[22:22]));
  MUXCY_L un1_fracta_i_s0_cry_22_cZ(.DI(prenorm_addsub_fractb_28_o[22:22]),.CI(un1_fracta_i_s0_cry_21),.S(un1_fracta_i_s0_axb_22),.LO(un1_fracta_i_s0_cry_22));
  XORCY un1_fracta_i_s0_s_21(.LI(un1_fracta_i_s0_axb_21),.CI(un1_fracta_i_s0_cry_20),.O(un1_fracta_i_10[21:21]));
  MUXCY_L un1_fracta_i_s0_cry_21_cZ(.DI(prenorm_addsub_fractb_28_o[21:21]),.CI(un1_fracta_i_s0_cry_20),.S(un1_fracta_i_s0_axb_21),.LO(un1_fracta_i_s0_cry_21));
  XORCY un1_fracta_i_s0_s_20(.LI(un1_fracta_i_s0_axb_20),.CI(un1_fracta_i_s0_cry_19),.O(un1_fracta_i_10[20:20]));
  MUXCY_L un1_fracta_i_s0_cry_20_cZ(.DI(prenorm_addsub_fractb_28_o[20:20]),.CI(un1_fracta_i_s0_cry_19),.S(un1_fracta_i_s0_axb_20),.LO(un1_fracta_i_s0_cry_20));
  XORCY un1_fracta_i_s0_s_19(.LI(un1_fracta_i_s0_axb_19),.CI(un1_fracta_i_s0_cry_18),.O(un1_fracta_i_10[19:19]));
  MUXCY_L un1_fracta_i_s0_cry_19_cZ(.DI(prenorm_addsub_fractb_28_o[19:19]),.CI(un1_fracta_i_s0_cry_18),.S(un1_fracta_i_s0_axb_19),.LO(un1_fracta_i_s0_cry_19));
  XORCY un1_fracta_i_s0_s_18(.LI(un1_fracta_i_s0_axb_18),.CI(un1_fracta_i_s0_cry_17),.O(un1_fracta_i_10[18:18]));
  MUXCY_L un1_fracta_i_s0_cry_18_cZ(.DI(prenorm_addsub_fractb_28_o[18:18]),.CI(un1_fracta_i_s0_cry_17),.S(un1_fracta_i_s0_axb_18),.LO(un1_fracta_i_s0_cry_18));
  XORCY un1_fracta_i_s0_s_17(.LI(un1_fracta_i_s0_axb_17),.CI(un1_fracta_i_s0_cry_16),.O(un1_fracta_i_10[17:17]));
  MUXCY_L un1_fracta_i_s0_cry_17_cZ(.DI(prenorm_addsub_fractb_28_o[17:17]),.CI(un1_fracta_i_s0_cry_16),.S(un1_fracta_i_s0_axb_17),.LO(un1_fracta_i_s0_cry_17));
  XORCY un1_fracta_i_s0_s_16(.LI(un1_fracta_i_s0_axb_16),.CI(un1_fracta_i_s0_cry_15),.O(un1_fracta_i_10[16:16]));
  MUXCY_L un1_fracta_i_s0_cry_16_cZ(.DI(prenorm_addsub_fractb_28_o[16:16]),.CI(un1_fracta_i_s0_cry_15),.S(un1_fracta_i_s0_axb_16),.LO(un1_fracta_i_s0_cry_16));
  XORCY un1_fracta_i_s0_s_15(.LI(un1_fracta_i_s0_axb_15),.CI(un1_fracta_i_s0_cry_14),.O(un1_fracta_i_10[15:15]));
  MUXCY_L un1_fracta_i_s0_cry_15_cZ(.DI(prenorm_addsub_fractb_28_o[15:15]),.CI(un1_fracta_i_s0_cry_14),.S(un1_fracta_i_s0_axb_15),.LO(un1_fracta_i_s0_cry_15));
  XORCY un1_fracta_i_s0_s_14(.LI(un1_fracta_i_s0_axb_14),.CI(un1_fracta_i_s0_cry_13),.O(un1_fracta_i_10[14:14]));
  MUXCY_L un1_fracta_i_s0_cry_14_cZ(.DI(prenorm_addsub_fractb_28_o[14:14]),.CI(un1_fracta_i_s0_cry_13),.S(un1_fracta_i_s0_axb_14),.LO(un1_fracta_i_s0_cry_14));
  XORCY un1_fracta_i_s0_s_13(.LI(un1_fracta_i_s0_axb_13),.CI(un1_fracta_i_s0_cry_12),.O(un1_fracta_i_10[13:13]));
  MUXCY_L un1_fracta_i_s0_cry_13_cZ(.DI(prenorm_addsub_fractb_28_o[13:13]),.CI(un1_fracta_i_s0_cry_12),.S(un1_fracta_i_s0_axb_13),.LO(un1_fracta_i_s0_cry_13));
  XORCY un1_fracta_i_s0_s_12(.LI(un1_fracta_i_s0_axb_12),.CI(un1_fracta_i_s0_cry_11),.O(un1_fracta_i_10[12:12]));
  MUXCY_L un1_fracta_i_s0_cry_12_cZ(.DI(prenorm_addsub_fractb_28_o[12:12]),.CI(un1_fracta_i_s0_cry_11),.S(un1_fracta_i_s0_axb_12),.LO(un1_fracta_i_s0_cry_12));
  XORCY un1_fracta_i_s0_s_11(.LI(un1_fracta_i_s0_axb_11),.CI(un1_fracta_i_s0_cry_10),.O(un1_fracta_i_10[11:11]));
  MUXCY_L un1_fracta_i_s0_cry_11_cZ(.DI(prenorm_addsub_fractb_28_o[11:11]),.CI(un1_fracta_i_s0_cry_10),.S(un1_fracta_i_s0_axb_11),.LO(un1_fracta_i_s0_cry_11));
  XORCY un1_fracta_i_s0_s_10(.LI(un1_fracta_i_s0_axb_10),.CI(un1_fracta_i_s0_cry_9),.O(un1_fracta_i_10[10:10]));
  MUXCY_L un1_fracta_i_s0_cry_10_cZ(.DI(prenorm_addsub_fractb_28_o[10:10]),.CI(un1_fracta_i_s0_cry_9),.S(un1_fracta_i_s0_axb_10),.LO(un1_fracta_i_s0_cry_10));
  XORCY un1_fracta_i_s0_s_9(.LI(un1_fracta_i_s0_axb_9),.CI(un1_fracta_i_s0_cry_8),.O(un1_fracta_i_10[9:9]));
  MUXCY_L un1_fracta_i_s0_cry_9_cZ(.DI(prenorm_addsub_fractb_28_o[9:9]),.CI(un1_fracta_i_s0_cry_8),.S(un1_fracta_i_s0_axb_9),.LO(un1_fracta_i_s0_cry_9));
  XORCY un1_fracta_i_s0_s_8(.LI(un1_fracta_i_s0_axb_8),.CI(un1_fracta_i_s0_cry_7),.O(un1_fracta_i_10[8:8]));
  MUXCY_L un1_fracta_i_s0_cry_8_cZ(.DI(prenorm_addsub_fractb_28_o[8:8]),.CI(un1_fracta_i_s0_cry_7),.S(un1_fracta_i_s0_axb_8),.LO(un1_fracta_i_s0_cry_8));
  XORCY un1_fracta_i_s0_s_7(.LI(un1_fracta_i_s0_axb_7),.CI(un1_fracta_i_s0_cry_6),.O(un1_fracta_i_10[7:7]));
  MUXCY_L un1_fracta_i_s0_cry_7_cZ(.DI(prenorm_addsub_fractb_28_o[7:7]),.CI(un1_fracta_i_s0_cry_6),.S(un1_fracta_i_s0_axb_7),.LO(un1_fracta_i_s0_cry_7));
  XORCY un1_fracta_i_s0_s_6(.LI(un1_fracta_i_s0_axb_6),.CI(un1_fracta_i_s0_cry_5),.O(un1_fracta_i_10[6:6]));
  MUXCY_L un1_fracta_i_s0_cry_6_cZ(.DI(prenorm_addsub_fractb_28_o[6:6]),.CI(un1_fracta_i_s0_cry_5),.S(un1_fracta_i_s0_axb_6),.LO(un1_fracta_i_s0_cry_6));
  XORCY un1_fracta_i_s0_s_5(.LI(un1_fracta_i_s0_axb_5),.CI(un1_fracta_i_s0_cry_4),.O(un1_fracta_i_10[5:5]));
  MUXCY_L un1_fracta_i_s0_cry_5_cZ(.DI(prenorm_addsub_fractb_28_o[5:5]),.CI(un1_fracta_i_s0_cry_4),.S(un1_fracta_i_s0_axb_5),.LO(un1_fracta_i_s0_cry_5));
  XORCY un1_fracta_i_s0_s_4(.LI(un1_fracta_i_s0_axb_4),.CI(un1_fracta_i_s0_cry_3),.O(un1_fracta_i_10[4:4]));
  MUXCY_L un1_fracta_i_s0_cry_4_cZ(.DI(prenorm_addsub_fractb_28_o[4:4]),.CI(un1_fracta_i_s0_cry_3),.S(un1_fracta_i_s0_axb_4),.LO(un1_fracta_i_s0_cry_4));
  XORCY un1_fracta_i_s0_s_3(.LI(un1_fracta_i_s0_axb_3),.CI(un1_fracta_i_s0_cry_2),.O(un1_fracta_i_10[3:3]));
  MUXCY_L un1_fracta_i_s0_cry_3_cZ(.DI(prenorm_addsub_fractb_28_o[3:3]),.CI(un1_fracta_i_s0_cry_2),.S(un1_fracta_i_s0_axb_3),.LO(un1_fracta_i_s0_cry_3));
  XORCY un1_fracta_i_s0_s_2(.LI(un1_fracta_i_s0_axb_2),.CI(un1_fracta_i_s0_cry_1),.O(un1_fracta_i_10[2:2]));
  MUXCY_L un1_fracta_i_s0_cry_2_cZ(.DI(prenorm_addsub_fractb_28_o[2:2]),.CI(un1_fracta_i_s0_cry_1),.S(un1_fracta_i_s0_axb_2),.LO(un1_fracta_i_s0_cry_2));
  XORCY un1_fracta_i_s0_s_1(.LI(un1_fracta_i_s0_axb_1),.CI(un1_fracta_i_s0_cry_0),.O(un1_fracta_i_10[1:1]));
  MUXCY_L un1_fracta_i_s0_cry_1_cZ(.DI(prenorm_addsub_fractb_28_o[1:1]),.CI(un1_fracta_i_s0_cry_0),.S(un1_fracta_i_s0_axb_1),.LO(un1_fracta_i_s0_cry_1));
  XORCY un1_fracta_i_s0_s_0(.LI(un1_fracta_i_s0_axb_0),.CI(un1_fracta_i_s0_cry_0_cy),.O(un1_fracta_i_10[0:0]));
  MUXCY_L un1_fracta_i_s0_cry_0_cZ(.DI(prenorm_addsub_fractb_28_o[0:0]),.CI(un1_fracta_i_s0_cry_0_cy),.S(un1_fracta_i_s0_axb_0),.LO(un1_fracta_i_s0_cry_0));
  XORCY un1_fracta_i_0_s_27(.LI(un1_fracta_i_0_s_27_RNO),.CI(un1_fracta_i_0_cry_26),.O(un1_fracta_i_11[27:27]));
  XORCY un1_fracta_i_0_s_26(.LI(un1_fracta_i_0_axb_26),.CI(un1_fracta_i_0_cry_25),.O(un1_fracta_i_11[26:26]));
  MUXCY_L un1_fracta_i_0_cry_26_cZ(.DI(prenorm_addsub_fracta_28_o[26:26]),.CI(un1_fracta_i_0_cry_25),.S(un1_fracta_i_0_axb_26),.LO(un1_fracta_i_0_cry_26));
  XORCY un1_fracta_i_0_s_25(.LI(un1_fracta_i_0_axb_25),.CI(un1_fracta_i_0_cry_24),.O(un1_fracta_i_11[25:25]));
  MUXCY_L un1_fracta_i_0_cry_25_cZ(.DI(prenorm_addsub_fracta_28_o[25:25]),.CI(un1_fracta_i_0_cry_24),.S(un1_fracta_i_0_axb_25),.LO(un1_fracta_i_0_cry_25));
  XORCY un1_fracta_i_0_s_24(.LI(un1_fracta_i_0_axb_24),.CI(un1_fracta_i_0_cry_23),.O(un1_fracta_i_11[24:24]));
  MUXCY_L un1_fracta_i_0_cry_24_cZ(.DI(prenorm_addsub_fracta_28_o[24:24]),.CI(un1_fracta_i_0_cry_23),.S(un1_fracta_i_0_axb_24),.LO(un1_fracta_i_0_cry_24));
  XORCY un1_fracta_i_0_s_23(.LI(un1_fracta_i_0_axb_23),.CI(un1_fracta_i_0_cry_22),.O(un1_fracta_i_11[23:23]));
  MUXCY_L un1_fracta_i_0_cry_23_cZ(.DI(prenorm_addsub_fracta_28_o[23:23]),.CI(un1_fracta_i_0_cry_22),.S(un1_fracta_i_0_axb_23),.LO(un1_fracta_i_0_cry_23));
  XORCY un1_fracta_i_0_s_22(.LI(un1_fracta_i_0_axb_22),.CI(un1_fracta_i_0_cry_21),.O(un1_fracta_i_11[22:22]));
  MUXCY_L un1_fracta_i_0_cry_22_cZ(.DI(prenorm_addsub_fracta_28_o[22:22]),.CI(un1_fracta_i_0_cry_21),.S(un1_fracta_i_0_axb_22),.LO(un1_fracta_i_0_cry_22));
  XORCY un1_fracta_i_0_s_21(.LI(un1_fracta_i_0_axb_21),.CI(un1_fracta_i_0_cry_20),.O(un1_fracta_i_11[21:21]));
  MUXCY_L un1_fracta_i_0_cry_21_cZ(.DI(prenorm_addsub_fracta_28_o[21:21]),.CI(un1_fracta_i_0_cry_20),.S(un1_fracta_i_0_axb_21),.LO(un1_fracta_i_0_cry_21));
  XORCY un1_fracta_i_0_s_20(.LI(un1_fracta_i_0_axb_20),.CI(un1_fracta_i_0_cry_19),.O(un1_fracta_i_11[20:20]));
  MUXCY_L un1_fracta_i_0_cry_20_cZ(.DI(prenorm_addsub_fracta_28_o[20:20]),.CI(un1_fracta_i_0_cry_19),.S(un1_fracta_i_0_axb_20),.LO(un1_fracta_i_0_cry_20));
  XORCY un1_fracta_i_0_s_19(.LI(un1_fracta_i_0_axb_19),.CI(un1_fracta_i_0_cry_18),.O(un1_fracta_i_11[19:19]));
  MUXCY_L un1_fracta_i_0_cry_19_cZ(.DI(prenorm_addsub_fracta_28_o[19:19]),.CI(un1_fracta_i_0_cry_18),.S(un1_fracta_i_0_axb_19),.LO(un1_fracta_i_0_cry_19));
  XORCY un1_fracta_i_0_s_18(.LI(un1_fracta_i_0_axb_18),.CI(un1_fracta_i_0_cry_17),.O(un1_fracta_i_11[18:18]));
  MUXCY_L un1_fracta_i_0_cry_18_cZ(.DI(prenorm_addsub_fracta_28_o[18:18]),.CI(un1_fracta_i_0_cry_17),.S(un1_fracta_i_0_axb_18),.LO(un1_fracta_i_0_cry_18));
  XORCY un1_fracta_i_0_s_17(.LI(un1_fracta_i_0_axb_17),.CI(un1_fracta_i_0_cry_16),.O(un1_fracta_i_11[17:17]));
  MUXCY_L un1_fracta_i_0_cry_17_cZ(.DI(prenorm_addsub_fracta_28_o[17:17]),.CI(un1_fracta_i_0_cry_16),.S(un1_fracta_i_0_axb_17),.LO(un1_fracta_i_0_cry_17));
  XORCY un1_fracta_i_0_s_16(.LI(un1_fracta_i_0_axb_16),.CI(un1_fracta_i_0_cry_15),.O(un1_fracta_i_11[16:16]));
  MUXCY_L un1_fracta_i_0_cry_16_cZ(.DI(prenorm_addsub_fracta_28_o[16:16]),.CI(un1_fracta_i_0_cry_15),.S(un1_fracta_i_0_axb_16),.LO(un1_fracta_i_0_cry_16));
  XORCY un1_fracta_i_0_s_15(.LI(un1_fracta_i_0_axb_15),.CI(un1_fracta_i_0_cry_14),.O(un1_fracta_i_11[15:15]));
  MUXCY_L un1_fracta_i_0_cry_15_cZ(.DI(prenorm_addsub_fracta_28_o[15:15]),.CI(un1_fracta_i_0_cry_14),.S(un1_fracta_i_0_axb_15),.LO(un1_fracta_i_0_cry_15));
  XORCY un1_fracta_i_0_s_14(.LI(un1_fracta_i_0_axb_14),.CI(un1_fracta_i_0_cry_13),.O(un1_fracta_i_11[14:14]));
  MUXCY_L un1_fracta_i_0_cry_14_cZ(.DI(prenorm_addsub_fracta_28_o[14:14]),.CI(un1_fracta_i_0_cry_13),.S(un1_fracta_i_0_axb_14),.LO(un1_fracta_i_0_cry_14));
  XORCY un1_fracta_i_0_s_13(.LI(un1_fracta_i_0_axb_13),.CI(un1_fracta_i_0_cry_12),.O(un1_fracta_i_11[13:13]));
  MUXCY_L un1_fracta_i_0_cry_13_cZ(.DI(prenorm_addsub_fracta_28_o[13:13]),.CI(un1_fracta_i_0_cry_12),.S(un1_fracta_i_0_axb_13),.LO(un1_fracta_i_0_cry_13));
  XORCY un1_fracta_i_0_s_12(.LI(un1_fracta_i_0_axb_12),.CI(un1_fracta_i_0_cry_11),.O(un1_fracta_i_11[12:12]));
  MUXCY_L un1_fracta_i_0_cry_12_cZ(.DI(prenorm_addsub_fracta_28_o[12:12]),.CI(un1_fracta_i_0_cry_11),.S(un1_fracta_i_0_axb_12),.LO(un1_fracta_i_0_cry_12));
  XORCY un1_fracta_i_0_s_11(.LI(un1_fracta_i_0_axb_11),.CI(un1_fracta_i_0_cry_10),.O(un1_fracta_i_11[11:11]));
  MUXCY_L un1_fracta_i_0_cry_11_cZ(.DI(prenorm_addsub_fracta_28_o[11:11]),.CI(un1_fracta_i_0_cry_10),.S(un1_fracta_i_0_axb_11),.LO(un1_fracta_i_0_cry_11));
  XORCY un1_fracta_i_0_s_10(.LI(un1_fracta_i_0_axb_10),.CI(un1_fracta_i_0_cry_9),.O(un1_fracta_i_11[10:10]));
  MUXCY_L un1_fracta_i_0_cry_10_cZ(.DI(prenorm_addsub_fracta_28_o[10:10]),.CI(un1_fracta_i_0_cry_9),.S(un1_fracta_i_0_axb_10),.LO(un1_fracta_i_0_cry_10));
  XORCY un1_fracta_i_0_s_9(.LI(un1_fracta_i_0_axb_9),.CI(un1_fracta_i_0_cry_8),.O(un1_fracta_i_11[9:9]));
  MUXCY_L un1_fracta_i_0_cry_9_cZ(.DI(prenorm_addsub_fracta_28_o[9:9]),.CI(un1_fracta_i_0_cry_8),.S(un1_fracta_i_0_axb_9),.LO(un1_fracta_i_0_cry_9));
  XORCY un1_fracta_i_0_s_8(.LI(un1_fracta_i_0_axb_8),.CI(un1_fracta_i_0_cry_7),.O(un1_fracta_i_11[8:8]));
  MUXCY_L un1_fracta_i_0_cry_8_cZ(.DI(prenorm_addsub_fracta_28_o[8:8]),.CI(un1_fracta_i_0_cry_7),.S(un1_fracta_i_0_axb_8),.LO(un1_fracta_i_0_cry_8));
  XORCY un1_fracta_i_0_s_7(.LI(un1_fracta_i_0_axb_7),.CI(un1_fracta_i_0_cry_6),.O(un1_fracta_i_11[7:7]));
  MUXCY_L un1_fracta_i_0_cry_7_cZ(.DI(prenorm_addsub_fracta_28_o[7:7]),.CI(un1_fracta_i_0_cry_6),.S(un1_fracta_i_0_axb_7),.LO(un1_fracta_i_0_cry_7));
  XORCY un1_fracta_i_0_s_6(.LI(un1_fracta_i_0_axb_6),.CI(un1_fracta_i_0_cry_5),.O(un1_fracta_i_11[6:6]));
  MUXCY_L un1_fracta_i_0_cry_6_cZ(.DI(prenorm_addsub_fracta_28_o[6:6]),.CI(un1_fracta_i_0_cry_5),.S(un1_fracta_i_0_axb_6),.LO(un1_fracta_i_0_cry_6));
  XORCY un1_fracta_i_0_s_5(.LI(un1_fracta_i_0_axb_5),.CI(un1_fracta_i_0_cry_4),.O(un1_fracta_i_11[5:5]));
  MUXCY_L un1_fracta_i_0_cry_5_cZ(.DI(prenorm_addsub_fracta_28_o[5:5]),.CI(un1_fracta_i_0_cry_4),.S(un1_fracta_i_0_axb_5),.LO(un1_fracta_i_0_cry_5));
  XORCY un1_fracta_i_0_s_4(.LI(un1_fracta_i_0_axb_4),.CI(un1_fracta_i_0_cry_3),.O(un1_fracta_i_11[4:4]));
  MUXCY_L un1_fracta_i_0_cry_4_cZ(.DI(prenorm_addsub_fracta_28_o[4:4]),.CI(un1_fracta_i_0_cry_3),.S(un1_fracta_i_0_axb_4),.LO(un1_fracta_i_0_cry_4));
  XORCY un1_fracta_i_0_s_3(.LI(un1_fracta_i_0_axb_3),.CI(un1_fracta_i_0_cry_2),.O(un1_fracta_i_11[3:3]));
  MUXCY_L un1_fracta_i_0_cry_3_cZ(.DI(prenorm_addsub_fracta_28_o[3:3]),.CI(un1_fracta_i_0_cry_2),.S(un1_fracta_i_0_axb_3),.LO(un1_fracta_i_0_cry_3));
  XORCY un1_fracta_i_0_s_2(.LI(un1_fracta_i_0_axb_2),.CI(un1_fracta_i_0_cry_1),.O(un1_fracta_i_11[2:2]));
  MUXCY_L un1_fracta_i_0_cry_2_cZ(.DI(prenorm_addsub_fracta_28_o[2:2]),.CI(un1_fracta_i_0_cry_1),.S(un1_fracta_i_0_axb_2),.LO(un1_fracta_i_0_cry_2));
  XORCY un1_fracta_i_0_s_1(.LI(un1_fracta_i_0_axb_1),.CI(un1_fracta_i_0_cry_0),.O(un1_fracta_i_11[1:1]));
  MUXCY_L un1_fracta_i_0_cry_1_cZ(.DI(prenorm_addsub_fracta_28_o[1:1]),.CI(un1_fracta_i_0_cry_0),.S(un1_fracta_i_0_axb_1),.LO(un1_fracta_i_0_cry_1));
  XORCY un1_fracta_i_0_s_0(.LI(un1_fracta_i_0_axb_0),.CI(un1_fracta_i_0_cry_0_cy),.O(un1_fracta_i_11[0:0]));
  MUXCY_L un1_fracta_i_0_cry_0_cZ(.DI(prenorm_addsub_fracta_28_o[0:0]),.CI(un1_fracta_i_0_cry_0_cy),.S(un1_fracta_i_0_axb_0),.LO(un1_fracta_i_0_cry_0));
  MUXCY_L desc290(.DI(fracta_lt_fractb_lt24),.CI(fracta_lt_fractb_cry[22:22]),.S(fracta_lt_fractb_df24),.LO(fracta_lt_fractb_cry[24:24]));
  MUXCY_L desc291(.DI(fracta_lt_fractb_lt22),.CI(fracta_lt_fractb_cry[20:20]),.S(fracta_lt_fractb_df22),.LO(fracta_lt_fractb_cry[22:22]));
  MUXCY_L desc292(.DI(fracta_lt_fractb_lt20),.CI(fracta_lt_fractb_cry[18:18]),.S(fracta_lt_fractb_df20),.LO(fracta_lt_fractb_cry[20:20]));
  MUXCY_L desc293(.DI(fracta_lt_fractb_lt18),.CI(fracta_lt_fractb_cry[16:16]),.S(fracta_lt_fractb_df18),.LO(fracta_lt_fractb_cry[18:18]));
  MUXCY_L desc294(.DI(fracta_lt_fractb_lt16),.CI(fracta_lt_fractb_cry[14:14]),.S(fracta_lt_fractb_df16),.LO(fracta_lt_fractb_cry[16:16]));
  MUXCY_L desc295(.DI(fracta_lt_fractb_lt14),.CI(fracta_lt_fractb_cry[12:12]),.S(fracta_lt_fractb_df14),.LO(fracta_lt_fractb_cry[14:14]));
  MUXCY_L desc296(.DI(fracta_lt_fractb_lt12),.CI(fracta_lt_fractb_cry[10:10]),.S(fracta_lt_fractb_df12),.LO(fracta_lt_fractb_cry[12:12]));
  MUXCY_L desc297(.DI(fracta_lt_fractb_lt10),.CI(fracta_lt_fractb_cry[8:8]),.S(fracta_lt_fractb_df10),.LO(fracta_lt_fractb_cry[10:10]));
  MUXCY_L desc298(.DI(fracta_lt_fractb_lt8),.CI(fracta_lt_fractb_cry[6:6]),.S(fracta_lt_fractb_df8),.LO(fracta_lt_fractb_cry[8:8]));
  MUXCY_L desc299(.DI(fracta_lt_fractb_lt6),.CI(fracta_lt_fractb_cry[4:4]),.S(fracta_lt_fractb_df6),.LO(fracta_lt_fractb_cry[6:6]));
  MUXCY_L desc300(.DI(fracta_lt_fractb_lt4),.CI(fracta_lt_fractb_cry[2:2]),.S(fracta_lt_fractb_df4),.LO(fracta_lt_fractb_cry[4:4]));
  MUXCY_L desc301(.DI(fracta_lt_fractb_lt2),.CI(fracta_lt_fractb_cry[0:0]),.S(fracta_lt_fractb_df2),.LO(fracta_lt_fractb_cry[2:2]));
  MUXCY_L desc302(.DI(fracta_lt_fractb_lt0),.CI(GND),.S(fracta_lt_fractb_df0),.LO(fracta_lt_fractb_cry[0:0]));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT2 m1_lut6_2_o6(.I0(s_fpu_op_i),.I1(s_opb_i_26),.O(N_1941));
defparam m1_lut6_2_o6.INIT=4'h9;
  LUT2 m1_lut6_2_o5(.I0(s_opa_i_27),.I1(s_opb_i_26),.O(N_1942_i));
defparam m1_lut6_2_o5.INIT=4'h6;
  LUT3 un1_fracta_i_s0_s_13_RNIB3IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[9:9]),.I2(un1_fracta_i_11[9:9]),.O(N_2599_i));
defparam un1_fracta_i_s0_s_13_RNIB3IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_13_RNIB3IC1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[13:13]),.I2(un1_fracta_i_11[13:13]),.O(N_2603_i));
defparam un1_fracta_i_s0_s_13_RNIB3IC1_o5.INIT=8'hE4;
  LUT5 un1_fracta_i_0_s_8_RNIJ1TA1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[8:8]),.I2(un1_fracta_i_11[8:8]),.I3(un1_fracta_i_10[9:9]),.I4(un1_fracta_i_11[9:9]),.O(m33_1_1));
defparam un1_fracta_i_0_s_8_RNIJ1TA1_o6.INIT=32'h00110A1B;
  LUT3 un1_fracta_i_0_s_8_RNIJ1TA1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[8:8]),.I2(un1_fracta_i_11[8:8]),.O(N_2598_i));
defparam un1_fracta_i_0_s_8_RNIJ1TA1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_12_RNI53IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[7:7]),.I2(un1_fracta_i_11[7:7]),.O(N_2597_i));
defparam un1_fracta_i_s0_s_12_RNI53IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_12_RNI53IC1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[12:12]),.I2(un1_fracta_i_11[12:12]),.O(N_2602_i));
defparam un1_fracta_i_s0_s_12_RNI53IC1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_11_RNI13IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[6:6]),.I2(un1_fracta_i_11[6:6]),.O(N_2596_i));
defparam un1_fracta_i_s0_s_11_RNI13IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_11_RNI13IC1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[11:11]),.I2(un1_fracta_i_11[11:11]),.O(N_2601_i));
defparam un1_fracta_i_s0_s_11_RNI13IC1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_10_RNIT2IC1_o6(.I0(un1_fracta_i_10[5:5]),.I1(un1_fracta_i_11[5:5]),.I2(fracta_lt_fractb),.O(N_2595_i));
defparam un1_fracta_i_s0_s_10_RNIT2IC1_o6.INIT=8'hCA;
  LUT3 un1_fracta_i_s0_s_10_RNIT2IC1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[10:10]),.I2(un1_fracta_i_11[10:10]),.O(N_2600_i));
defparam un1_fracta_i_s0_s_10_RNIT2IC1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_24_RNI55IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[24:24]),.I2(un1_fracta_i_11[24:24]),.O(un1_fracta_i_s0_s_24_RNI55IC1_O6));
defparam un1_fracta_i_s0_s_24_RNI55IC1_o6.INIT=8'h1B;
  LUT3 un1_fracta_i_s0_s_24_RNI55IC1_o5(.I0(un1_fracta_i_10[4:4]),.I1(un1_fracta_i_11[4:4]),.I2(fracta_lt_fractb),.O(N_65_0_i));
defparam un1_fracta_i_s0_s_24_RNI55IC1_o5.INIT=8'hCA;
  LUT5 un1_fracta_i_0_s_3_RNIR0TA1_o6(.I0(un1_fracta_i_10[2:2]),.I1(un1_fracta_i_11[2:2]),.I2(un1_fracta_i_10[3:3]),.I3(un1_fracta_i_11[3:3]),.I4(fracta_lt_fractb),.O(m33_0_1));
defparam un1_fracta_i_0_s_3_RNIR0TA1_o6.INIT=32'h00330505;
  LUT3 un1_fracta_i_0_s_3_RNIR0TA1_o5(.I0(un1_fracta_i_10[3:3]),.I1(un1_fracta_i_11[3:3]),.I2(fracta_lt_fractb),.O(N_62_0_i));
defparam un1_fracta_i_0_s_3_RNIR0TA1_o5.INIT=8'hCA;
  LUT3 un1_fracta_i_s0_s_27_RNI55IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[27:27]),.I2(un1_fracta_i_11[27:27]),.O(N_2617_i));
defparam un1_fracta_i_s0_s_27_RNI55IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_27_RNI55IC1_o5(.I0(un1_fracta_i_10[1:1]),.I1(un1_fracta_i_11[1:1]),.I2(fracta_lt_fractb),.O(N_2591_i));
defparam un1_fracta_i_s0_s_27_RNI55IC1_o5.INIT=8'hCA;
  LUT3 un1_fracta_i_s0_s_26_RNI15IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[26:26]),.I2(un1_fracta_i_11[26:26]),.O(N_2616_i));
defparam un1_fracta_i_s0_s_26_RNI15IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_26_RNI15IC1_o5(.I0(un1_fracta_i_10[0:0]),.I1(un1_fracta_i_11[0:0]),.I2(fracta_lt_fractb),.O(N_2590_i));
defparam un1_fracta_i_s0_s_26_RNI15IC1_o5.INIT=8'hCA;
  LUT5 un1_fracta_i_s0_s_25_RNIF97E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[25:25]),.I2(un1_fracta_i_11[25:25]),.I3(un1_fracta_i_10[26:26]),.I4(un1_fracta_i_11[26:26]),.O(m33_4_1));
defparam un1_fracta_i_s0_s_25_RNIF97E1_o6.INIT=32'h00110A1B;
  LUT3 un1_fracta_i_s0_s_25_RNIF97E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[25:25]),.I2(un1_fracta_i_11[25:25]),.O(N_2615_i));
defparam un1_fracta_i_s0_s_25_RNIF97E1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_22_RNI597E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[22:22]),.I2(un1_fracta_i_11[22:22]),.O(N_2612_i));
defparam un1_fracta_i_s0_s_22_RNI597E1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_22_RNI597E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[24:24]),.I2(un1_fracta_i_11[24:24]),.O(N_2614_i));
defparam un1_fracta_i_s0_s_22_RNI597E1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_21_RNI197E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[21:21]),.I2(un1_fracta_i_11[21:21]),.O(N_2611_i));
defparam un1_fracta_i_s0_s_21_RNI197E1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_21_RNI197E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[23:23]),.I2(un1_fracta_i_11[23:23]),.O(N_2613_i));
defparam un1_fracta_i_s0_s_21_RNI197E1_o5.INIT=8'hE4;
  LUT5 un1_fracta_i_s0_s_20_RNIR87E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[20:20]),.I2(un1_fracta_i_11[20:20]),.I3(un1_fracta_i_10[21:21]),.I4(un1_fracta_i_11[21:21]),.O(m33_3_1));
defparam un1_fracta_i_s0_s_20_RNIR87E1_o6.INIT=32'h00110A1B;
  LUT3 un1_fracta_i_s0_s_20_RNIR87E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[20:20]),.I2(un1_fracta_i_11[20:20]),.O(N_2610_i));
defparam un1_fracta_i_s0_s_20_RNIR87E1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_17_RNIL57E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[17:17]),.I2(un1_fracta_i_11[17:17]),.O(N_2607_i));
defparam un1_fracta_i_s0_s_17_RNIL57E1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_17_RNIL57E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[19:19]),.I2(un1_fracta_i_11[19:19]),.O(N_2609_i));
defparam un1_fracta_i_s0_s_17_RNIL57E1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_16_RNI33IC1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[16:16]),.I2(un1_fracta_i_11[16:16]),.O(N_2606_i));
defparam un1_fracta_i_s0_s_16_RNI33IC1_o6.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_16_RNI33IC1_o5(.I0(un1_fracta_i_10[2:2]),.I1(un1_fracta_i_11[2:2]),.I2(fracta_lt_fractb),.O(N_59_0_i));
defparam un1_fracta_i_s0_s_16_RNI33IC1_o5.INIT=8'hCA;
  LUT5 un1_fracta_i_s0_s_15_RNI757E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[14:14]),.I2(un1_fracta_i_11[14:14]),.I3(un1_fracta_i_10[15:15]),.I4(un1_fracta_i_11[15:15]),.O(m33_2_1));
defparam un1_fracta_i_s0_s_15_RNI757E1_o6.INIT=32'h00110A1B;
  LUT3 un1_fracta_i_s0_s_15_RNI757E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[15:15]),.I2(un1_fracta_i_11[15:15]),.O(N_2605_i));
defparam un1_fracta_i_s0_s_15_RNI757E1_o5.INIT=8'hE4;
  LUT3 un1_fracta_i_s0_s_14_RNID77E1_o6(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[27:27]),.I2(un1_fracta_i_11[27:27]),.O(un1_fracta_i_s0_s_14_RNID77E1_O6));
defparam un1_fracta_i_s0_s_14_RNID77E1_o6.INIT=8'h1B;
  LUT3 un1_fracta_i_s0_s_14_RNID77E1_o5(.I0(fracta_lt_fractb),.I1(un1_fracta_i_10[14:14]),.I2(un1_fracta_i_11[14:14]),.O(N_2604_i));
defparam un1_fracta_i_s0_s_14_RNID77E1_o5.INIT=8'hE4;
  LUT2 fracta_lt_fractb_df26_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[26:26]),.I1(prenorm_addsub_fractb_28_o[26:26]),.O(fracta_lt_fractb_df26));
defparam fracta_lt_fractb_df26_lut6_2_o6.INIT=4'h9;
  LUT2 fracta_lt_fractb_df26_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[26:26]),.I1(prenorm_addsub_fractb_28_o[26:26]),.O(fracta_lt_fractb_lt26));
defparam fracta_lt_fractb_df26_lut6_2_o5.INIT=4'h2;
  LUT4 fracta_lt_fractb_df24_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[24:24]),.I1(prenorm_addsub_fracta_28_o[25:25]),.I2(prenorm_addsub_fractb_28_o[24:24]),.I3(prenorm_addsub_fractb_28_o[25:25]),.O(fracta_lt_fractb_df24));
defparam fracta_lt_fractb_df24_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df24_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[24:24]),.I1(prenorm_addsub_fracta_28_o[25:25]),.I2(prenorm_addsub_fractb_28_o[24:24]),.I3(prenorm_addsub_fractb_28_o[25:25]),.O(fracta_lt_fractb_lt24));
defparam fracta_lt_fractb_df24_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df22_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[22:22]),.I1(prenorm_addsub_fracta_28_o[23:23]),.I2(prenorm_addsub_fractb_28_o[22:22]),.I3(prenorm_addsub_fractb_28_o[23:23]),.O(fracta_lt_fractb_df22));
defparam fracta_lt_fractb_df22_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df22_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[22:22]),.I1(prenorm_addsub_fracta_28_o[23:23]),.I2(prenorm_addsub_fractb_28_o[22:22]),.I3(prenorm_addsub_fractb_28_o[23:23]),.O(fracta_lt_fractb_lt22));
defparam fracta_lt_fractb_df22_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df20_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[20:20]),.I1(prenorm_addsub_fracta_28_o[21:21]),.I2(prenorm_addsub_fractb_28_o[20:20]),.I3(prenorm_addsub_fractb_28_o[21:21]),.O(fracta_lt_fractb_df20));
defparam fracta_lt_fractb_df20_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df20_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[20:20]),.I1(prenorm_addsub_fracta_28_o[21:21]),.I2(prenorm_addsub_fractb_28_o[20:20]),.I3(prenorm_addsub_fractb_28_o[21:21]),.O(fracta_lt_fractb_lt20));
defparam fracta_lt_fractb_df20_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df18_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[18:18]),.I1(prenorm_addsub_fracta_28_o[19:19]),.I2(prenorm_addsub_fractb_28_o[18:18]),.I3(prenorm_addsub_fractb_28_o[19:19]),.O(fracta_lt_fractb_df18));
defparam fracta_lt_fractb_df18_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df18_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[18:18]),.I1(prenorm_addsub_fracta_28_o[19:19]),.I2(prenorm_addsub_fractb_28_o[18:18]),.I3(prenorm_addsub_fractb_28_o[19:19]),.O(fracta_lt_fractb_lt18));
defparam fracta_lt_fractb_df18_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df16_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[16:16]),.I1(prenorm_addsub_fracta_28_o[17:17]),.I2(prenorm_addsub_fractb_28_o[16:16]),.I3(prenorm_addsub_fractb_28_o[17:17]),.O(fracta_lt_fractb_df16));
defparam fracta_lt_fractb_df16_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df16_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[16:16]),.I1(prenorm_addsub_fracta_28_o[17:17]),.I2(prenorm_addsub_fractb_28_o[16:16]),.I3(prenorm_addsub_fractb_28_o[17:17]),.O(fracta_lt_fractb_lt16));
defparam fracta_lt_fractb_df16_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df14_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[14:14]),.I1(prenorm_addsub_fracta_28_o[15:15]),.I2(prenorm_addsub_fractb_28_o[14:14]),.I3(prenorm_addsub_fractb_28_o[15:15]),.O(fracta_lt_fractb_df14));
defparam fracta_lt_fractb_df14_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df14_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[14:14]),.I1(prenorm_addsub_fracta_28_o[15:15]),.I2(prenorm_addsub_fractb_28_o[14:14]),.I3(prenorm_addsub_fractb_28_o[15:15]),.O(fracta_lt_fractb_lt14));
defparam fracta_lt_fractb_df14_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df12_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[12:12]),.I1(prenorm_addsub_fracta_28_o[13:13]),.I2(prenorm_addsub_fractb_28_o[12:12]),.I3(prenorm_addsub_fractb_28_o[13:13]),.O(fracta_lt_fractb_df12));
defparam fracta_lt_fractb_df12_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df12_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[12:12]),.I1(prenorm_addsub_fracta_28_o[13:13]),.I2(prenorm_addsub_fractb_28_o[12:12]),.I3(prenorm_addsub_fractb_28_o[13:13]),.O(fracta_lt_fractb_lt12));
defparam fracta_lt_fractb_df12_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df10_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[10:10]),.I1(prenorm_addsub_fracta_28_o[11:11]),.I2(prenorm_addsub_fractb_28_o[10:10]),.I3(prenorm_addsub_fractb_28_o[11:11]),.O(fracta_lt_fractb_df10));
defparam fracta_lt_fractb_df10_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df10_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[10:10]),.I1(prenorm_addsub_fracta_28_o[11:11]),.I2(prenorm_addsub_fractb_28_o[10:10]),.I3(prenorm_addsub_fractb_28_o[11:11]),.O(fracta_lt_fractb_lt10));
defparam fracta_lt_fractb_df10_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df8_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[8:8]),.I1(prenorm_addsub_fracta_28_o[9:9]),.I2(prenorm_addsub_fractb_28_o[8:8]),.I3(prenorm_addsub_fractb_28_o[9:9]),.O(fracta_lt_fractb_df8));
defparam fracta_lt_fractb_df8_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df8_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[8:8]),.I1(prenorm_addsub_fracta_28_o[9:9]),.I2(prenorm_addsub_fractb_28_o[8:8]),.I3(prenorm_addsub_fractb_28_o[9:9]),.O(fracta_lt_fractb_lt8));
defparam fracta_lt_fractb_df8_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df6_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[6:6]),.I1(prenorm_addsub_fracta_28_o[7:7]),.I2(prenorm_addsub_fractb_28_o[6:6]),.I3(prenorm_addsub_fractb_28_o[7:7]),.O(fracta_lt_fractb_df6));
defparam fracta_lt_fractb_df6_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df6_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[6:6]),.I1(prenorm_addsub_fracta_28_o[7:7]),.I2(prenorm_addsub_fractb_28_o[6:6]),.I3(prenorm_addsub_fractb_28_o[7:7]),.O(fracta_lt_fractb_lt6));
defparam fracta_lt_fractb_df6_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df4_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[4:4]),.I1(prenorm_addsub_fracta_28_o[5:5]),.I2(prenorm_addsub_fractb_28_o[4:4]),.I3(prenorm_addsub_fractb_28_o[5:5]),.O(fracta_lt_fractb_df4));
defparam fracta_lt_fractb_df4_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df4_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[4:4]),.I1(prenorm_addsub_fracta_28_o[5:5]),.I2(prenorm_addsub_fractb_28_o[4:4]),.I3(prenorm_addsub_fractb_28_o[5:5]),.O(fracta_lt_fractb_lt4));
defparam fracta_lt_fractb_df4_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df2_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[2:2]),.I1(prenorm_addsub_fracta_28_o[3:3]),.I2(prenorm_addsub_fractb_28_o[2:2]),.I3(prenorm_addsub_fractb_28_o[3:3]),.O(fracta_lt_fractb_df2));
defparam fracta_lt_fractb_df2_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df2_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[2:2]),.I1(prenorm_addsub_fracta_28_o[3:3]),.I2(prenorm_addsub_fractb_28_o[2:2]),.I3(prenorm_addsub_fractb_28_o[3:3]),.O(fracta_lt_fractb_lt2));
defparam fracta_lt_fractb_df2_lut6_2_o5.INIT=16'h08CE;
  LUT4 fracta_lt_fractb_df0_lut6_2_o6(.I0(prenorm_addsub_fracta_28_o[0:0]),.I1(prenorm_addsub_fracta_28_o[1:1]),.I2(prenorm_addsub_fractb_28_o[0:0]),.I3(prenorm_addsub_fractb_28_o[1:1]),.O(fracta_lt_fractb_df0));
defparam fracta_lt_fractb_df0_lut6_2_o6.INIT=16'h8421;
  LUT4 fracta_lt_fractb_df0_lut6_2_o5(.I0(prenorm_addsub_fracta_28_o[0:0]),.I1(prenorm_addsub_fracta_28_o[1:1]),.I2(prenorm_addsub_fractb_28_o[0:0]),.I3(prenorm_addsub_fractb_28_o[1:1]),.O(fracta_lt_fractb_lt0));
defparam fracta_lt_fractb_df0_lut6_2_o5.INIT=16'h08CE;
endmodule
module post_norm_addsub_inj (addsub_fract_o,v_count_2_0,pre_norm_div_dvsor,s_opa_i,s_output_o_0_0,s_output_o_0_9,postnorm_addsub_output_o,s_output1,s_output_o_1,s_rmode_i,s_fpu_op_i,prenorm_addsub_exp_o,s_opb_i_15,s_opb_i_14,s_opb_i_2,s_opb_i_1,s_opb_i_3,s_opb_i_17,s_opb_i_0,s_opb_i_16,s_opb_i_18,s_opb_i_27,un4_s_infa,un1_s_infb,div_zero_o_0,un3_s_snan_o_0,N_9_i_0_e,N_54,result_2_10,result_i_0_0,s_ine_o,un2_s_qnan_o_0_a2_0_e,N_6_i_0_e,clk_i,N_765_i_0_e,N_763_i_0_e,N_12_i_0_e,N_773_i_0_e,N_1941,un3_s_underflow_o_0,postnorm_addsub_ine_o,result_2_2,N_1055,result_2,result_2_16,N_1051,N_764_i,N_766_i,N_767_i,N_768_i,N_769_i,N_770_i,N_771_i,N_772_i,N_774_i,N_775_i,N_776_i,N_777_i,N_778_i,N_779_i,N_780_i,N_14_i,N_18_i,N_20_i,addsub_sign_o,N_1979,N_36_0,N_1948);
input [27:0] addsub_fract_o ;
input [4:4] v_count_2_0 ;
output [5:5] pre_norm_div_dvsor ;
input [31:31] s_opa_i ;
output s_output_o_0_0 ;
output s_output_o_0_9 ;
output [31:0] postnorm_addsub_output_o ;
input [31:0] s_output1 ;
output s_output_o_1 ;
input [1:0] s_rmode_i ;
input [2:1] s_fpu_op_i ;
input [7:0] prenorm_addsub_exp_o ;
input s_opb_i_15 ;
input s_opb_i_14 ;
input s_opb_i_2 ;
input s_opb_i_1 ;
input s_opb_i_3 ;
input s_opb_i_17 ;
input s_opb_i_0 ;
input s_opb_i_16 ;
input s_opb_i_18 ;
input s_opb_i_27 ;
input un4_s_infa ;
input un1_s_infb ;
input div_zero_o_0 ;
input un3_s_snan_o_0 ;
output N_9_i_0_e ;
input N_54 ;
output result_2_10 ;
output result_i_0_0 ;
input s_ine_o ;
output un2_s_qnan_o_0_a2_0_e ;
output N_6_i_0_e ;
input clk_i ;
output N_765_i_0_e ;
output N_763_i_0_e ;
output N_12_i_0_e ;
output N_773_i_0_e ;
input N_1941 ;
output un3_s_underflow_o_0 ;
output postnorm_addsub_ine_o ;
output result_2_2 ;
input N_1055 ;
output result_2 ;
input result_2_16 ;
input N_1051 ;
output N_764_i ;
output N_766_i ;
output N_767_i ;
output N_768_i ;
output N_769_i ;
output N_770_i ;
output N_771_i ;
output N_772_i ;
output N_774_i ;
output N_775_i ;
output N_776_i ;
output N_777_i ;
output N_778_i ;
output N_779_i ;
output N_780_i ;
output N_14_i ;
output N_18_i ;
output N_20_i ;
input addsub_sign_o ;
input N_1979 ;
input N_36_0 ;
input N_1948 ;
wire s_output_o_0_0 ;
wire s_output_o_0_9 ;
wire s_output_o_1 ;
wire s_opb_i_15 ;
wire s_opb_i_14 ;
wire s_opb_i_2 ;
wire s_opb_i_1 ;
wire s_opb_i_3 ;
wire s_opb_i_17 ;
wire s_opb_i_0 ;
wire s_opb_i_16 ;
wire s_opb_i_18 ;
wire s_opb_i_27 ;
wire un4_s_infa ;
wire un1_s_infb ;
wire div_zero_o_0 ;
wire un3_s_snan_o_0 ;
wire N_9_i_0_e ;
wire N_54 ;
wire result_2_10 ;
wire result_i_0_0 ;
wire s_ine_o ;
wire un2_s_qnan_o_0_a2_0_e ;
wire N_6_i_0_e ;
wire clk_i ;
wire N_765_i_0_e ;
wire N_763_i_0_e ;
wire N_12_i_0_e ;
wire N_773_i_0_e ;
wire N_1941 ;
wire un3_s_underflow_o_0 ;
wire postnorm_addsub_ine_o ;
wire result_2_2 ;
wire N_1055 ;
wire result_2 ;
wire result_2_16 ;
wire N_1051 ;
wire N_764_i ;
wire N_766_i ;
wire N_767_i ;
wire N_768_i ;
wire N_769_i ;
wire N_770_i ;
wire N_771_i ;
wire N_772_i ;
wire N_774_i ;
wire N_775_i ;
wire N_776_i ;
wire N_777_i ;
wire N_778_i ;
wire N_779_i ;
wire N_780_i ;
wire N_14_i ;
wire N_18_i ;
wire N_20_i ;
wire addsub_sign_o ;
wire N_1979 ;
wire N_36_0 ;
wire N_1948 ;
wire [9:0] s_exp10 ;
wire [7:3] s_expo9_3 ;
wire [30:24] s_output_o_0_e ;
wire [25:25] s_output_o_m0 ;
wire s_zeros_0_8 ;
wire s_zeros_0_1 ;
wire s_zeros_0_2 ;
wire [4:0] s_zeros ;
wire [4:4] s_zeros_0_a2_3 ;
wire [1:1] s_zeros_0_i_1_RNI027Q1 ;
wire [4:1] s_exp10_5 ;
wire [4:0] s_shl1 ;
wire [7:0] s_expo9_1_4 ;
wire [7:0] s_expo9_1 ;
wire [27:0] s_fracto28_1 ;
wire [3:3] s_zeros_0_a2_0_2 ;
wire [23:23] s_output_o_1_e ;
wire [5:4] s_expo9_2 ;
wire s_shr1_0_0 ;
wire s_shr1 ;
wire [27:27] s_fracto28_1_3_0 ;
wire [27:3] s_fracto28_rnd ;
wire [16:0] s_fracto28_1_3 ;
wire [22:22] s_output_o ;
wire un1_s_exp10_1 ;
wire [25:3] s_fracto28_2 ;
wire [1:1] s_zeros_0_i_a2_2 ;
wire [1:1] s_zeros_0_i_1 ;
wire [3:0] s_zeros_0_0 ;
wire s_zeros_0_8_tz ;
wire s_zeros_0_4 ;
wire [7:5] s_exp10_5_i ;
wire GND ;
wire s_exp10_s_9_true ;
wire un11_s_exp10_7_3 ;
wire un1_s_exp10_3_i ;
wire un15_s_zero_fract_sn ;
wire s_overflow ;
wire VCC ;
wire N_473_i ;
wire N_2203 ;
wire N_84 ;
wire N_311 ;
wire N_388 ;
wire N_329 ;
wire N_345 ;
wire un1_s_exp10_3 ;
wire N_389 ;
wire N_1832 ;
wire N_1803 ;
wire N_1815 ;
wire N_68 ;
wire N_1833 ;
wire N_1816 ;
wire N_1821 ;
wire N_1822 ;
wire N_1807 ;
wire N_1808 ;
wire N_1823 ;
wire N_1809 ;
wire N_91 ;
wire N_835 ;
wire N_92 ;
wire s_exp10_5_c4 ;
wire s_exp10_5_c3 ;
wire N_1697 ;
wire N_1696 ;
wire N_1686 ;
wire N_1727 ;
wire N_1726 ;
wire N_1720 ;
wire N_1684 ;
wire N_1685 ;
wire N_1812 ;
wire N_1725_i ;
wire N_1683 ;
wire N_1729 ;
wire N_1693 ;
wire N_331 ;
wire N_1776 ;
wire N_58 ;
wire s_exp10_5_c2 ;
wire result_1 ;
wire N_1861 ;
wire m149_0 ;
wire N_289 ;
wire N_1709 ;
wire N_1869 ;
wire N_6 ;
wire N_844_0_4 ;
wire N_91_0_0_1 ;
wire m149_e_1 ;
wire N_1705 ;
wire N_8 ;
wire N_1700 ;
wire N_1855 ;
wire N_1712 ;
wire N_1842 ;
wire N_1711 ;
wire N_1774 ;
wire N_1713 ;
wire N_1708 ;
wire N_1676 ;
wire N_1707 ;
wire N_1701 ;
wire N_299_2 ;
wire N_1706 ;
wire un6_s_expo9_3_c4 ;
wire un6_s_expo9_3_c6 ;
wire un2_s_expo9_2 ;
wire N_811_4 ;
wire N_811_1 ;
wire N_1872 ;
wire un1_s_expo9_3 ;
wire N_82 ;
wire N_836 ;
wire N_811_0_4 ;
wire N_1800 ;
wire N_1857 ;
wire un2_s_ine_o_i_a5_1 ;
wire N_2179_i_0 ;
wire un3_s_fracto28_rnd_1_axb_1 ;
wire un3_s_fracto28_rnd_1_axb_2 ;
wire un3_s_fracto28_rnd_1_axb_3 ;
wire un3_s_fracto28_rnd_1_axb_4 ;
wire un3_s_fracto28_rnd_1_axb_5 ;
wire un3_s_fracto28_rnd_1_axb_6 ;
wire un3_s_fracto28_rnd_1_axb_7 ;
wire un3_s_fracto28_rnd_1_axb_8 ;
wire un3_s_fracto28_rnd_1_axb_9 ;
wire un3_s_fracto28_rnd_1_axb_10 ;
wire un3_s_fracto28_rnd_1_axb_11 ;
wire un3_s_fracto28_rnd_1_axb_12 ;
wire un3_s_fracto28_rnd_1_axb_13 ;
wire un3_s_fracto28_rnd_1_axb_14 ;
wire un3_s_fracto28_rnd_1_axb_15 ;
wire un3_s_fracto28_rnd_1_axb_16 ;
wire un3_s_fracto28_rnd_1_axb_17 ;
wire un3_s_fracto28_rnd_1_axb_18 ;
wire un3_s_fracto28_rnd_1_axb_19 ;
wire un3_s_fracto28_rnd_1_axb_20 ;
wire un3_s_fracto28_rnd_1_axb_21 ;
wire un3_s_fracto28_rnd_1_axb_22 ;
wire un3_s_fracto28_rnd_1_axb_23 ;
wire N_1806_i ;
wire N_1811_i ;
wire N_1814_i ;
wire N_1818_i ;
wire N_1820_i ;
wire N_1825_i ;
wire N_1831_i ;
wire N_1835_i ;
wire N_1841_i ;
wire N_1848_i ;
wire N_1854_i ;
wire N_1779_i ;
wire N_1781_i ;
wire N_1784_i ;
wire N_1787_i ;
wire N_1790_i ;
wire N_28_0_i ;
wire N_1795_i ;
wire N_1796_i ;
wire N_1799_i ;
wire N_1802_i ;
wire N_3392_mux ;
wire N_390 ;
wire N_391 ;
wire N_392 ;
wire un12_s_exp10_iso ;
wire s_overflow_1 ;
wire s_expo9_0_c4 ;
wire N_1770 ;
wire s_exp10_axb_1 ;
wire N_60 ;
wire N_1723 ;
wire s_roundup_1_3_i_a2_0 ;
wire N_85 ;
wire un3_s_fracto28_rnd_1_s_1 ;
wire un3_s_fracto28_rnd_1_s_24 ;
wire N_4 ;
wire s_exp10_5_axb0 ;
wire un3_s_fracto28_rnd_1_axb_24 ;
wire N_835_1_4 ;
wire N_835_3_4 ;
wire N_338 ;
wire N_835_0 ;
wire N_835_2 ;
wire N_1692 ;
wire N_1695 ;
wire N_1721 ;
wire N_1722 ;
wire N_1827 ;
wire N_1837 ;
wire N_1850 ;
wire N_1673 ;
wire N_61 ;
wire N_1844 ;
wire N_62 ;
wire N_64 ;
wire N_337 ;
wire N_1877 ;
wire N_63 ;
wire N_1769 ;
wire N_1797 ;
wire N_1829 ;
wire N_105 ;
wire N_1852 ;
wire N_1839 ;
wire un12_s_exp10 ;
wire N_93 ;
wire un3_s_fracto28_rnd_1_s_23 ;
wire un3_s_fracto28_rnd_1_s_22 ;
wire un3_s_fracto28_rnd_1_s_2 ;
wire un3_s_fracto28_rnd_1_s_3 ;
wire un3_s_fracto28_rnd_1_s_4 ;
wire un3_s_fracto28_rnd_1_s_5 ;
wire un3_s_fracto28_rnd_1_s_6 ;
wire un3_s_fracto28_rnd_1_s_7 ;
wire un3_s_fracto28_rnd_1_s_8 ;
wire un3_s_fracto28_rnd_1_s_9 ;
wire un3_s_fracto28_rnd_1_s_10 ;
wire un3_s_fracto28_rnd_1_s_11 ;
wire un3_s_fracto28_rnd_1_s_12 ;
wire un3_s_fracto28_rnd_1_s_13 ;
wire un3_s_fracto28_rnd_1_s_14 ;
wire un3_s_fracto28_rnd_1_s_15 ;
wire un3_s_fracto28_rnd_1_s_19 ;
wire un3_s_fracto28_rnd_1_s_20 ;
wire un3_s_fracto28_rnd_1_s_21 ;
wire un3_s_fracto28_rnd_1_s_18 ;
wire un3_s_fracto28_rnd_1_s_17 ;
wire un3_s_fracto28_rnd_1_s_16 ;
wire N_1847 ;
wire s_exp10_5_ac0_13_i ;
wire s_overflow_0_0 ;
wire s_overflow_2 ;
wire s_exp10_axb_2 ;
wire s_exp10_axb_3 ;
wire s_exp10_axb_4 ;
wire un3_s_fracto28_rnd_1_cry_23 ;
wire un3_s_fracto28_rnd_1_cry_22 ;
wire un3_s_fracto28_rnd_1_cry_21 ;
wire un3_s_fracto28_rnd_1_cry_20 ;
wire un3_s_fracto28_rnd_1_cry_19 ;
wire un3_s_fracto28_rnd_1_cry_18 ;
wire un3_s_fracto28_rnd_1_cry_17 ;
wire un3_s_fracto28_rnd_1_cry_16 ;
wire un3_s_fracto28_rnd_1_cry_15 ;
wire un3_s_fracto28_rnd_1_cry_14 ;
wire un3_s_fracto28_rnd_1_cry_13 ;
wire un3_s_fracto28_rnd_1_cry_12 ;
wire un3_s_fracto28_rnd_1_cry_11 ;
wire un3_s_fracto28_rnd_1_cry_10 ;
wire un3_s_fracto28_rnd_1_cry_9 ;
wire un3_s_fracto28_rnd_1_cry_8 ;
wire un3_s_fracto28_rnd_1_cry_7 ;
wire un3_s_fracto28_rnd_1_cry_6 ;
wire un3_s_fracto28_rnd_1_cry_5 ;
wire un3_s_fracto28_rnd_1_cry_4 ;
wire un3_s_fracto28_rnd_1_cry_3 ;
wire un3_s_fracto28_rnd_1_cry_2 ;
wire un3_s_fracto28_rnd_1_cry_1 ;
wire s_exp10_cry_8 ;
wire s_exp10_cry_7 ;
wire s_exp10_cry_6 ;
wire s_exp10_cry_5 ;
wire s_exp10_cry_4 ;
wire s_exp10_cry_3 ;
wire s_exp10_cry_2 ;
wire s_exp10_cry_1 ;
wire s_exp10_cry_0 ;
// instances
  LUT1 s_exp10_s_9_true_cZ(.I0(GND),.O(s_exp10_s_9_true));
defparam s_exp10_s_9_true_cZ.INIT=2'h3;
  LUT5 un1_s_exp10_3_i_cZ(.I0(s_exp10[3:3]),.I1(s_exp10[4:4]),.I2(s_exp10[7:7]),.I3(s_exp10[8:8]),.I4(un11_s_exp10_7_3),.O(un1_s_exp10_3_i));
defparam un1_s_exp10_3_i_cZ.INIT=32'hFF01FF00;
  LUT6_2 desc303(.I0(prenorm_addsub_exp_o[0:0]),.I1(s_zeros_0_8),.I2(s_zeros_0_1),.I3(N_311),.I4(s_zeros_0_2),.I5(un1_s_exp10_3_i),.O6(N_388),.O5(s_zeros[0:0]));
defparam desc303.INIT=64'h55555555FFFFFFFC;
  LUT6_2 desc304(.I0(addsub_fract_o[12:12]),.I1(addsub_fract_o[20:20]),.I2(addsub_fract_o[16:16]),.I3(addsub_fract_o[18:18]),.I4(N_329),.I5(s_zeros_0_a2_3[4:4]),.O6(s_zeros[4:4]),.O5(N_345));
defparam desc304.INIT=64'h0000000000010000;
  LUT6_2 desc305(.I0(s_shl1[1:1]),.I1(N_1720),.I2(N_1696),.I3(N_1684),.I4(N_1685),.I5(s_shl1[3:3]),.O6(N_1812),.O5(N_1725_i));
defparam desc305.INIT=64'h05AF05AF1111BBBB;
  LUT6_2 desc306(.I0(s_shl1[1:1]),.I1(N_1683),.I2(N_1686),.I3(N_1684),.I4(N_1685),.I5(s_shl1[3:3]),.O6(N_1729),.O5(N_1693));
defparam desc306.INIT=64'hDD88DD88F5F5A0A0;
  FD desc307(.Q(postnorm_addsub_output_o[30:30]),.D(s_output_o_0_e[30:30]),.C(clk_i));
  FD desc308(.Q(postnorm_addsub_output_o[29:29]),.D(s_output_o_0_e[29:29]),.C(clk_i));
  FD desc309(.Q(postnorm_addsub_output_o[28:28]),.D(s_output_o_0_e[28:28]),.C(clk_i));
  FD desc310(.Q(postnorm_addsub_output_o[27:27]),.D(s_output_o_0_e[27:27]),.C(clk_i));
  FD desc311(.Q(postnorm_addsub_output_o[26:26]),.D(s_output_o_0_e[26:26]),.C(clk_i));
  FD desc312(.Q(postnorm_addsub_output_o[25:25]),.D(s_output_o_0_e[25:25]),.C(clk_i));
  FD desc313(.Q(postnorm_addsub_output_o[24:24]),.D(s_output_o_0_e[24:24]),.C(clk_i));
  FD desc314(.Q(postnorm_addsub_output_o[23:23]),.D(s_output_o_1_e[23:23]),.C(clk_i));
  LUT6 desc315(.I0(N_2203),.I1(s_expo9_2[4:4]),.I2(s_expo9_2[5:5]),.I3(un1_s_expo9_3),.I4(un6_s_expo9_3_c4),.I5(un15_s_zero_fract_sn),.O(s_output_o_0_e[28:28]));
defparam desc315.INIT=64'h555555557DF5F5F5;
  LUT6 desc316(.I0(N_2203),.I1(s_expo9_1[0:0]),.I2(s_expo9_1[1:1]),.I3(un1_s_expo9_3),.I4(un2_s_expo9_2),.I5(un15_s_zero_fract_sn),.O(s_output_o_0_e[24:24]));
defparam desc316.INIT=64'h55555555F5D77DF5;
  LUT5 desc317(.I0(N_2203),.I1(s_expo9_2[4:4]),.I2(un1_s_expo9_3),.I3(un6_s_expo9_3_c4),.I4(un15_s_zero_fract_sn),.O(s_output_o_0_e[27:27]));
defparam desc317.INIT=32'h55557DDD;
  LUT6 desc318(.I0(N_2203),.I1(s_expo9_1[0:0]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(un1_s_expo9_3),.I5(un15_s_zero_fract_sn),.O(s_output_o_1_e[23:23]));
defparam desc318.INIT=64'h55555555777DDDD7;
  LUT6 un2_s_inf_o_i_a2_RNI66FI1(.I0(N_82),.I1(N_84),.I2(N_92),.I3(s_output1[6:6]),.I4(s_rmode_i[0:0]),.I5(N_836),.O(N_765_i_0_e));
defparam un2_s_inf_o_i_a2_RNI66FI1.INIT=64'h00000000FF02FF01;
  LUT6 un2_s_inf_o_i_a2_RNI22FI1(.I0(N_82),.I1(N_84),.I2(N_92),.I3(s_output1[2:2]),.I4(s_rmode_i[0:0]),.I5(N_836),.O(N_763_i_0_e));
defparam un2_s_inf_o_i_a2_RNI22FI1.INIT=64'h00000000FF02FF01;
  LUT6 un2_s_inf_o_i_a2_RNI00FI1(.I0(N_82),.I1(N_84),.I2(N_92),.I3(s_output1[0:0]),.I4(s_rmode_i[0:0]),.I5(N_836),.O(N_12_i_0_e));
defparam un2_s_inf_o_i_a2_RNI00FI1.INIT=64'h00000000FF02FF01;
  LUT6 un2_s_inf_o_i_a2_RNILM7S1(.I0(N_82),.I1(N_84),.I2(N_92),.I3(s_output1[14:14]),.I4(s_rmode_i[0:0]),.I5(N_836),.O(N_773_i_0_e));
defparam un2_s_inf_o_i_a2_RNILM7S1.INIT=64'h00000000FF02FF01;
  LUT5 desc319(.I0(s_expo9_3[7:7]),.I1(s_overflow),.I2(un15_s_zero_fract_sn),.I3(un1_s_infb),.I4(un4_s_infa),.O(s_output_o_0_e[30:30]));
defparam desc319.INIT=32'hFFFFFFCE;
  LUT6 desc320(.I0(N_82),.I1(N_84),.I2(N_91),.I3(s_output1[22:22]),.I4(s_output1[23:23]),.I5(s_rmode_i[0:0]),.O(s_output_o_0_0));
defparam desc320.INIT=64'hFF02FF00FF01FF00;
  LUT6 desc321(.I0(N_811_0_4),.I1(N_811_1),.I2(N_1941),.I3(s_fpu_op_i[2:2]),.I4(s_opa_i[31:31]),.I5(s_output1[31:31]),.O(s_output_o_0_9));
defparam desc321.INIT=64'hFFFFFFFF00880008;
  LUT6 un3_s_underflow_o_0_a2_0_0_4_lut6_2_RNI6FO72(.I0(N_844_0_4),.I1(s_ine_o),.I2(s_output1[24:24]),.I3(s_output1[25:25]),.I4(s_output1[26:26]),.I5(s_output1[30:30]),.O(un3_s_underflow_o_0));
defparam un3_s_underflow_o_0_a2_0_0_4_lut6_2_RNI6FO72.INIT=64'h0000000000000008;
  LUT6 desc322(.I0(addsub_fract_o[27:27]),.I1(s_exp10[3:3]),.I2(s_exp10[4:4]),.I3(s_exp10[7:7]),.I4(s_exp10[8:8]),.I5(un11_s_exp10_7_3),.O(s_shr1_0_0));
defparam desc322.INIT=64'h0000AAA80000AAAA;
  LUT6 desc323(.I0(N_1800),.I1(N_1815),.I2(N_1857),.I3(s_shl1[3:3]),.I4(s_shl1[4:4]),.I5(s_shr1),.O(s_fracto28_1_3_0[27:27]));
defparam desc323.INIT=64'h000000005555330F;
  LUT6 ine_o_RNO(.I0(s_fracto28_rnd[3:3]),.I1(s_fracto28_rnd[27:27]),.I2(s_overflow),.I3(un2_s_ine_o_i_a5_1),.I4(un1_s_infb),.I5(un4_s_infa),.O(N_2179_i_0));
defparam ine_o_RNO.INIT=64'h000000000000F8FF;
  LUT1 un3_s_fracto28_rnd_1_axb_1_cZ(.I0(s_fracto28_1[4:4]),.O(un3_s_fracto28_rnd_1_axb_1));
defparam un3_s_fracto28_rnd_1_axb_1_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_2_cZ(.I0(s_fracto28_1[5:5]),.O(un3_s_fracto28_rnd_1_axb_2));
defparam un3_s_fracto28_rnd_1_axb_2_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_3_cZ(.I0(s_fracto28_1[6:6]),.O(un3_s_fracto28_rnd_1_axb_3));
defparam un3_s_fracto28_rnd_1_axb_3_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_4_cZ(.I0(s_fracto28_1[7:7]),.O(un3_s_fracto28_rnd_1_axb_4));
defparam un3_s_fracto28_rnd_1_axb_4_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_5_cZ(.I0(s_fracto28_1[8:8]),.O(un3_s_fracto28_rnd_1_axb_5));
defparam un3_s_fracto28_rnd_1_axb_5_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_6_cZ(.I0(s_fracto28_1[9:9]),.O(un3_s_fracto28_rnd_1_axb_6));
defparam un3_s_fracto28_rnd_1_axb_6_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_7_cZ(.I0(s_fracto28_1[10:10]),.O(un3_s_fracto28_rnd_1_axb_7));
defparam un3_s_fracto28_rnd_1_axb_7_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_8_cZ(.I0(s_fracto28_1[11:11]),.O(un3_s_fracto28_rnd_1_axb_8));
defparam un3_s_fracto28_rnd_1_axb_8_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_9_cZ(.I0(s_fracto28_1[12:12]),.O(un3_s_fracto28_rnd_1_axb_9));
defparam un3_s_fracto28_rnd_1_axb_9_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_10_cZ(.I0(s_fracto28_1[13:13]),.O(un3_s_fracto28_rnd_1_axb_10));
defparam un3_s_fracto28_rnd_1_axb_10_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_11_cZ(.I0(s_fracto28_1[14:14]),.O(un3_s_fracto28_rnd_1_axb_11));
defparam un3_s_fracto28_rnd_1_axb_11_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_12_cZ(.I0(s_fracto28_1[15:15]),.O(un3_s_fracto28_rnd_1_axb_12));
defparam un3_s_fracto28_rnd_1_axb_12_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_13_cZ(.I0(s_fracto28_1[16:16]),.O(un3_s_fracto28_rnd_1_axb_13));
defparam un3_s_fracto28_rnd_1_axb_13_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_14_cZ(.I0(s_fracto28_1[17:17]),.O(un3_s_fracto28_rnd_1_axb_14));
defparam un3_s_fracto28_rnd_1_axb_14_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_15_cZ(.I0(s_fracto28_1[18:18]),.O(un3_s_fracto28_rnd_1_axb_15));
defparam un3_s_fracto28_rnd_1_axb_15_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_16_cZ(.I0(s_fracto28_1[19:19]),.O(un3_s_fracto28_rnd_1_axb_16));
defparam un3_s_fracto28_rnd_1_axb_16_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_17_cZ(.I0(s_fracto28_1[20:20]),.O(un3_s_fracto28_rnd_1_axb_17));
defparam un3_s_fracto28_rnd_1_axb_17_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_18_cZ(.I0(s_fracto28_1[21:21]),.O(un3_s_fracto28_rnd_1_axb_18));
defparam un3_s_fracto28_rnd_1_axb_18_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_19_cZ(.I0(s_fracto28_1[22:22]),.O(un3_s_fracto28_rnd_1_axb_19));
defparam un3_s_fracto28_rnd_1_axb_19_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_20_cZ(.I0(s_fracto28_1[23:23]),.O(un3_s_fracto28_rnd_1_axb_20));
defparam un3_s_fracto28_rnd_1_axb_20_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_21_cZ(.I0(s_fracto28_1[24:24]),.O(un3_s_fracto28_rnd_1_axb_21));
defparam un3_s_fracto28_rnd_1_axb_21_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_22_cZ(.I0(s_fracto28_1[25:25]),.O(un3_s_fracto28_rnd_1_axb_22));
defparam un3_s_fracto28_rnd_1_axb_22_cZ.INIT=2'h2;
  LUT1 un3_s_fracto28_rnd_1_axb_23_cZ(.I0(s_fracto28_1[26:26]),.O(un3_s_fracto28_rnd_1_axb_23));
defparam un3_s_fracto28_rnd_1_axb_23_cZ.INIT=2'h2;
  FD desc324(.Q(s_fracto28_1[27:27]),.D(s_fracto28_1_3_0[27:27]),.C(clk_i));
  FD desc325(.Q(s_fracto28_1[12:12]),.D(s_fracto28_1_3[12:12]),.C(clk_i));
  FD desc326(.Q(s_fracto28_1[13:13]),.D(s_fracto28_1_3[13:13]),.C(clk_i));
  FD desc327(.Q(s_fracto28_1[14:14]),.D(s_fracto28_1_3[14:14]),.C(clk_i));
  FD desc328(.Q(s_fracto28_1[15:15]),.D(N_1806_i),.C(clk_i));
  FD desc329(.Q(s_fracto28_1[16:16]),.D(s_fracto28_1_3[16:16]),.C(clk_i));
  FD desc330(.Q(s_fracto28_1[17:17]),.D(N_1811_i),.C(clk_i));
  FD desc331(.Q(s_fracto28_1[18:18]),.D(N_1814_i),.C(clk_i));
  FD desc332(.Q(s_fracto28_1[19:19]),.D(N_1818_i),.C(clk_i));
  FD desc333(.Q(s_fracto28_1[20:20]),.D(N_1820_i),.C(clk_i));
  FD desc334(.Q(s_fracto28_1[21:21]),.D(N_1825_i),.C(clk_i));
  FD desc335(.Q(s_fracto28_1[22:22]),.D(N_1831_i),.C(clk_i));
  FD desc336(.Q(s_fracto28_1[23:23]),.D(N_1835_i),.C(clk_i));
  FD desc337(.Q(s_fracto28_1[24:24]),.D(N_1841_i),.C(clk_i));
  FD desc338(.Q(s_fracto28_1[25:25]),.D(N_1848_i),.C(clk_i));
  FD desc339(.Q(s_fracto28_1[26:26]),.D(N_1854_i),.C(clk_i));
  FD desc340(.Q(s_fracto28_1[0:0]),.D(s_fracto28_1_3[0:0]),.C(clk_i));
  FD desc341(.Q(s_fracto28_1[1:1]),.D(N_1779_i),.C(clk_i));
  FD desc342(.Q(s_fracto28_1[2:2]),.D(N_1781_i),.C(clk_i));
  FD desc343(.Q(s_fracto28_1[3:3]),.D(N_1784_i),.C(clk_i));
  FD desc344(.Q(s_fracto28_1[4:4]),.D(N_1787_i),.C(clk_i));
  FD desc345(.Q(s_fracto28_1[5:5]),.D(N_1790_i),.C(clk_i));
  FD desc346(.Q(s_fracto28_1[6:6]),.D(N_28_0_i),.C(clk_i));
  FD desc347(.Q(s_fracto28_1[7:7]),.D(N_1795_i),.C(clk_i));
  FD desc348(.Q(s_fracto28_1[8:8]),.D(N_1796_i),.C(clk_i));
  FD desc349(.Q(s_fracto28_1[9:9]),.D(s_fracto28_1_3[9:9]),.C(clk_i));
  FD desc350(.Q(s_fracto28_1[10:10]),.D(N_1799_i),.C(clk_i));
  FD desc351(.Q(s_fracto28_1[11:11]),.D(N_1802_i),.C(clk_i));
  FD desc352(.Q(postnorm_addsub_output_o[31:31]),.D(N_3392_mux),.C(clk_i));
  FD desc353(.Q(postnorm_addsub_output_o[22:22]),.D(s_output_o[22:22]),.C(clk_i));
  FD ine_o_Z(.Q(postnorm_addsub_ine_o),.D(N_2179_i_0),.C(clk_i));
  FDR desc354(.Q(s_shl1[0:0]),.D(N_388),.C(clk_i),.R(un1_s_exp10_1));
  FDR desc355(.Q(s_shl1[1:1]),.D(N_389),.C(clk_i),.R(un1_s_exp10_1));
  FDR desc356(.Q(s_shl1[2:2]),.D(N_390),.C(clk_i),.R(un1_s_exp10_1));
  FDR desc357(.Q(s_shl1[3:3]),.D(N_391),.C(clk_i),.R(un1_s_exp10_1));
  FDR desc358(.Q(s_shl1[4:4]),.D(N_392),.C(clk_i),.R(un1_s_exp10_1));
  FDR desc359(.Q(postnorm_addsub_output_o[16:16]),.D(s_fracto28_2[19:19]),.C(clk_i),.R(N_473_i));
  FDR desc360(.Q(postnorm_addsub_output_o[17:17]),.D(s_fracto28_2[20:20]),.C(clk_i),.R(N_473_i));
  FDR desc361(.Q(postnorm_addsub_output_o[18:18]),.D(s_fracto28_2[21:21]),.C(clk_i),.R(N_473_i));
  FDR desc362(.Q(postnorm_addsub_output_o[19:19]),.D(s_fracto28_2[22:22]),.C(clk_i),.R(N_473_i));
  FDR desc363(.Q(postnorm_addsub_output_o[20:20]),.D(s_fracto28_2[23:23]),.C(clk_i),.R(N_473_i));
  FDR desc364(.Q(postnorm_addsub_output_o[21:21]),.D(s_fracto28_2[24:24]),.C(clk_i),.R(N_473_i));
  FDR desc365(.Q(postnorm_addsub_output_o[1:1]),.D(s_fracto28_2[4:4]),.C(clk_i),.R(N_473_i));
  FDR desc366(.Q(postnorm_addsub_output_o[2:2]),.D(s_fracto28_2[5:5]),.C(clk_i),.R(N_473_i));
  FDR desc367(.Q(postnorm_addsub_output_o[3:3]),.D(s_fracto28_2[6:6]),.C(clk_i),.R(N_473_i));
  FDR desc368(.Q(postnorm_addsub_output_o[4:4]),.D(s_fracto28_2[7:7]),.C(clk_i),.R(N_473_i));
  FDR desc369(.Q(postnorm_addsub_output_o[5:5]),.D(s_fracto28_2[8:8]),.C(clk_i),.R(N_473_i));
  FDR desc370(.Q(postnorm_addsub_output_o[6:6]),.D(s_fracto28_2[9:9]),.C(clk_i),.R(N_473_i));
  FDR desc371(.Q(postnorm_addsub_output_o[7:7]),.D(s_fracto28_2[10:10]),.C(clk_i),.R(N_473_i));
  FDR desc372(.Q(postnorm_addsub_output_o[8:8]),.D(s_fracto28_2[11:11]),.C(clk_i),.R(N_473_i));
  FDR desc373(.Q(postnorm_addsub_output_o[9:9]),.D(s_fracto28_2[12:12]),.C(clk_i),.R(N_473_i));
  FDR desc374(.Q(postnorm_addsub_output_o[10:10]),.D(s_fracto28_2[13:13]),.C(clk_i),.R(N_473_i));
  FDR desc375(.Q(postnorm_addsub_output_o[11:11]),.D(s_fracto28_2[14:14]),.C(clk_i),.R(N_473_i));
  FDR desc376(.Q(postnorm_addsub_output_o[12:12]),.D(s_fracto28_2[15:15]),.C(clk_i),.R(N_473_i));
  FDR desc377(.Q(postnorm_addsub_output_o[13:13]),.D(s_fracto28_2[16:16]),.C(clk_i),.R(N_473_i));
  FDR desc378(.Q(postnorm_addsub_output_o[14:14]),.D(s_fracto28_2[17:17]),.C(clk_i),.R(N_473_i));
  FDR desc379(.Q(postnorm_addsub_output_o[15:15]),.D(s_fracto28_2[18:18]),.C(clk_i),.R(N_473_i));
  FDR desc380(.Q(postnorm_addsub_output_o[0:0]),.D(s_fracto28_2[3:3]),.C(clk_i),.R(N_473_i));
  LUT6 un12_s_exp10_iso_cZ(.I0(s_exp10[3:3]),.I1(s_exp10[4:4]),.I2(s_exp10[9:9]),.I3(s_exp10[7:7]),.I4(s_exp10[8:8]),.I5(un11_s_exp10_7_3),.O(un12_s_exp10_iso));
defparam un12_s_exp10_iso_cZ.INIT=64'hF0F0F0F1F0F0F0F0;
  LUT6 s_overflow_1_cZ(.I0(s_expo9_1[2:2]),.I1(s_expo9_1[1:1]),.I2(s_expo9_1[0:0]),.I3(s_fracto28_1[26:26]),.I4(s_fracto28_1[27:27]),.I5(un1_s_expo9_3),.O(s_overflow_1));
defparam s_overflow_1_cZ.INIT=64'h2828288888888881;
  LUT6 un1_s_expo9_3_cZ(.I0(s_expo9_1[6:6]),.I1(s_expo9_1[7:7]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(un6_s_expo9_3_c6),.I5(s_fracto28_rnd[27:27]),.O(un1_s_expo9_3));
defparam un1_s_expo9_3_cZ.INIT=64'h777EFFFF00000000;
  LUT6 desc381(.I0(s_expo9_1[6:6]),.I1(s_expo9_1[7:7]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(un6_s_expo9_3_c6),.I5(s_fracto28_rnd[27:27]),.O(s_expo9_3[7:7]));
defparam desc381.INIT=64'hEEEDCCCCCCC9CCCC;
  LUT6 desc382(.I0(s_expo9_1[6:6]),.I1(s_expo9_1[7:7]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(un6_s_expo9_3_c6),.I5(s_fracto28_rnd[27:27]),.O(s_expo9_3[6:6]));
defparam desc382.INIT=64'hDDDBAAAAAAA5AAAA;
  LUT5 desc383(.I0(s_expo9_1[5:5]),.I1(s_expo9_1[4:4]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(s_expo9_0_c4),.O(s_expo9_2[5:5]));
defparam desc383.INIT=32'hAAAAAAA9;
  LUT5 desc384(.I0(addsub_fract_o[17:17]),.I1(addsub_fract_o[18:18]),.I2(s_zeros_0_i_a2_2[1:1]),.I3(s_zeros_0_i_1[1:1]),.I4(N_1770),.O(s_zeros_0_i_1_RNI027Q1[1:1]));
defparam desc384.INIT=32'hFFF0FFE0;
  LUT6 s_exp10_5_axbxc1_lut6_2_RNIVR242(.I0(addsub_fract_o[17:17]),.I1(addsub_fract_o[18:18]),.I2(s_exp10_5[1:1]),.I3(s_zeros_0_i_a2_2[1:1]),.I4(s_zeros_0_i_1[1:1]),.I5(N_1770),.O(s_exp10_axb_1));
defparam s_exp10_5_axbxc1_lut6_2_RNIVR242.INIT=64'h0F0F0FF00F0F1EF0;
  LUT5 desc385(.I0(s_opb_i_2),.I1(s_opb_i_1),.I2(s_opb_i_3),.I3(result_2_2),.I4(N_1055),.O(result_2));
defparam desc385.INIT=32'hFFFEFFFF;
  LUT6 desc386(.I0(prenorm_addsub_exp_o[0:0]),.I1(addsub_fract_o[27:27]),.I2(s_zeros_0_8),.I3(s_zeros_0_1),.I4(N_311),.I5(s_zeros_0_2),.O(s_exp10[0:0]));
defparam desc386.INIT=64'h9999999999999996;
  LUT6 desc387(.I0(addsub_fract_o[2:2]),.I1(addsub_fract_o[3:3]),.I2(s_shl1[2:2]),.I3(s_shl1[1:1]),.I4(s_shl1[0:0]),.I5(N_1711),.O(N_60));
defparam desc387.INIT=64'h0F0A0F0C000A000C;
  LUT6 desc388(.I0(s_opb_i_17),.I1(s_opb_i_0),.I2(s_opb_i_16),.I3(s_opb_i_18),.I4(result_2_16),.I5(N_1051),.O(result_2_2));
defparam desc388.INIT=64'hFFFFFFFEFFFFFFFF;
  LUT5 s_exp10_cry_3_RNO(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[3:3]),.I2(prenorm_addsub_exp_o[0:0]),.I3(prenorm_addsub_exp_o[2:2]),.I4(addsub_fract_o[27:27]),.O(s_exp10_5[3:3]));
defparam s_exp10_cry_3_RNO.INIT=32'h66CC6CCC;
  LUT4 s_exp10_cry_2_RNO(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.I2(prenorm_addsub_exp_o[2:2]),.I3(addsub_fract_o[27:27]),.O(s_exp10_5[2:2]));
defparam s_exp10_cry_2_RNO.INIT=16'h5A78;
  LUT6_L desc389(.I0(addsub_fract_o[1:1]),.I1(addsub_fract_o[2:2]),.I2(addsub_fract_o[4:4]),.I3(addsub_fract_o[3:3]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.LO(N_1723));
defparam desc389.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc390(.I0(addsub_fract_o[4:4]),.I1(addsub_fract_o[7:7]),.I2(addsub_fract_o[3:3]),.I3(addsub_fract_o[8:8]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1684));
defparam desc390.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6_L desc391(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(s_shl1[3:3]),.I3(N_1711),.I4(N_1712),.I5(N_68),.LO(N_1800));
defparam desc391.INIT=64'hA0E0B0F0AFEFBFFF;
  LUT6 s_exp10_cry_4_RNO(.I0(prenorm_addsub_exp_o[4:4]),.I1(prenorm_addsub_exp_o[1:1]),.I2(prenorm_addsub_exp_o[3:3]),.I3(prenorm_addsub_exp_o[0:0]),.I4(prenorm_addsub_exp_o[2:2]),.I5(addsub_fract_o[27:27]),.O(s_exp10_5[4:4]));
defparam s_exp10_cry_4_RNO.INIT=64'h6A6AAAAA6AAAAAAA;
  LUT4 s_roundup_1_3_i_a2_0_0(.I0(s_fracto28_1[0:0]),.I1(s_fracto28_1[1:1]),.I2(addsub_fract_o[0:0]),.I3(addsub_fract_o[27:27]),.O(s_roundup_1_3_i_a2_0));
defparam s_roundup_1_3_i_a2_0_0.INIT=16'h0111;
  LUT5 un2_s_ine_o_i_a5_1_cZ(.I0(s_fracto28_1[0:0]),.I1(s_fracto28_1[1:1]),.I2(s_fracto28_1[2:2]),.I3(addsub_fract_o[0:0]),.I4(s_shr1),.O(un2_s_ine_o_i_a5_1));
defparam un2_s_ine_o_i_a5_1_cZ.INIT=32'h00010101;
  LUT6_L desc392(.I0(s_output1[5:5]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_764_i));
defparam desc392.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc393(.I0(s_output1[7:7]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_766_i));
defparam desc393.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc394(.I0(s_output1[8:8]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_767_i));
defparam desc394.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc395(.I0(s_output1[9:9]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_768_i));
defparam desc395.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc396(.I0(s_output1[10:10]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_769_i));
defparam desc396.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc397(.I0(s_output1[11:11]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_770_i));
defparam desc397.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc398(.I0(s_output1[12:12]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_771_i));
defparam desc398.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc399(.I0(s_output1[13:13]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_772_i));
defparam desc399.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc400(.I0(s_output1[15:15]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_774_i));
defparam desc400.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc401(.I0(s_output1[16:16]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_775_i));
defparam desc401.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc402(.I0(s_output1[17:17]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_776_i));
defparam desc402.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc403(.I0(s_output1[18:18]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_777_i));
defparam desc403.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc404(.I0(s_output1[19:19]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_778_i));
defparam desc404.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc405(.I0(s_output1[20:20]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_779_i));
defparam desc405.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc406(.I0(s_output1[21:21]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_780_i));
defparam desc406.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc407(.I0(s_output1[1:1]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_14_i));
defparam desc407.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc408(.I0(s_output1[3:3]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_18_i));
defparam desc408.INIT=64'h2222AAAA2232AAFA;
  LUT6_L desc409(.I0(s_output1[4:4]),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.I4(N_835),.I5(N_85),.LO(N_20_i));
defparam desc409.INIT=64'h2222AAAA2232AAFA;
  LUT5_L desc410(.I0(s_output1[22:22]),.I1(s_output1[23:23]),.I2(N_91),.I3(N_835),.I4(N_85),.LO(s_output_o_1));
defparam desc410.INIT=32'hCCCCC8C0;
  LUT6_L desc411(.I0(addsub_fract_o[12:12]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_60),.I5(N_68),.LO(N_1802_i));
defparam desc411.INIT=64'hA3A3A0A3A3A0A0A0;
  LUT6_L desc412(.I0(s_fracto28_1[4:4]),.I1(s_fracto28_1[27:27]),.I2(un3_s_fracto28_rnd_1_s_1),.I3(s_fracto28_rnd[3:3]),.I4(un3_s_fracto28_rnd_1_s_24),.I5(N_4),.LO(s_fracto28_2[3:3]));
defparam desc412.INIT=64'hBB88BB88F0F0FF00;
  LUT6 desc413(.I0(addsub_sign_o),.I1(s_fracto28_1[2:2]),.I2(s_fracto28_1[3:3]),.I3(s_rmode_i[1:1]),.I4(s_rmode_i[0:0]),.I5(s_roundup_1_3_i_a2_0),.O(s_fracto28_rnd[3:3]));
defparam desc413.INIT=64'h78F0B4305AF0A53C;
  LUT6_L desc414(.I0(s_fpu_op_i[1:1]),.I1(s_rmode_i[1:1]),.I2(un4_s_infa),.I3(un1_s_infb),.I4(div_zero_o_0),.I5(N_811_4),.LO(N_811_0_4));
defparam desc414.INIT=64'h0000000400000000;
  LUT6_L desc415(.I0(s_exp10_5_axb0),.I1(s_zeros_0_8),.I2(s_zeros_0_1),.I3(N_311),.I4(s_zeros_0_2),.I5(s_exp10[8:8]),.LO(s_expo9_1_4[0:0]));
defparam desc415.INIT=64'hFFFFFFFFAAAAAAA9;
  LUT6 desc416(.I0(s_output1[31:31]),.I1(s_rmode_i[1:1]),.I2(s_rmode_i[0:0]),.I3(un4_s_infa),.I4(un1_s_infb),.I5(div_zero_o_0),.O(N_85));
defparam desc416.INIT=64'hFFFFFFFFFFFFFF87;
  FD desc417(.Q(s_shr1),.D(s_shr1_0_0),.C(clk_i));
  LUT4 desc418(.I0(s_zeros_0_0[3:3]),.I1(s_zeros[4:4]),.I2(s_zeros_0_i_1_RNI027Q1[1:1]),.I3(s_zeros[0:0]),.O(un15_s_zero_fract_sn));
defparam desc418.INIT=16'h0800;
  LUT1 un3_s_fracto28_rnd_1_axb_24_cZ(.I0(s_fracto28_1[27:27]),.O(un3_s_fracto28_rnd_1_axb_24));
defparam un3_s_fracto28_rnd_1_axb_24_cZ.INIT=2'h2;
  LUT2 s_exp10_5_axb0_cZ(.I0(prenorm_addsub_exp_o[0:0]),.I1(addsub_fract_o[27:27]),.O(s_exp10_5_axb0));
defparam s_exp10_5_axb0_cZ.INIT=4'h9;
  LUT2 desc419(.I0(s_output1[31:31]),.I1(s_rmode_i[1:1]),.O(N_82));
defparam desc419.INIT=4'h7;
  LUT2_L desc420(.I0(s_exp10[1:1]),.I1(s_exp10[8:8]),.LO(s_expo9_1_4[1:1]));
defparam desc420.INIT=4'hE;
  LUT4 desc421(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[23:23]),.I2(addsub_fract_o[20:20]),.I3(addsub_fract_o[24:24]),.O(s_zeros_0_i_a2_2[1:1]));
defparam desc421.INIT=16'h0001;
  LUT4 desc422(.I0(s_output1[4:4]),.I1(s_output1[5:5]),.I2(s_output1[18:18]),.I3(s_output1[19:19]),.O(N_835_1_4));
defparam desc422.INIT=16'h0001;
  LUT4 desc423(.I0(s_output1[0:0]),.I1(s_output1[1:1]),.I2(s_output1[2:2]),.I3(s_output1[3:3]),.O(N_835_3_4));
defparam desc423.INIT=16'h0001;
  LUT4 desc424(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[19:19]),.I2(addsub_fract_o[21:21]),.I3(addsub_fract_o[23:23]),.O(N_338));
defparam desc424.INIT=16'h0001;
  LUT5 un11_s_exp10_7_3_cZ(.I0(s_exp10[0:0]),.I1(s_exp10[1:1]),.I2(s_exp10[2:2]),.I3(s_exp10[5:5]),.I4(s_exp10[6:6]),.O(un11_s_exp10_7_3));
defparam un11_s_exp10_7_3_cZ.INIT=32'h00000001;
  LUT6 desc425(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[21:21]),.I2(addsub_fract_o[23:23]),.I3(addsub_fract_o[22:22]),.I4(addsub_fract_o[24:24]),.I5(N_1861),.O(s_zeros_0_i_1[1:1]));
defparam desc425.INIT=64'hAAAAAFAEFFFFFFFF;
  LUT6 desc426(.I0(s_output1[7:7]),.I1(s_output1[8:8]),.I2(s_output1[9:9]),.I3(s_output1[10:10]),.I4(s_output1[11:11]),.I5(s_output1[12:12]),.O(N_835_0));
defparam desc426.INIT=64'h0000000000000001;
  LUT6 desc427(.I0(s_output1[6:6]),.I1(s_output1[13:13]),.I2(s_output1[14:14]),.I3(s_output1[15:15]),.I4(s_output1[16:16]),.I5(s_output1[17:17]),.O(N_835_2));
defparam desc427.INIT=64'h0000000000000001;
  LUT6_L desc428(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[6:6]),.I2(addsub_fract_o[1:1]),.I3(addsub_fract_o[2:2]),.I4(addsub_fract_o[4:4]),.I5(addsub_fract_o[3:3]),.LO(N_1692));
defparam desc428.INIT=64'hEEEEEEEEEEEEFFFE;
  LUT6 desc429(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[6:6]),.I2(addsub_fract_o[1:1]),.I3(addsub_fract_o[2:2]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1683));
defparam desc429.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6 desc430(.I0(addsub_fract_o[11:11]),.I1(addsub_fract_o[15:15]),.I2(addsub_fract_o[12:12]),.I3(addsub_fract_o[16:16]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1685));
defparam desc430.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc431(.I0(addsub_fract_o[9:9]),.I1(addsub_fract_o[13:13]),.I2(addsub_fract_o[10:10]),.I3(addsub_fract_o[14:14]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1686));
defparam desc431.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc432(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[17:17]),.I2(addsub_fract_o[20:20]),.I3(addsub_fract_o[18:18]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1695));
defparam desc432.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc433(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[6:6]),.I2(addsub_fract_o[9:9]),.I3(addsub_fract_o[10:10]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1696));
defparam desc433.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc434(.I0(addsub_fract_o[7:7]),.I1(addsub_fract_o[11:11]),.I2(addsub_fract_o[8:8]),.I3(addsub_fract_o[12:12]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1697));
defparam desc434.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc435(.I0(addsub_fract_o[13:13]),.I1(addsub_fract_o[17:17]),.I2(addsub_fract_o[14:14]),.I3(addsub_fract_o[18:18]),.I4(s_shl1[2:2]),.I5(s_shl1[0:0]),.O(N_1720));
defparam desc435.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc436(.I0(addsub_fract_o[15:15]),.I1(addsub_fract_o[17:17]),.I2(addsub_fract_o[16:16]),.I3(addsub_fract_o[18:18]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1721));
defparam desc436.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc437(.I0(addsub_fract_o[13:13]),.I1(addsub_fract_o[15:15]),.I2(addsub_fract_o[14:14]),.I3(addsub_fract_o[16:16]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1722));
defparam desc437.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc438(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[21:21]),.I2(addsub_fract_o[22:22]),.I3(addsub_fract_o[20:20]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1827));
defparam desc438.INIT=64'h5555333300FF0F0F;
  LUT6 desc439(.I0(addsub_fract_o[21:21]),.I1(addsub_fract_o[23:23]),.I2(addsub_fract_o[22:22]),.I3(addsub_fract_o[24:24]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1837));
defparam desc439.INIT=64'h555533330F0F00FF;
  LUT6 desc440(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[26:26]),.I2(addsub_fract_o[23:23]),.I3(addsub_fract_o[24:24]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1850));
defparam desc440.INIT=64'h0F0F555500FF3333;
  LUT6 desc441(.I0(addsub_fract_o[11:11]),.I1(addsub_fract_o[13:13]),.I2(addsub_fract_o[15:15]),.I3(addsub_fract_o[17:17]),.I4(addsub_fract_o[14:14]),.I5(N_338),.O(s_zeros_0_a2_3[4:4]));
defparam desc441.INIT=64'hFFFFFFFEFFFFFFFF;
  LUT6 desc442(.I0(addsub_fract_o[1:1]),.I1(addsub_fract_o[2:2]),.I2(addsub_fract_o[0:0]),.I3(s_shl1[2:2]),.I4(s_shl1[1:1]),.I5(s_shl1[0:0]),.O(N_1673));
defparam desc442.INIT=64'hFFFFFF55FF0FFF33;
  LUT6 un2_s_overflow_o_i_o2_0_1(.I0(s_output1[27:27]),.I1(s_output1[28:28]),.I2(s_output1[25:25]),.I3(s_output1[26:26]),.I4(s_output1[30:30]),.I5(N_91_0_0_1),.O(N_91));
defparam un2_s_overflow_o_i_o2_0_1.INIT=64'hFFFFFFFF7FFFFFFF;
  LUT6 s_roundup_1_3_i(.I0(addsub_sign_o),.I1(s_fracto28_1[2:2]),.I2(s_fracto28_1[3:3]),.I3(s_rmode_i[1:1]),.I4(s_rmode_i[0:0]),.I5(s_roundup_1_3_i_a2_0),.O(N_4));
defparam s_roundup_1_3_i.INIT=64'h77FFBB3F55FFAA33;
  LUT5 desc443(.I0(addsub_fract_o[0:0]),.I1(s_shl1[2:2]),.I2(s_shl1[1:1]),.I3(s_shl1[0:0]),.I4(N_1723),.O(N_61));
defparam desc443.INIT=32'h333B0008;
  LUT6 desc444(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1701),.I3(N_1713),.I4(N_1709),.I5(N_1708),.O(N_1803));
defparam desc444.INIT=64'h028A46CE139B57DF;
  LUT6 desc445(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1701),.I3(N_1709),.I4(N_1708),.I5(N_1707),.O(N_1807));
defparam desc445.INIT=64'h082A4C6E193B5D7F;
  LUT6 desc446(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_6),.I3(N_8),.I4(N_1712),.I5(N_1713),.O(N_1808));
defparam desc446.INIT=64'h02468ACE13579BDF;
  LUT6 desc447(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1706),.I3(N_1709),.I4(N_1708),.I5(N_1707),.O(N_1815));
defparam desc447.INIT=64'h018923AB45CD67EF;
  LUT6 desc448(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1705),.I3(N_1706),.I4(N_1708),.I5(N_1707),.O(N_1821));
defparam desc448.INIT=64'h014589CD2367ABEF;
  LUT6 desc449(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_8),.I3(N_1701),.I4(N_1713),.I5(N_1709),.O(N_1822));
defparam desc449.INIT=64'h084C2A6E195D3B7F;
  LUT6 desc450(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1700),.I3(N_1705),.I4(N_1706),.I5(N_1707),.O(N_1832));
defparam desc450.INIT=64'h0145236789CDABEF;
  LUT6 desc451(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1842),.I3(N_1700),.I4(N_1705),.I5(N_1706),.O(N_1844));
defparam desc451.INIT=64'h1054327698DCBAFE;
  LUT6 desc452(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_1855),.I3(N_1842),.I4(N_1700),.I5(N_1705),.O(N_1857));
defparam desc452.INIT=64'h54107632DC98FEBA;
  LUT5 desc453(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_6),.I3(N_1711),.I4(N_1712),.O(N_62));
defparam desc453.INIT=32'h76543210;
  LUT6 desc454(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_6),.I3(N_8),.I4(N_1711),.I5(N_1712),.O(N_64));
defparam desc454.INIT=64'hFBEA7362D9C85140;
  LUT6 desc455(.I0(s_shl1[2:2]),.I1(s_shl1[1:1]),.I2(N_6),.I3(N_8),.I4(N_1701),.I5(N_1713),.O(N_68));
defparam desc455.INIT=64'hF7D5E6C4B391A280;
  LUT6 desc456(.I0(addsub_fract_o[15:15]),.I1(addsub_fract_o[16:16]),.I2(N_299_2),.I3(N_338),.I4(N_289),.I5(s_zeros_0_a2_0_2[3:3]),.O(s_zeros_0_0[3:3]));
defparam desc456.INIT=64'hFF00FF00FF00FE00;
  LUT6 desc457(.I0(addsub_fract_o[22:22]),.I1(addsub_fract_o[20:20]),.I2(addsub_fract_o[24:24]),.I3(addsub_fract_o[16:16]),.I4(addsub_fract_o[18:18]),.I5(N_1861),.O(N_337));
defparam desc457.INIT=64'h0000000100000000;
  LUT6 desc458(.I0(addsub_fract_o[15:15]),.I1(addsub_fract_o[17:17]),.I2(addsub_fract_o[16:16]),.I3(addsub_fract_o[18:18]),.I4(N_289),.I5(N_1872),.O(N_1877));
defparam desc458.INIT=64'h0001000100010000;
  LUT6 desc459(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[1:1]),.I2(addsub_fract_o[2:2]),.I3(addsub_fract_o[4:4]),.I4(addsub_fract_o[0:0]),.I5(addsub_fract_o[3:3]),.O(s_zeros_0_8_tz));
defparam desc459.INIT=64'hAAFFAAFFAAAEAAAF;
  LUT5 un1_s_exp10_3_cZ(.I0(s_exp10[3:3]),.I1(s_exp10[4:4]),.I2(s_exp10[7:7]),.I3(s_exp10[8:8]),.I4(un11_s_exp10_7_3),.O(un1_s_exp10_3));
defparam un1_s_exp10_3_cZ.INIT=32'h00FE00FF;
  LUT3 desc460(.I0(s_fracto28_1[27:27]),.I1(un3_s_fracto28_rnd_1_s_24),.I2(N_4),.O(s_fracto28_rnd[27:27]));
defparam desc460.INIT=8'hAC;
  LUT6 desc461(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[21:21]),.I2(addsub_fract_o[23:23]),.I3(addsub_fract_o[22:22]),.I4(addsub_fract_o[24:24]),.I5(N_1861),.O(s_zeros_0_0[0:0]));
defparam desc461.INIT=64'hAAAAFAFE00000000;
  LUT6 desc462(.I0(addsub_fract_o[0:0]),.I1(s_shl1[2:2]),.I2(s_shl1[1:1]),.I3(s_shl1[0:0]),.I4(N_1676),.I5(N_1683),.O(N_63));
defparam desc462.INIT=64'h3FBF0F8F30B00080;
  LUT6 desc463(.I0(s_output1[20:20]),.I1(s_output1[21:21]),.I2(N_835_1_4),.I3(N_835_3_4),.I4(N_835_0),.I5(N_835_2),.O(N_835));
defparam desc463.INIT=64'h1000000000000000;
  LUT6_L desc464(.I0(addsub_fract_o[13:13]),.I1(addsub_fract_o[15:15]),.I2(addsub_fract_o[14:14]),.I3(addsub_fract_o[16:16]),.I4(addsub_fract_o[18:18]),.I5(N_331),.LO(s_zeros_0_4));
defparam desc464.INIT=64'h000000CE00000000;
  LUT4_L desc465(.I0(s_expo9_1[3:3]),.I1(s_expo9_1[2:2]),.I2(s_expo9_1[1:1]),.I3(s_expo9_1[0:0]),.LO(s_expo9_0_c4));
defparam desc465.INIT=16'hFFFE;
  LUT6_L desc466(.I0(addsub_fract_o[9:9]),.I1(addsub_fract_o[11:11]),.I2(addsub_fract_o[10:10]),.I3(addsub_fract_o[12:12]),.I4(N_1774),.I5(N_1692),.LO(N_1769));
defparam desc466.INIT=64'h0033003200320032;
  LUT5_L desc467(.I0(addsub_fract_o[1:1]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_1776),.LO(s_fracto28_1_3[0:0]));
defparam desc467.INIT=32'hA0A3A0A0;
  LUT5 desc468(.I0(s_shl1[1:1]),.I1(s_shl1[3:3]),.I2(N_1696),.I3(N_1673),.I4(N_1684),.O(N_1797));
defparam desc468.INIT=32'hCD01EF23;
  LUT5_L desc469(.I0(s_shl1[2:2]),.I1(s_shl1[3:3]),.I2(N_1721),.I3(N_1827),.I4(N_1727),.LO(N_1829));
defparam desc469.INIT=32'h1302DFCE;
  LUT5 desc470(.I0(s_shl1[2:2]),.I1(s_shl1[3:3]),.I2(N_1722),.I3(N_1695),.I4(N_1726),.O(N_105));
defparam desc470.INIT=32'hFDEC3120;
  LUT5_L desc471(.I0(s_shl1[2:2]),.I1(s_shl1[3:3]),.I2(N_1850),.I3(N_1827),.I4(N_1725_i),.LO(N_1852));
defparam desc471.INIT=32'hFEDC3210;
  LUT5_L desc472(.I0(s_shl1[2:2]),.I1(s_shl1[3:3]),.I2(N_1837),.I3(N_1695),.I4(N_1693),.LO(N_1839));
defparam desc472.INIT=32'h1032DCFE;
  LUT6_L un12_s_exp10_cZ(.I0(s_exp10[3:3]),.I1(s_exp10[4:4]),.I2(s_exp10[9:9]),.I3(s_exp10[7:7]),.I4(s_exp10[8:8]),.I5(un11_s_exp10_7_3),.LO(un12_s_exp10));
defparam un12_s_exp10_cZ.INIT=64'hF0F0F0F1F0F0F0F0;
  LUT5 desc473(.I0(s_shl1[1:1]),.I1(s_shl1[3:3]),.I2(N_1776),.I3(N_1683),.I4(N_1684),.O(N_93));
defparam desc473.INIT=32'hF3D1E2C0;
  LUT6 desc474(.I0(s_fracto28_1[25:25]),.I1(s_fracto28_1[26:26]),.I2(un3_s_fracto28_rnd_1_s_23),.I3(un3_s_fracto28_rnd_1_s_22),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.O(s_fracto28_2[25:25]));
defparam desc474.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6_L desc475(.I0(s_fracto28_1[4:4]),.I1(s_fracto28_1[5:5]),.I2(un3_s_fracto28_rnd_1_s_1),.I3(un3_s_fracto28_rnd_1_s_2),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[4:4]));
defparam desc475.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc476(.I0(s_fracto28_1[5:5]),.I1(s_fracto28_1[6:6]),.I2(un3_s_fracto28_rnd_1_s_2),.I3(un3_s_fracto28_rnd_1_s_3),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[5:5]));
defparam desc476.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc477(.I0(s_fracto28_1[6:6]),.I1(s_fracto28_1[7:7]),.I2(un3_s_fracto28_rnd_1_s_3),.I3(un3_s_fracto28_rnd_1_s_4),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[6:6]));
defparam desc477.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc478(.I0(s_fracto28_1[7:7]),.I1(s_fracto28_1[8:8]),.I2(un3_s_fracto28_rnd_1_s_4),.I3(un3_s_fracto28_rnd_1_s_5),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[7:7]));
defparam desc478.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc479(.I0(s_fracto28_1[8:8]),.I1(s_fracto28_1[9:9]),.I2(un3_s_fracto28_rnd_1_s_5),.I3(un3_s_fracto28_rnd_1_s_6),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[8:8]));
defparam desc479.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc480(.I0(s_fracto28_1[9:9]),.I1(s_fracto28_1[10:10]),.I2(un3_s_fracto28_rnd_1_s_6),.I3(un3_s_fracto28_rnd_1_s_7),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[9:9]));
defparam desc480.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc481(.I0(s_fracto28_1[10:10]),.I1(s_fracto28_1[11:11]),.I2(un3_s_fracto28_rnd_1_s_7),.I3(un3_s_fracto28_rnd_1_s_8),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[10:10]));
defparam desc481.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc482(.I0(s_fracto28_1[11:11]),.I1(s_fracto28_1[12:12]),.I2(un3_s_fracto28_rnd_1_s_8),.I3(un3_s_fracto28_rnd_1_s_9),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[11:11]));
defparam desc482.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc483(.I0(s_fracto28_1[12:12]),.I1(s_fracto28_1[13:13]),.I2(un3_s_fracto28_rnd_1_s_9),.I3(un3_s_fracto28_rnd_1_s_10),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[12:12]));
defparam desc483.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc484(.I0(s_fracto28_1[13:13]),.I1(s_fracto28_1[14:14]),.I2(un3_s_fracto28_rnd_1_s_10),.I3(un3_s_fracto28_rnd_1_s_11),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[13:13]));
defparam desc484.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc485(.I0(s_fracto28_1[14:14]),.I1(s_fracto28_1[15:15]),.I2(un3_s_fracto28_rnd_1_s_11),.I3(un3_s_fracto28_rnd_1_s_12),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[14:14]));
defparam desc485.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc486(.I0(s_fracto28_1[15:15]),.I1(s_fracto28_1[16:16]),.I2(un3_s_fracto28_rnd_1_s_12),.I3(un3_s_fracto28_rnd_1_s_13),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[15:15]));
defparam desc486.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc487(.I0(s_fracto28_1[16:16]),.I1(s_fracto28_1[17:17]),.I2(un3_s_fracto28_rnd_1_s_13),.I3(un3_s_fracto28_rnd_1_s_14),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[16:16]));
defparam desc487.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc488(.I0(s_fracto28_1[17:17]),.I1(s_fracto28_1[18:18]),.I2(un3_s_fracto28_rnd_1_s_14),.I3(un3_s_fracto28_rnd_1_s_15),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[17:17]));
defparam desc488.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc489(.I0(s_fracto28_1[22:22]),.I1(s_fracto28_1[23:23]),.I2(un3_s_fracto28_rnd_1_s_19),.I3(un3_s_fracto28_rnd_1_s_20),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[22:22]));
defparam desc489.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc490(.I0(s_fracto28_1[23:23]),.I1(s_fracto28_1[24:24]),.I2(un3_s_fracto28_rnd_1_s_20),.I3(un3_s_fracto28_rnd_1_s_21),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[23:23]));
defparam desc490.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc491(.I0(s_fracto28_1[24:24]),.I1(s_fracto28_1[25:25]),.I2(un3_s_fracto28_rnd_1_s_21),.I3(un3_s_fracto28_rnd_1_s_22),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[24:24]));
defparam desc491.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6 desc492(.I0(s_output1[24:24]),.I1(s_output1[25:25]),.I2(s_output1[26:26]),.I3(s_output1[30:30]),.I4(N_844_0_4),.I5(N_835),.O(N_811_4));
defparam desc492.INIT=64'h0001000000000000;
  LUT2 un2_s_inf_o_i_a2(.I0(s_output1[22:22]),.I1(N_835),.O(N_836));
defparam un2_s_inf_o_i_a2.INIT=4'h8;
  LUT6_L desc493(.I0(s_fracto28_1[21:21]),.I1(s_fracto28_1[22:22]),.I2(un3_s_fracto28_rnd_1_s_18),.I3(un3_s_fracto28_rnd_1_s_19),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[21:21]));
defparam desc493.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc494(.I0(s_fracto28_1[20:20]),.I1(s_fracto28_1[21:21]),.I2(un3_s_fracto28_rnd_1_s_17),.I3(un3_s_fracto28_rnd_1_s_18),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[20:20]));
defparam desc494.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc495(.I0(s_fracto28_1[19:19]),.I1(s_fracto28_1[20:20]),.I2(un3_s_fracto28_rnd_1_s_16),.I3(un3_s_fracto28_rnd_1_s_17),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[19:19]));
defparam desc495.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L desc496(.I0(s_fracto28_1[18:18]),.I1(s_fracto28_1[19:19]),.I2(un3_s_fracto28_rnd_1_s_15),.I3(un3_s_fracto28_rnd_1_s_16),.I4(N_4),.I5(s_fracto28_rnd[27:27]),.LO(s_fracto28_2[18:18]));
defparam desc496.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6 un6_s_expo9_3_ac0_5(.I0(s_expo9_1[3:3]),.I1(s_expo9_1[2:2]),.I2(s_expo9_1[1:1]),.I3(s_expo9_1[0:0]),.I4(s_fracto28_1[26:26]),.I5(s_fracto28_1[27:27]),.O(un6_s_expo9_3_c4));
defparam un6_s_expo9_3_ac0_5.INIT=64'h8000800080000001;
  LUT6 desc497(.I0(prenorm_addsub_exp_o[4:4]),.I1(prenorm_addsub_exp_o[3:3]),.I2(prenorm_addsub_exp_o[2:2]),.I3(result_1),.I4(s_exp10[8:8]),.I5(un12_s_exp10),.O(un1_s_exp10_1));
defparam desc497.INIT=64'h00010001FFFF0000;
  LUT6_L desc498(.I0(prenorm_addsub_exp_o[3:3]),.I1(prenorm_addsub_exp_o[2:2]),.I2(result_1),.I3(N_331),.I4(s_zeros_0_0[3:3]),.I5(un1_s_exp10_3),.LO(N_391));
defparam desc498.INIT=64'hFF000000A9A9A9A9;
  LUT6_L desc499(.I0(s_shl1[4:4]),.I1(s_shl1[3:3]),.I2(N_58),.I3(N_1844),.I4(N_1807),.I5(N_1808),.LO(N_1847));
defparam desc499.INIT=64'h7F6E3B2A5D4C1908;
  LUT6 desc500(.I0(addsub_fract_o[9:9]),.I1(addsub_fract_o[11:11]),.I2(addsub_fract_o[10:10]),.I3(addsub_fract_o[12:12]),.I4(addsub_fract_o[14:14]),.I5(N_337),.O(s_zeros_0_2));
defparam desc500.INIT=64'h000000CE00000000;
  LUT6 desc501(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[17:17]),.I2(addsub_fract_o[18:18]),.I3(N_331),.I4(s_zeros_0_0[0:0]),.I5(s_zeros_0_4),.O(s_zeros_0_1));
defparam desc501.INIT=64'hFFFFFFFFFFFFAE00;
  LUT6 desc502(.I0(addsub_fract_o[6:6]),.I1(addsub_fract_o[8:8]),.I2(addsub_fract_o[10:10]),.I3(addsub_fract_o[14:14]),.I4(s_zeros_0_8_tz),.I5(N_345),.O(s_zeros_0_8));
defparam desc502.INIT=64'h0001000000000000;
  LUT6 desc503(.I0(addsub_fract_o[7:7]),.I1(addsub_fract_o[8:8]),.I2(addsub_fract_o[10:10]),.I3(addsub_fract_o[12:12]),.I4(addsub_fract_o[14:14]),.I5(N_337),.O(N_311));
defparam desc503.INIT=64'h0000000200000000;
  LUT5 desc504(.I0(prenorm_addsub_exp_o[5:5]),.I1(prenorm_addsub_exp_o[4:4]),.I2(prenorm_addsub_exp_o[3:3]),.I3(prenorm_addsub_exp_o[2:2]),.I4(s_exp10_5_c2),.O(s_exp10_5_i[5:5]));
defparam desc504.INIT=32'h95555555;
  LUT5 desc505(.I0(addsub_fract_o[13:13]),.I1(addsub_fract_o[15:15]),.I2(addsub_fract_o[14:14]),.I3(addsub_fract_o[16:16]),.I4(N_1769),.O(N_1770));
defparam desc505.INIT=32'h00330032;
  LUT5_L desc506(.I0(addsub_fract_o[2:2]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_58),.LO(N_1779_i));
defparam desc506.INIT=32'hA0A3A0A0;
  LUT6_L desc507(.I0(prenorm_addsub_exp_o[2:2]),.I1(result_1),.I2(m149_e_1),.I3(m149_0),.I4(N_1877),.I5(un1_s_exp10_3),.LO(N_390));
defparam desc507.INIT=64'hFF000F0099999999;
  LUT6_L desc508(.I0(prenorm_addsub_exp_o[4:4]),.I1(prenorm_addsub_exp_o[3:3]),.I2(prenorm_addsub_exp_o[2:2]),.I3(result_1),.I4(s_zeros[4:4]),.I5(un1_s_exp10_3),.LO(N_392));
defparam desc508.INIT=64'hFFFF0000AAA9AAA9;
  LUT6_L desc509(.I0(addsub_fract_o[10:10]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_58),.I5(N_1808),.LO(s_fracto28_1_3[9:9]));
defparam desc509.INIT=64'hA3A0A0A0A3A3A0A3;
  LUT6_L desc510(.I0(addsub_fract_o[13:13]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_61),.I5(N_1726),.LO(s_fracto28_1_3[12:12]));
defparam desc510.INIT=64'hA3A3A0A3A3A0A0A0;
  LUT6_L desc511(.I0(addsub_fract_o[14:14]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_62),.I5(N_1822),.LO(s_fracto28_1_3[13:13]));
defparam desc511.INIT=64'hA3A0A0A0A3A3A0A3;
  LUT6 desc512(.I0(s_expo9_1[4:4]),.I1(s_expo9_1[3:3]),.I2(s_expo9_1[2:2]),.I3(s_expo9_1[1:1]),.I4(s_expo9_1[0:0]),.I5(un2_s_expo9_2),.O(s_expo9_2[4:4]));
defparam desc512.INIT=64'hAAAAAAA9AAAAAAAA;
  LUT5_L desc513(.I0(addsub_fract_o[4:4]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_60),.LO(N_1784_i));
defparam desc513.INIT=32'hA0A3A0A0;
  LUT5_L desc514(.I0(addsub_fract_o[3:3]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_1673),.LO(N_1781_i));
defparam desc514.INIT=32'hA0A0A0A3;
  LUT6_L desc515(.I0(addsub_fract_o[17:17]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_1776),.I5(N_1729),.LO(s_fracto28_1_3[16:16]));
defparam desc515.INIT=64'hA3AFA3A3A0ACA0A0;
  LUT6 desc516(.I0(prenorm_addsub_exp_o[6:6]),.I1(prenorm_addsub_exp_o[5:5]),.I2(prenorm_addsub_exp_o[4:4]),.I3(prenorm_addsub_exp_o[3:3]),.I4(prenorm_addsub_exp_o[2:2]),.I5(s_exp10_5_c2),.O(s_exp10_5_i[6:6]));
defparam desc516.INIT=64'h9555555555555555;
  LUT5_L desc517(.I0(addsub_fract_o[8:8]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_64),.LO(N_1795_i));
defparam desc517.INIT=32'hA0A3A0A0;
  LUT5_L desc518(.I0(addsub_fract_o[6:6]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_62),.LO(N_1790_i));
defparam desc518.INIT=32'hA0A3A0A0;
  LUT5_L desc519(.I0(addsub_fract_o[5:5]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_61),.LO(N_1787_i));
defparam desc519.INIT=32'hA0A3A0A0;
  LUT4_L desc520(.I0(addsub_fract_o[11:11]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(N_1797),.LO(N_1799_i));
defparam desc520.INIT=16'hA0A3;
  LUT6_L desc521(.I0(addsub_fract_o[16:16]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_1803),.I5(N_64),.LO(N_1806_i));
defparam desc521.INIT=64'hA3A0A3A3A0A0A0A3;
  LUT6 s_exp10_5_ac0_13_i_cZ(.I0(prenorm_addsub_exp_o[7:7]),.I1(prenorm_addsub_exp_o[6:6]),.I2(prenorm_addsub_exp_o[5:5]),.I3(prenorm_addsub_exp_o[4:4]),.I4(prenorm_addsub_exp_o[3:3]),.I5(s_exp10_5_c3),.O(s_exp10_5_ac0_13_i));
defparam s_exp10_5_ac0_13_i_cZ.INIT=64'h7FFFFFFFFFFFFFFF;
  LUT6 desc522(.I0(prenorm_addsub_exp_o[7:7]),.I1(prenorm_addsub_exp_o[6:6]),.I2(prenorm_addsub_exp_o[5:5]),.I3(prenorm_addsub_exp_o[4:4]),.I4(prenorm_addsub_exp_o[3:3]),.I5(s_exp10_5_c3),.O(s_exp10_5_i[7:7]));
defparam desc522.INIT=64'h9555555555555555;
  LUT6_L desc523(.I0(addsub_fract_o[15:15]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_63),.I5(N_1727),.LO(s_fracto28_1_3[14:14]));
defparam desc523.INIT=64'hA3A3A0A3A3A0A0A0;
  LUT4_L desc524(.I0(addsub_fract_o[9:9]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(N_93),.LO(N_1796_i));
defparam desc524.INIT=16'hA3A0;
  LUT5_L desc525(.I0(addsub_fract_o[27:27]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(N_1797),.I4(N_1852),.LO(N_1854_i));
defparam desc525.INIT=32'hA0ACA3AF;
  LUT3_L desc526(.I0(addsub_fract_o[26:26]),.I1(s_shr1),.I2(N_1847),.LO(N_1848_i));
defparam desc526.INIT=8'h8B;
  LUT6_L desc527(.I0(addsub_fract_o[24:24]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_64),.I5(N_1833),.LO(N_1835_i));
defparam desc527.INIT=64'hA0ACA0A0A3AFA3A3;
  LUT6_L desc528(.I0(addsub_fract_o[22:22]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_62),.I5(N_1823),.LO(N_1825_i));
defparam desc528.INIT=64'hA0ACA0A0A3AFA3A3;
  LUT6_L desc529(.I0(addsub_fract_o[21:21]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_61),.I5(N_105),.LO(N_1820_i));
defparam desc529.INIT=64'hA3AFA3A3A0ACA0A0;
  LUT6_L desc530(.I0(addsub_fract_o[20:20]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_60),.I5(N_1816),.LO(N_1818_i));
defparam desc530.INIT=64'hA0ACA0A0A3AFA3A3;
  LUT6_L desc531(.I0(addsub_fract_o[19:19]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_1673),.I5(N_1812),.LO(N_1814_i));
defparam desc531.INIT=64'hA0A0A0ACA3A3A3AF;
  LUT6_L desc532(.I0(addsub_fract_o[18:18]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_58),.I5(N_1809),.LO(N_1811_i));
defparam desc532.INIT=64'hA0ACA0A0A3AFA3A3;
  LUT5_L desc533(.I0(addsub_fract_o[7:7]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_63),.LO(N_28_0_i));
defparam desc533.INIT=32'hA0A3A0A0;
  LUT5_L desc534(.I0(addsub_fract_o[25:25]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(N_93),.I4(N_1839),.LO(N_1841_i));
defparam desc534.INIT=32'hACA0AFA3;
  LUT6_L desc535(.I0(addsub_fract_o[23:23]),.I1(s_shl1[4:4]),.I2(s_shr1),.I3(s_shl1[3:3]),.I4(N_63),.I5(N_1829),.LO(N_1831_i));
defparam desc535.INIT=64'hA0ACA0A0A3AFA3A3;
  LUT6_L desc536(.I0(addsub_sign_o),.I1(s_opa_i[31:31]),.I2(s_opb_i_27),.I3(N_1979),.I4(N_36_0),.I5(N_1948),.LO(N_3392_mux));
defparam desc536.INIT=64'hAAAAAAAAAACCF0F0;
  LUT6 desc537(.I0(s_expo9_1[3:3]),.I1(s_expo9_1[2:2]),.I2(s_expo9_1[1:1]),.I3(s_expo9_1[0:0]),.I4(un2_s_expo9_2),.I5(un1_s_expo9_3),.O(s_expo9_3[3:3]));
defparam desc537.INIT=64'hAAAA6AAAAAA9AAAA;
  LUT4 s_overflow_0_0_cZ(.I0(un6_s_expo9_3_c4),.I1(s_expo9_2[5:5]),.I2(s_expo9_2[4:4]),.I3(un1_s_expo9_3),.O(s_overflow_0_0));
defparam s_overflow_0_0_cZ.INIT=16'h48C0;
  LUT6 desc538(.I0(s_expo9_1[2:2]),.I1(s_expo9_1[1:1]),.I2(s_expo9_1[0:0]),.I3(un2_s_expo9_2),.I4(un1_s_expo9_3),.I5(un15_s_zero_fract_sn),.O(s_output_o_m0[25:25]));
defparam desc538.INIT=64'h00000000AA6AA9AA;
  LUT3_L s_overflow_2_cZ(.I0(s_expo9_3[6:6]),.I1(s_expo9_3[7:7]),.I2(s_expo9_3[3:3]),.LO(s_overflow_2));
defparam s_overflow_2_cZ.INIT=8'h80;
  LUT6 s_overflow_cZ(.I0(s_expo9_1[0:0]),.I1(un2_s_expo9_2),.I2(un1_s_expo9_3),.I3(s_overflow_0_0),.I4(s_overflow_1),.I5(s_overflow_2),.O(s_overflow));
defparam s_overflow_cZ.INIT=64'h9600000000000000;
  LUT6_L desc539(.I0(un4_s_infa),.I1(un1_s_infb),.I2(s_fracto28_2[25:25]),.I3(N_1948),.I4(un15_s_zero_fract_sn),.I5(s_overflow),.LO(s_output_o[22:22]));
defparam desc539.INIT=64'h00FF00FF00EE10FE;
  LUT5 s_exp10_5_ac0_1_lut6_2_RNI8F6F6(.I0(prenorm_addsub_exp_o[2:2]),.I1(m149_e_1),.I2(s_exp10_5_c2),.I3(m149_0),.I4(N_1877),.O(s_exp10_axb_2));
defparam s_exp10_5_ac0_1_lut6_2_RNI8F6F6.INIT=32'h5AA596A5;
  LUT5 desc540(.I0(addsub_fract_o[20:20]),.I1(prenorm_addsub_exp_o[3:3]),.I2(N_329),.I3(s_exp10_5_c3),.I4(s_zeros_0_0[3:3]),.O(s_exp10_axb_3));
defparam desc540.INIT=32'h9C63CC33;
  LUT5 s_exp10_5_ac0_5_lut6_2_RNIEJ5Q(.I0(prenorm_addsub_exp_o[4:4]),.I1(addsub_fract_o[12:12]),.I2(s_exp10_5_c4),.I3(s_zeros_0_a2_3[4:4]),.I4(N_337),.O(s_exp10_axb_4));
defparam s_exp10_5_ac0_5_lut6_2_RNIEJ5Q.INIT=32'hA596A5A5;
  XORCY un3_s_fracto28_rnd_1_s_24_cZ(.LI(un3_s_fracto28_rnd_1_axb_24),.CI(un3_s_fracto28_rnd_1_cry_23),.O(un3_s_fracto28_rnd_1_s_24));
  XORCY un3_s_fracto28_rnd_1_s_23_cZ(.LI(un3_s_fracto28_rnd_1_axb_23),.CI(un3_s_fracto28_rnd_1_cry_22),.O(un3_s_fracto28_rnd_1_s_23));
  MUXCY_L un3_s_fracto28_rnd_1_cry_23_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_22),.S(un3_s_fracto28_rnd_1_axb_23),.LO(un3_s_fracto28_rnd_1_cry_23));
  XORCY un3_s_fracto28_rnd_1_s_22_cZ(.LI(un3_s_fracto28_rnd_1_axb_22),.CI(un3_s_fracto28_rnd_1_cry_21),.O(un3_s_fracto28_rnd_1_s_22));
  MUXCY_L un3_s_fracto28_rnd_1_cry_22_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_21),.S(un3_s_fracto28_rnd_1_axb_22),.LO(un3_s_fracto28_rnd_1_cry_22));
  XORCY un3_s_fracto28_rnd_1_s_21_cZ(.LI(un3_s_fracto28_rnd_1_axb_21),.CI(un3_s_fracto28_rnd_1_cry_20),.O(un3_s_fracto28_rnd_1_s_21));
  MUXCY_L un3_s_fracto28_rnd_1_cry_21_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_20),.S(un3_s_fracto28_rnd_1_axb_21),.LO(un3_s_fracto28_rnd_1_cry_21));
  XORCY un3_s_fracto28_rnd_1_s_20_cZ(.LI(un3_s_fracto28_rnd_1_axb_20),.CI(un3_s_fracto28_rnd_1_cry_19),.O(un3_s_fracto28_rnd_1_s_20));
  MUXCY_L un3_s_fracto28_rnd_1_cry_20_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_19),.S(un3_s_fracto28_rnd_1_axb_20),.LO(un3_s_fracto28_rnd_1_cry_20));
  XORCY un3_s_fracto28_rnd_1_s_19_cZ(.LI(un3_s_fracto28_rnd_1_axb_19),.CI(un3_s_fracto28_rnd_1_cry_18),.O(un3_s_fracto28_rnd_1_s_19));
  MUXCY_L un3_s_fracto28_rnd_1_cry_19_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_18),.S(un3_s_fracto28_rnd_1_axb_19),.LO(un3_s_fracto28_rnd_1_cry_19));
  XORCY un3_s_fracto28_rnd_1_s_18_cZ(.LI(un3_s_fracto28_rnd_1_axb_18),.CI(un3_s_fracto28_rnd_1_cry_17),.O(un3_s_fracto28_rnd_1_s_18));
  MUXCY_L un3_s_fracto28_rnd_1_cry_18_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_17),.S(un3_s_fracto28_rnd_1_axb_18),.LO(un3_s_fracto28_rnd_1_cry_18));
  XORCY un3_s_fracto28_rnd_1_s_17_cZ(.LI(un3_s_fracto28_rnd_1_axb_17),.CI(un3_s_fracto28_rnd_1_cry_16),.O(un3_s_fracto28_rnd_1_s_17));
  MUXCY_L un3_s_fracto28_rnd_1_cry_17_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_16),.S(un3_s_fracto28_rnd_1_axb_17),.LO(un3_s_fracto28_rnd_1_cry_17));
  XORCY un3_s_fracto28_rnd_1_s_16_cZ(.LI(un3_s_fracto28_rnd_1_axb_16),.CI(un3_s_fracto28_rnd_1_cry_15),.O(un3_s_fracto28_rnd_1_s_16));
  MUXCY_L un3_s_fracto28_rnd_1_cry_16_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_15),.S(un3_s_fracto28_rnd_1_axb_16),.LO(un3_s_fracto28_rnd_1_cry_16));
  XORCY un3_s_fracto28_rnd_1_s_15_cZ(.LI(un3_s_fracto28_rnd_1_axb_15),.CI(un3_s_fracto28_rnd_1_cry_14),.O(un3_s_fracto28_rnd_1_s_15));
  MUXCY_L un3_s_fracto28_rnd_1_cry_15_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_14),.S(un3_s_fracto28_rnd_1_axb_15),.LO(un3_s_fracto28_rnd_1_cry_15));
  XORCY un3_s_fracto28_rnd_1_s_14_cZ(.LI(un3_s_fracto28_rnd_1_axb_14),.CI(un3_s_fracto28_rnd_1_cry_13),.O(un3_s_fracto28_rnd_1_s_14));
  MUXCY_L un3_s_fracto28_rnd_1_cry_14_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_13),.S(un3_s_fracto28_rnd_1_axb_14),.LO(un3_s_fracto28_rnd_1_cry_14));
  XORCY un3_s_fracto28_rnd_1_s_13_cZ(.LI(un3_s_fracto28_rnd_1_axb_13),.CI(un3_s_fracto28_rnd_1_cry_12),.O(un3_s_fracto28_rnd_1_s_13));
  MUXCY_L un3_s_fracto28_rnd_1_cry_13_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_12),.S(un3_s_fracto28_rnd_1_axb_13),.LO(un3_s_fracto28_rnd_1_cry_13));
  XORCY un3_s_fracto28_rnd_1_s_12_cZ(.LI(un3_s_fracto28_rnd_1_axb_12),.CI(un3_s_fracto28_rnd_1_cry_11),.O(un3_s_fracto28_rnd_1_s_12));
  MUXCY_L un3_s_fracto28_rnd_1_cry_12_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_11),.S(un3_s_fracto28_rnd_1_axb_12),.LO(un3_s_fracto28_rnd_1_cry_12));
  XORCY un3_s_fracto28_rnd_1_s_11_cZ(.LI(un3_s_fracto28_rnd_1_axb_11),.CI(un3_s_fracto28_rnd_1_cry_10),.O(un3_s_fracto28_rnd_1_s_11));
  MUXCY_L un3_s_fracto28_rnd_1_cry_11_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_10),.S(un3_s_fracto28_rnd_1_axb_11),.LO(un3_s_fracto28_rnd_1_cry_11));
  XORCY un3_s_fracto28_rnd_1_s_10_cZ(.LI(un3_s_fracto28_rnd_1_axb_10),.CI(un3_s_fracto28_rnd_1_cry_9),.O(un3_s_fracto28_rnd_1_s_10));
  MUXCY_L un3_s_fracto28_rnd_1_cry_10_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_9),.S(un3_s_fracto28_rnd_1_axb_10),.LO(un3_s_fracto28_rnd_1_cry_10));
  XORCY un3_s_fracto28_rnd_1_s_9_cZ(.LI(un3_s_fracto28_rnd_1_axb_9),.CI(un3_s_fracto28_rnd_1_cry_8),.O(un3_s_fracto28_rnd_1_s_9));
  MUXCY_L un3_s_fracto28_rnd_1_cry_9_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_8),.S(un3_s_fracto28_rnd_1_axb_9),.LO(un3_s_fracto28_rnd_1_cry_9));
  XORCY un3_s_fracto28_rnd_1_s_8_cZ(.LI(un3_s_fracto28_rnd_1_axb_8),.CI(un3_s_fracto28_rnd_1_cry_7),.O(un3_s_fracto28_rnd_1_s_8));
  MUXCY_L un3_s_fracto28_rnd_1_cry_8_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_7),.S(un3_s_fracto28_rnd_1_axb_8),.LO(un3_s_fracto28_rnd_1_cry_8));
  XORCY un3_s_fracto28_rnd_1_s_7_cZ(.LI(un3_s_fracto28_rnd_1_axb_7),.CI(un3_s_fracto28_rnd_1_cry_6),.O(un3_s_fracto28_rnd_1_s_7));
  MUXCY_L un3_s_fracto28_rnd_1_cry_7_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_6),.S(un3_s_fracto28_rnd_1_axb_7),.LO(un3_s_fracto28_rnd_1_cry_7));
  XORCY un3_s_fracto28_rnd_1_s_6_cZ(.LI(un3_s_fracto28_rnd_1_axb_6),.CI(un3_s_fracto28_rnd_1_cry_5),.O(un3_s_fracto28_rnd_1_s_6));
  MUXCY_L un3_s_fracto28_rnd_1_cry_6_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_5),.S(un3_s_fracto28_rnd_1_axb_6),.LO(un3_s_fracto28_rnd_1_cry_6));
  XORCY un3_s_fracto28_rnd_1_s_5_cZ(.LI(un3_s_fracto28_rnd_1_axb_5),.CI(un3_s_fracto28_rnd_1_cry_4),.O(un3_s_fracto28_rnd_1_s_5));
  MUXCY_L un3_s_fracto28_rnd_1_cry_5_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_4),.S(un3_s_fracto28_rnd_1_axb_5),.LO(un3_s_fracto28_rnd_1_cry_5));
  XORCY un3_s_fracto28_rnd_1_s_4_cZ(.LI(un3_s_fracto28_rnd_1_axb_4),.CI(un3_s_fracto28_rnd_1_cry_3),.O(un3_s_fracto28_rnd_1_s_4));
  MUXCY_L un3_s_fracto28_rnd_1_cry_4_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_3),.S(un3_s_fracto28_rnd_1_axb_4),.LO(un3_s_fracto28_rnd_1_cry_4));
  XORCY un3_s_fracto28_rnd_1_s_3_cZ(.LI(un3_s_fracto28_rnd_1_axb_3),.CI(un3_s_fracto28_rnd_1_cry_2),.O(un3_s_fracto28_rnd_1_s_3));
  MUXCY_L un3_s_fracto28_rnd_1_cry_3_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_2),.S(un3_s_fracto28_rnd_1_axb_3),.LO(un3_s_fracto28_rnd_1_cry_3));
  XORCY un3_s_fracto28_rnd_1_s_2_cZ(.LI(un3_s_fracto28_rnd_1_axb_2),.CI(un3_s_fracto28_rnd_1_cry_1),.O(un3_s_fracto28_rnd_1_s_2));
  MUXCY_L un3_s_fracto28_rnd_1_cry_2_cZ(.DI(GND),.CI(un3_s_fracto28_rnd_1_cry_1),.S(un3_s_fracto28_rnd_1_axb_2),.LO(un3_s_fracto28_rnd_1_cry_2));
  XORCY un3_s_fracto28_rnd_1_s_1_cZ(.LI(un3_s_fracto28_rnd_1_axb_1),.CI(s_fracto28_1[3:3]),.O(un3_s_fracto28_rnd_1_s_1));
  MUXCY_L un3_s_fracto28_rnd_1_cry_1_cZ(.DI(GND),.CI(s_fracto28_1[3:3]),.S(un3_s_fracto28_rnd_1_axb_1),.LO(un3_s_fracto28_rnd_1_cry_1));
  XORCY s_exp10_s_9(.LI(s_exp10_s_9_true),.CI(s_exp10_cry_8),.O(s_exp10[9:9]));
  XORCY s_exp10_s_8(.LI(s_exp10_5_ac0_13_i),.CI(s_exp10_cry_7),.O(s_exp10[8:8]));
  MUXCY_L s_exp10_cry_8_cZ(.DI(VCC),.CI(s_exp10_cry_7),.S(s_exp10_5_ac0_13_i),.LO(s_exp10_cry_8));
  XORCY s_exp10_s_7(.LI(s_exp10_5_i[7:7]),.CI(s_exp10_cry_6),.O(s_exp10[7:7]));
  MUXCY_L s_exp10_cry_7_cZ(.DI(VCC),.CI(s_exp10_cry_6),.S(s_exp10_5_i[7:7]),.LO(s_exp10_cry_7));
  XORCY s_exp10_s_6(.LI(s_exp10_5_i[6:6]),.CI(s_exp10_cry_5),.O(s_exp10[6:6]));
  MUXCY_L s_exp10_cry_6_cZ(.DI(VCC),.CI(s_exp10_cry_5),.S(s_exp10_5_i[6:6]),.LO(s_exp10_cry_6));
  XORCY s_exp10_s_5(.LI(s_exp10_5_i[5:5]),.CI(s_exp10_cry_4),.O(s_exp10[5:5]));
  MUXCY_L s_exp10_cry_5_cZ(.DI(VCC),.CI(s_exp10_cry_4),.S(s_exp10_5_i[5:5]),.LO(s_exp10_cry_5));
  XORCY s_exp10_s_4(.LI(s_exp10_axb_4),.CI(s_exp10_cry_3),.O(s_exp10[4:4]));
  MUXCY_L s_exp10_cry_4_cZ(.DI(s_exp10_5[4:4]),.CI(s_exp10_cry_3),.S(s_exp10_axb_4),.LO(s_exp10_cry_4));
  XORCY s_exp10_s_3(.LI(s_exp10_axb_3),.CI(s_exp10_cry_2),.O(s_exp10[3:3]));
  MUXCY_L s_exp10_cry_3_cZ(.DI(s_exp10_5[3:3]),.CI(s_exp10_cry_2),.S(s_exp10_axb_3),.LO(s_exp10_cry_3));
  XORCY s_exp10_s_2(.LI(s_exp10_axb_2),.CI(s_exp10_cry_1),.O(s_exp10[2:2]));
  MUXCY_L s_exp10_cry_2_cZ(.DI(s_exp10_5[2:2]),.CI(s_exp10_cry_1),.S(s_exp10_axb_2),.LO(s_exp10_cry_2));
  XORCY s_exp10_s_1(.LI(s_exp10_axb_1),.CI(s_exp10_cry_0),.O(s_exp10[1:1]));
  MUXCY_L s_exp10_cry_1_cZ(.DI(s_zeros_0_i_1_RNI027Q1[1:1]),.CI(s_exp10_cry_0),.S(s_exp10_axb_1),.LO(s_exp10_cry_1));
  MUXCY_L s_exp10_cry_0_cZ(.DI(s_exp10_5_axb0),.CI(GND),.S(s_exp10[0:0]),.LO(s_exp10_cry_0));
  FDR desc541(.Q(s_expo9_1[7:7]),.D(s_expo9_1_4[7:7]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc542(.Q(s_expo9_1[6:6]),.D(s_expo9_1_4[6:6]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc543(.Q(s_expo9_1[5:5]),.D(s_expo9_1_4[5:5]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc544(.Q(s_expo9_1[4:4]),.D(s_expo9_1_4[4:4]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc545(.Q(s_expo9_1[3:3]),.D(s_expo9_1_4[3:3]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc546(.Q(s_expo9_1[2:2]),.D(s_expo9_1_4[2:2]),.C(clk_i),.R(un12_s_exp10_iso));
  FDR desc547(.Q(s_expo9_1[1:1]),.D(s_expo9_1_4[1:1]),.C(clk_i),.R(un12_s_exp10_iso));
  FDS desc548(.Q(s_expo9_1[0:0]),.D(s_expo9_1_4[0:0]),.C(clk_i),.S(un12_s_exp10_iso));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT4 un2_s_overflow_o_i_o2_0_1_RNIMTS61_o6(.I0(N_835),.I1(s_output1[22:22]),.I2(s_output1[23:23]),.I3(N_91),.O(un2_s_qnan_o_0_a2_0_e));
defparam un2_s_overflow_o_i_o2_0_1_RNIMTS61_o6.INIT=16'h0080;
  LUT3 un2_s_overflow_o_i_o2_0_1_RNIMTS61_o5(.I0(s_output1[23:23]),.I1(N_91),.I2(s_ine_o),.O(N_6_i_0_e));
defparam un2_s_overflow_o_i_o2_0_1_RNIMTS61_o5.INIT=8'h20;
  LUT5 desc549(.I0(addsub_fract_o[7:7]),.I1(addsub_fract_o[9:9]),.I2(addsub_fract_o[8:8]),.I3(addsub_fract_o[10:10]),.I4(N_1869),.O(s_zeros_0_a2_0_2[3:3]));
defparam desc549.INIT=32'h00010000;
  LUT5 desc550(.I0(addsub_fract_o[7:7]),.I1(addsub_fract_o[9:9]),.I2(addsub_fract_o[8:8]),.I3(addsub_fract_o[10:10]),.I4(N_1869),.O(N_1872));
defparam desc550.INIT=32'h00000001;
  LUT2 desc551(.I0(s_rmode_i[0:0]),.I1(s_output1[22:22]),.O(N_811_1));
defparam desc551.INIT=4'h2;
  LUT2 desc552(.I0(N_811_4),.I1(s_output1[22:22]),.O(result_i_0_0));
defparam desc552.INIT=4'h2;
  LUT2 desc553(.I0(s_opb_i_15),.I1(s_opb_i_14),.O(result_2_10));
defparam desc553.INIT=4'hE;
  LUT3 desc554(.I0(s_opb_i_14),.I1(v_count_2_0[4:4]),.I2(N_54),.O(pre_norm_div_dvsor[5:5]));
defparam desc554.INIT=8'hB0;
  LUT5 un6_s_expo9_3_ac0_9_lut6_2_o6(.I0(s_expo9_1[5:5]),.I1(s_expo9_1[4:4]),.I2(s_fracto28_1[26:26]),.I3(s_fracto28_1[27:27]),.I4(un6_s_expo9_3_c4),.O(un6_s_expo9_3_c6));
defparam un6_s_expo9_3_ac0_9_lut6_2_o6.INIT=32'h88810000;
  LUT2 un6_s_expo9_3_ac0_9_lut6_2_o5(.I0(s_fracto28_1[26:26]),.I1(s_fracto28_1[27:27]),.O(un2_s_expo9_2));
defparam un6_s_expo9_3_ac0_9_lut6_2_o5.INIT=4'h1;
  LUT2 desc555(.I0(s_exp10[6:6]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[6:6]));
defparam desc555.INIT=4'hE;
  LUT2 desc556(.I0(s_exp10[7:7]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[7:7]));
defparam desc556.INIT=4'hE;
  LUT2 desc557(.I0(s_exp10[4:4]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[4:4]));
defparam desc557.INIT=4'hE;
  LUT2 desc558(.I0(s_exp10[5:5]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[5:5]));
defparam desc558.INIT=4'hE;
  LUT2 desc559(.I0(s_exp10[2:2]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[2:2]));
defparam desc559.INIT=4'hE;
  LUT2 desc560(.I0(s_exp10[3:3]),.I1(s_exp10[8:8]),.O(s_expo9_1_4[3:3]));
defparam desc560.INIT=4'hE;
  LUT2 desc561(.I0(addsub_fract_o[17:17]),.I1(addsub_fract_o[18:18]),.O(N_299_2));
defparam desc561.INIT=4'hE;
  LUT3 desc562(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[18:18]),.I2(s_shl1[0:0]),.O(N_1706));
defparam desc562.INIT=8'hCA;
  LUT3 desc563(.I0(addsub_fract_o[17:17]),.I1(addsub_fract_o[16:16]),.I2(s_shl1[0:0]),.O(N_1707));
defparam desc563.INIT=8'hCA;
  LUT3 desc564(.I0(addsub_fract_o[11:11]),.I1(addsub_fract_o[10:10]),.I2(s_shl1[0:0]),.O(N_1701));
defparam desc564.INIT=8'hCA;
  LUT3 desc565(.I0(addsub_fract_o[15:15]),.I1(addsub_fract_o[14:14]),.I2(s_shl1[0:0]),.O(N_1708));
defparam desc565.INIT=8'hCA;
  LUT3 desc566(.I0(addsub_fract_o[4:4]),.I1(addsub_fract_o[3:3]),.I2(s_shl1[0:0]),.O(N_1676));
defparam desc566.INIT=8'hCA;
  LUT2 desc567(.I0(addsub_fract_o[7:7]),.I1(addsub_fract_o[8:8]),.O(N_1774));
defparam desc567.INIT=4'h1;
  LUT3 desc568(.I0(addsub_fract_o[9:9]),.I1(addsub_fract_o[8:8]),.I2(s_shl1[0:0]),.O(N_1713));
defparam desc568.INIT=8'hCA;
  LUT3 desc569(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[24:24]),.I2(s_shl1[0:0]),.O(N_1842));
defparam desc569.INIT=8'h35;
  LUT3 desc570(.I0(addsub_fract_o[1:1]),.I1(addsub_fract_o[0:0]),.I2(s_shl1[0:0]),.O(N_1711));
defparam desc570.INIT=8'hCA;
  LUT3 desc571(.I0(addsub_fract_o[26:26]),.I1(addsub_fract_o[27:27]),.I2(s_shl1[0:0]),.O(N_1855));
defparam desc571.INIT=8'h53;
  LUT3 desc572(.I0(addsub_fract_o[2:2]),.I1(addsub_fract_o[3:3]),.I2(s_shl1[0:0]),.O(N_1712));
defparam desc572.INIT=8'hAC;
  LUT3 desc573(.I0(addsub_fract_o[6:6]),.I1(addsub_fract_o[7:7]),.I2(s_shl1[0:0]),.O(N_8));
defparam desc573.INIT=8'hAC;
  LUT3 desc574(.I0(addsub_fract_o[23:23]),.I1(addsub_fract_o[22:22]),.I2(s_shl1[0:0]),.O(N_1700));
defparam desc574.INIT=8'hCA;
  LUT4 desc575(.I0(addsub_fract_o[19:19]),.I1(addsub_fract_o[21:21]),.I2(addsub_fract_o[22:22]),.I3(addsub_fract_o[20:20]),.O(m149_e_1));
defparam desc575.INIT=16'h0001;
  LUT3 desc576(.I0(addsub_fract_o[21:21]),.I1(addsub_fract_o[20:20]),.I2(s_shl1[0:0]),.O(N_1705));
defparam desc576.INIT=8'hCA;
  LUT4 un3_s_underflow_o_0_a2_0_0_4_lut6_2_o6(.I0(s_output1[27:27]),.I1(s_output1[28:28]),.I2(s_output1[29:29]),.I3(s_output1[23:23]),.O(N_844_0_4));
defparam un3_s_underflow_o_0_a2_0_0_4_lut6_2_o6.INIT=16'h0001;
  LUT2 un3_s_underflow_o_0_a2_0_0_4_lut6_2_o5(.I0(s_output1[29:29]),.I1(s_output1[24:24]),.O(N_91_0_0_1));
defparam un3_s_underflow_o_0_a2_0_0_4_lut6_2_o5.INIT=4'h7;
  LUT4 desc577(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[6:6]),.I2(addsub_fract_o[4:4]),.I3(addsub_fract_o[3:3]),.O(N_1869));
defparam desc577.INIT=16'h0001;
  LUT3 desc578(.I0(addsub_fract_o[5:5]),.I1(addsub_fract_o[4:4]),.I2(s_shl1[0:0]),.O(N_6));
defparam desc578.INIT=8'hCA;
  LUT4 desc579(.I0(addsub_fract_o[11:11]),.I1(addsub_fract_o[13:13]),.I2(addsub_fract_o[12:12]),.I3(addsub_fract_o[14:14]),.O(N_289));
defparam desc579.INIT=16'hFFFE;
  LUT3 desc580(.I0(addsub_fract_o[13:13]),.I1(addsub_fract_o[12:12]),.I2(s_shl1[0:0]),.O(N_1709));
defparam desc580.INIT=8'hCA;
  LUT2 m133_lut6_2_o6(.I0(addsub_fract_o[26:26]),.I1(addsub_fract_o[27:27]),.O(N_1861));
defparam m133_lut6_2_o6.INIT=4'h1;
  LUT5 m133_lut6_2_o5(.I0(addsub_fract_o[25:25]),.I1(addsub_fract_o[26:26]),.I2(addsub_fract_o[23:23]),.I3(addsub_fract_o[24:24]),.I4(addsub_fract_o[27:27]),.O(m149_0));
defparam m133_lut6_2_o5.INIT=32'h00000001;
  LUT3 s_exp10_5_ac0_1_lut6_2_o6(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.I2(addsub_fract_o[27:27]),.O(s_exp10_5_c2));
defparam s_exp10_5_ac0_1_lut6_2_o6.INIT=8'hA8;
  LUT2 s_exp10_5_ac0_1_lut6_2_o5(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.O(result_1));
defparam s_exp10_5_ac0_1_lut6_2_o5.INIT=4'hE;
  LUT4 desc581(.I0(addsub_fract_o[0:0]),.I1(s_shl1[2:2]),.I2(s_shl1[1:1]),.I3(s_shl1[0:0]),.O(N_1776));
defparam desc581.INIT=16'h0002;
  LUT5 desc582(.I0(addsub_fract_o[1:1]),.I1(addsub_fract_o[0:0]),.I2(s_shl1[2:2]),.I3(s_shl1[1:1]),.I4(s_shl1[0:0]),.O(N_58));
defparam desc582.INIT=32'h000C000A;
  LUT5 desc583(.I0(addsub_fract_o[26:26]),.I1(addsub_fract_o[22:22]),.I2(addsub_fract_o[20:20]),.I3(addsub_fract_o[24:24]),.I4(addsub_fract_o[27:27]),.O(N_331));
defparam desc583.INIT=32'h00000001;
  LUT4 desc584(.I0(addsub_fract_o[26:26]),.I1(addsub_fract_o[22:22]),.I2(addsub_fract_o[24:24]),.I3(addsub_fract_o[27:27]),.O(N_329));
defparam desc584.INIT=16'h0001;
  LUT3 desc585(.I0(s_shl1[1:1]),.I1(N_1697),.I2(N_1686),.O(N_1727));
defparam desc585.INIT=8'hD8;
  LUT3 desc586(.I0(s_shl1[1:1]),.I1(N_1697),.I2(N_1696),.O(N_1726));
defparam desc586.INIT=8'hE4;
  LUT5 s_exp10_5_ac0_5_lut6_2_o6(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[3:3]),.I2(prenorm_addsub_exp_o[0:0]),.I3(prenorm_addsub_exp_o[2:2]),.I4(addsub_fract_o[27:27]),.O(s_exp10_5_c4));
defparam s_exp10_5_ac0_5_lut6_2_o6.INIT=32'h88008000;
  LUT4 s_exp10_5_ac0_5_lut6_2_o5(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.I2(prenorm_addsub_exp_o[2:2]),.I3(addsub_fract_o[27:27]),.O(s_exp10_5_c3));
defparam s_exp10_5_ac0_5_lut6_2_o5.INIT=16'hA080;
  LUT2 un2_s_overflow_o_i_o2_lut6_2_o6(.I0(s_output1[23:23]),.I1(N_91),.O(N_92));
defparam un2_s_overflow_o_i_o2_lut6_2_o6.INIT=4'hD;
  LUT5 un2_s_overflow_o_i_o2_lut6_2_o5(.I0(s_output1[23:23]),.I1(N_91),.I2(N_835),.I3(s_output1[22:22]),.I4(un3_s_snan_o_0),.O(N_9_i_0_e));
defparam un2_s_overflow_o_i_o2_lut6_2_o5.INIT=32'h00000222;
  LUT3 desc587(.I0(s_shl1[3:3]),.I1(N_1821),.I2(N_1822),.O(N_1823));
defparam desc587.INIT=8'hE4;
  LUT3 desc588(.I0(s_shl1[3:3]),.I1(N_1807),.I2(N_1808),.O(N_1809));
defparam desc588.INIT=8'hE4;
  LUT3 desc589(.I0(s_shl1[3:3]),.I1(N_1832),.I2(N_1803),.O(N_1833));
defparam desc589.INIT=8'hE4;
  LUT3 desc590(.I0(s_shl1[3:3]),.I1(N_1815),.I2(N_68),.O(N_1816));
defparam desc590.INIT=8'h4E;
  LUT3 s_exp10_5_axbxc1_lut6_2_o6(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.I2(addsub_fract_o[27:27]),.O(s_exp10_5[1:1]));
defparam s_exp10_5_axbxc1_lut6_2_o6.INIT=8'h56;
  LUT4 s_exp10_5_axbxc1_lut6_2_o5(.I0(prenorm_addsub_exp_o[1:1]),.I1(prenorm_addsub_exp_o[0:0]),.I2(s_zeros_0_i_1_RNI027Q1[1:1]),.I3(un1_s_exp10_3),.O(N_389));
defparam s_exp10_5_axbxc1_lut6_2_o5.INIT=16'h0F99;
  LUT3 desc591(.I0(un4_s_infa),.I1(un1_s_infb),.I2(div_zero_o_0),.O(N_84));
defparam desc591.INIT=8'hFE;
  LUT4 desc592(.I0(un4_s_infa),.I1(un1_s_infb),.I2(s_output_o_m0[25:25]),.I3(s_overflow),.O(s_output_o_0_e[25:25]));
defparam desc592.INIT=16'hFFFE;
  LUT3 s_output_os2_i_a5_lut6_2_o6(.I0(un4_s_infa),.I1(un1_s_infb),.I2(s_overflow),.O(N_2203));
defparam s_output_os2_i_a5_lut6_2_o6.INIT=8'h01;
  LUT5 s_output_os2_i_a5_lut6_2_o5(.I0(un4_s_infa),.I1(un1_s_infb),.I2(s_overflow),.I3(s_expo9_3[6:6]),.I4(un15_s_zero_fract_sn),.O(s_output_o_0_e[29:29]));
defparam s_output_os2_i_a5_lut6_2_o5.INIT=32'hFEFEFFFE;
  LUT4 desc593(.I0(un4_s_infa),.I1(un1_s_infb),.I2(un15_s_zero_fract_sn),.I3(s_overflow),.O(N_473_i));
defparam desc593.INIT=16'hFFFE;
  LUT5 desc594(.I0(s_expo9_3[3:3]),.I1(un4_s_infa),.I2(un1_s_infb),.I3(un15_s_zero_fract_sn),.I4(s_overflow),.O(s_output_o_0_e[26:26]));
defparam desc594.INIT=32'hFFFFFCFE;
endmodule
module pre_norm_mul_inj (v_count,s_fracta_52_o_0_e,pre_norm_mul_exp_10,s_exp_10_o_1,s_exp_10_o_0_d0,s_exp_10_o_0_0,s_exp_10_o_0_1,s_opb_i,s_opa_i,un4_s_expb_in_2_i_o2_0,N_48_0,N_1245,clk_i,un4_s_expb_in_2_i_o2_1,N_1077,result_i_o3_lut6_2_O6,N_1084_i,p_desc595_p_O_FD,p_desc596_p_O_FD,p_desc597_p_O_FD,p_desc598_p_O_FD,p_desc599_p_O_FD,p_desc600_p_O_FD,p_desc601_p_O_FD,p_desc602_p_O_FD,p_desc603_p_O_FD,p_desc604_p_O_FD);
input [4:4] v_count ;
output [29:29] s_fracta_52_o_0_e ;
output [9:0] pre_norm_mul_exp_10 ;
input s_exp_10_o_1 ;
input s_exp_10_o_0_d0 ;
output s_exp_10_o_0_0 ;
output s_exp_10_o_0_1 ;
input [30:23] s_opb_i ;
input [30:23] s_opa_i ;
output un4_s_expb_in_2_i_o2_0 ;
input N_48_0 ;
input N_1245 ;
input clk_i ;
input un4_s_expb_in_2_i_o2_1 ;
input N_1077 ;
input result_i_o3_lut6_2_O6 ;
input N_1084_i ;
wire s_exp_10_o_1 ;
wire s_exp_10_o_0_d0 ;
wire s_exp_10_o_0_0 ;
wire s_exp_10_o_0_1 ;
wire un4_s_expb_in_2_i_o2_0 ;
wire N_48_0 ;
wire N_1245 ;
wire clk_i ;
wire un4_s_expb_in_2_i_o2_1 ;
wire N_1077 ;
wire result_i_o3_lut6_2_O6 ;
wire N_1084_i ;
wire [9:2] s_exp_10_o_0 ;
wire [9:2] s_exp_10_o ;
wire [23:23] s_opa_i_0 ;
wire s_exp_10_o_c5 ;
wire VCC ;
wire GND ;
wire s_exp_10_o_6_c4 ;
wire s_exp_10_o_0_axb_0 ;
wire s_exp_10_o_0_axb_1 ;
wire s_exp_10_o_0_axb_2 ;
wire s_exp_10_o_0_axb_5 ;
wire s_exp_10_o_0_cry_0_RNO ;
wire s_exp_10_o_0_cry_0_cy ;
wire s_exp_10_o_0_axb_4 ;
wire s_exp_10_o_0_axb_3 ;
wire s_exp_10_o_0_axb_6 ;
wire s_exp_10_o_0_axb_7 ;
wire s_exp_10_o_0_axb_9 ;
wire s_exp_10_o_0_axb_8 ;
wire s_exp_10_o_0_cry_8 ;
wire s_exp_10_o_0_cry_7 ;
wire s_exp_10_o_0_cry_6 ;
wire s_exp_10_o_0_cry_5 ;
wire s_exp_10_o_0_cry_4 ;
wire s_exp_10_o_0_cry_3 ;
wire s_exp_10_o_0_cry_2 ;
wire s_exp_10_o_0_cry_1 ;
wire s_exp_10_o_0_cry_0 ;
input p_desc595_p_O_FD ;
input p_desc596_p_O_FD ;
input p_desc597_p_O_FD ;
input p_desc598_p_O_FD ;
input p_desc599_p_O_FD ;
input p_desc600_p_O_FD ;
input p_desc601_p_O_FD ;
input p_desc602_p_O_FD ;
input p_desc603_p_O_FD ;
input p_desc604_p_O_FD ;
// instances
  LUT3 s_exp_10_o_0_axb_1_cZ(.I0(s_opa_i[24:24]),.I1(s_opb_i[23:23]),.I2(s_opb_i[24:24]),.O(s_exp_10_o_0_axb_1));
defparam s_exp_10_o_0_axb_1_cZ.INIT=8'h96;
  LUT4 s_exp_10_o_0_axb_2_cZ(.I0(s_opa_i[25:25]),.I1(s_opb_i[23:23]),.I2(s_opb_i[24:24]),.I3(s_opb_i[25:25]),.O(s_exp_10_o_0_axb_2));
defparam s_exp_10_o_0_axb_2_cZ.INIT=16'h956A;
  LUT4 s_exp_10_o_0_axb_5_cZ(.I0(s_exp_10_o_6_c4),.I1(s_opa_i[28:28]),.I2(s_opb_i[27:27]),.I3(s_opb_i[28:28]),.O(s_exp_10_o_0_axb_5));
defparam s_exp_10_o_0_axb_5_cZ.INIT=16'h936C;
  LUT1 s_exp_10_o_0_cry_0_thru(.I0(s_opa_i[23:23]),.O(s_opa_i_0[23:23]));
defparam s_exp_10_o_0_cry_0_thru.INIT=2'h2;
  p_O_FD desc595(.Q(pre_norm_mul_exp_10[1:1]),.D(s_exp_10_o_1),.C(clk_i),.E(p_desc595_p_O_FD));
  p_O_FD desc596(.Q(pre_norm_mul_exp_10[2:2]),.D(s_exp_10_o[2:2]),.C(clk_i),.E(p_desc596_p_O_FD));
  p_O_FD desc597(.Q(pre_norm_mul_exp_10[3:3]),.D(s_exp_10_o[3:3]),.C(clk_i),.E(p_desc597_p_O_FD));
  p_O_FD desc598(.Q(pre_norm_mul_exp_10[4:4]),.D(s_exp_10_o[4:4]),.C(clk_i),.E(p_desc598_p_O_FD));
  p_O_FD desc599(.Q(pre_norm_mul_exp_10[5:5]),.D(s_exp_10_o[5:5]),.C(clk_i),.E(p_desc599_p_O_FD));
  p_O_FD desc600(.Q(pre_norm_mul_exp_10[6:6]),.D(s_exp_10_o[6:6]),.C(clk_i),.E(p_desc600_p_O_FD));
  p_O_FD desc601(.Q(pre_norm_mul_exp_10[7:7]),.D(s_exp_10_o[7:7]),.C(clk_i),.E(p_desc601_p_O_FD));
  p_O_FD desc602(.Q(pre_norm_mul_exp_10[8:8]),.D(s_exp_10_o[8:8]),.C(clk_i),.E(p_desc602_p_O_FD));
  p_O_FD desc603(.Q(pre_norm_mul_exp_10[9:9]),.D(s_exp_10_o[9:9]),.C(clk_i),.E(p_desc603_p_O_FD));
  p_O_FD desc604(.Q(pre_norm_mul_exp_10[0:0]),.D(s_exp_10_o_0_d0),.C(clk_i),.E(p_desc604_p_O_FD));
  LUT6 s_exp_10_o_0_cry_0_RNO_cZ(.I0(s_opb_i[24:24]),.I1(s_opb_i[28:28]),.I2(s_opb_i[27:27]),.I3(s_opb_i[23:23]),.I4(un4_s_expb_in_2_i_o2_0),.I5(un4_s_expb_in_2_i_o2_1),.O(s_exp_10_o_0_cry_0_RNO));
defparam s_exp_10_o_0_cry_0_RNO_cZ.INIT=64'h00FF00FF00FF00FE;
  MUXCY_L s_exp_10_o_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(s_opa_i_0[23:23]),.LO(s_exp_10_o_0_cry_0_cy));
  LUT6 s_exp_10_o_0_s_0_lut6_2_RNO(.I0(s_opb_i[24:24]),.I1(s_opb_i[28:28]),.I2(s_opb_i[27:27]),.I3(s_opb_i[23:23]),.I4(un4_s_expb_in_2_i_o2_0),.I5(un4_s_expb_in_2_i_o2_1),.O(s_exp_10_o_0_axb_0));
defparam s_exp_10_o_0_s_0_lut6_2_RNO.INIT=64'h00FF00FF00FF00FE;
  LUT6 s_exp_10_o_0_axb_4_cZ(.I0(s_opb_i[25:25]),.I1(s_opa_i[27:27]),.I2(s_opb_i[26:26]),.I3(s_opb_i[24:24]),.I4(s_opb_i[27:27]),.I5(s_opb_i[23:23]),.O(s_exp_10_o_0_axb_4));
defparam s_exp_10_o_0_axb_4_cZ.INIT=64'h93336CCC3333CCCC;
  LUT6_L s_exp_10_o_axbxc3(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_exp_10_o_0_0),.I3(s_exp_10_o_0[3:3]),.I4(s_exp_10_o_0_1),.I5(s_exp_10_o_0[2:2]),.LO(s_exp_10_o[3:3]));
defparam s_exp_10_o_axbxc3.INIT=64'hEF10FF00FF00FF00;
  LUT5_L s_exp_10_o_axbxc2(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_exp_10_o_0_0),.I3(s_exp_10_o_0_1),.I4(s_exp_10_o_0[2:2]),.LO(s_exp_10_o[2:2]));
defparam s_exp_10_o_axbxc2.INIT=32'hEFFF1000;
  LUT5 s_exp_10_o_0_axb_3_cZ(.I0(s_opb_i[25:25]),.I1(s_opa_i[26:26]),.I2(s_opb_i[26:26]),.I3(s_opb_i[24:24]),.I4(s_opb_i[23:23]),.O(s_exp_10_o_0_axb_3));
defparam s_exp_10_o_0_axb_3_cZ.INIT=32'h963C3C3C;
  LUT5 s_exp_10_o_0_axb_6_cZ(.I0(s_opa_i[29:29]),.I1(s_opb_i[29:29]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.I4(s_exp_10_o_6_c4),.O(s_exp_10_o_0_axb_6));
defparam s_exp_10_o_0_axb_6_cZ.INIT=32'h96666666;
  LUT6 s_exp_10_o_0_axb_7_cZ(.I0(s_opb_i[30:30]),.I1(s_opa_i[30:30]),.I2(s_opb_i[29:29]),.I3(s_opb_i[28:28]),.I4(s_opb_i[27:27]),.I5(s_exp_10_o_6_c4),.O(s_exp_10_o_0_axb_7));
defparam s_exp_10_o_0_axb_7_cZ.INIT=64'h6999999999999999;
  LUT6 s_exp_10_o_ac0_7(.I0(s_exp_10_o_0_0),.I1(result_i_o3_lut6_2_O6),.I2(s_exp_10_o_0[4:4]),.I3(s_exp_10_o_0[3:3]),.I4(s_exp_10_o_0_1),.I5(s_exp_10_o_0[2:2]),.O(s_exp_10_o_c5));
defparam s_exp_10_o_ac0_7.INIT=64'h2000000000000000;
  LUT6_L s_exp_10_o_axbxc4(.I0(s_exp_10_o_0_0),.I1(result_i_o3_lut6_2_O6),.I2(s_exp_10_o_0[4:4]),.I3(s_exp_10_o_0[3:3]),.I4(s_exp_10_o_0_1),.I5(s_exp_10_o_0[2:2]),.LO(s_exp_10_o[4:4]));
defparam s_exp_10_o_axbxc4.INIT=64'hD2F0F0F0F0F0F0F0;
  LUT5 s_exp_10_o_0_axb_9_cZ(.I0(s_opb_i[30:30]),.I1(s_opb_i[29:29]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.I4(s_exp_10_o_6_c4),.O(s_exp_10_o_0_axb_9));
defparam s_exp_10_o_0_axb_9_cZ.INIT=32'h15555555;
  LUT5 s_exp_10_o_0_axb_8_cZ(.I0(s_opb_i[30:30]),.I1(s_opb_i[29:29]),.I2(s_opb_i[28:28]),.I3(s_opb_i[27:27]),.I4(s_exp_10_o_6_c4),.O(s_exp_10_o_0_axb_8));
defparam s_exp_10_o_0_axb_8_cZ.INIT=32'h15555555;
  LUT6_L s_exp_10_o_axbxc9(.I0(s_exp_10_o_0[9:9]),.I1(s_exp_10_o_0[8:8]),.I2(s_exp_10_o_0[7:7]),.I3(s_exp_10_o_0[5:5]),.I4(s_exp_10_o_0[6:6]),.I5(s_exp_10_o_c5),.LO(s_exp_10_o[9:9]));
defparam s_exp_10_o_axbxc9.INIT=64'h6AAAAAAAAAAAAAAA;
  XORCY s_exp_10_o_0_s_9(.LI(s_exp_10_o_0_axb_9),.CI(s_exp_10_o_0_cry_8),.O(s_exp_10_o_0[9:9]));
  XORCY s_exp_10_o_0_s_8(.LI(s_exp_10_o_0_axb_8),.CI(s_exp_10_o_0_cry_7),.O(s_exp_10_o_0[8:8]));
  MUXCY_L s_exp_10_o_0_cry_8_cZ(.DI(GND),.CI(s_exp_10_o_0_cry_7),.S(s_exp_10_o_0_axb_8),.LO(s_exp_10_o_0_cry_8));
  XORCY s_exp_10_o_0_s_7(.LI(s_exp_10_o_0_axb_7),.CI(s_exp_10_o_0_cry_6),.O(s_exp_10_o_0[7:7]));
  MUXCY_L s_exp_10_o_0_cry_7_cZ(.DI(s_opa_i[30:30]),.CI(s_exp_10_o_0_cry_6),.S(s_exp_10_o_0_axb_7),.LO(s_exp_10_o_0_cry_7));
  XORCY s_exp_10_o_0_s_6(.LI(s_exp_10_o_0_axb_6),.CI(s_exp_10_o_0_cry_5),.O(s_exp_10_o_0[6:6]));
  MUXCY_L s_exp_10_o_0_cry_6_cZ(.DI(s_opa_i[29:29]),.CI(s_exp_10_o_0_cry_5),.S(s_exp_10_o_0_axb_6),.LO(s_exp_10_o_0_cry_6));
  XORCY s_exp_10_o_0_s_5(.LI(s_exp_10_o_0_axb_5),.CI(s_exp_10_o_0_cry_4),.O(s_exp_10_o_0[5:5]));
  MUXCY_L s_exp_10_o_0_cry_5_cZ(.DI(s_opa_i[28:28]),.CI(s_exp_10_o_0_cry_4),.S(s_exp_10_o_0_axb_5),.LO(s_exp_10_o_0_cry_5));
  XORCY s_exp_10_o_0_s_4(.LI(s_exp_10_o_0_axb_4),.CI(s_exp_10_o_0_cry_3),.O(s_exp_10_o_0[4:4]));
  MUXCY_L s_exp_10_o_0_cry_4_cZ(.DI(s_opa_i[27:27]),.CI(s_exp_10_o_0_cry_3),.S(s_exp_10_o_0_axb_4),.LO(s_exp_10_o_0_cry_4));
  XORCY s_exp_10_o_0_s_3(.LI(s_exp_10_o_0_axb_3),.CI(s_exp_10_o_0_cry_2),.O(s_exp_10_o_0[3:3]));
  MUXCY_L s_exp_10_o_0_cry_3_cZ(.DI(s_opa_i[26:26]),.CI(s_exp_10_o_0_cry_2),.S(s_exp_10_o_0_axb_3),.LO(s_exp_10_o_0_cry_3));
  XORCY s_exp_10_o_0_s_2(.LI(s_exp_10_o_0_axb_2),.CI(s_exp_10_o_0_cry_1),.O(s_exp_10_o_0[2:2]));
  MUXCY_L s_exp_10_o_0_cry_2_cZ(.DI(s_opa_i[25:25]),.CI(s_exp_10_o_0_cry_1),.S(s_exp_10_o_0_axb_2),.LO(s_exp_10_o_0_cry_2));
  XORCY s_exp_10_o_0_s_1(.LI(s_exp_10_o_0_axb_1),.CI(s_exp_10_o_0_cry_0),.O(s_exp_10_o_0_1));
  MUXCY_L s_exp_10_o_0_cry_1_cZ(.DI(s_opa_i[24:24]),.CI(s_exp_10_o_0_cry_0),.S(s_exp_10_o_0_axb_1),.LO(s_exp_10_o_0_cry_1));
  MUXCY_L s_exp_10_o_0_cry_0_cZ(.DI(N_1084_i),.CI(s_exp_10_o_0_cry_0_cy),.S(s_exp_10_o_0_cry_0_RNO),.LO(s_exp_10_o_0_cry_0));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT2 s_exp_10_o_0_s_0_lut6_2_o6(.I0(s_opa_i[23:23]),.I1(s_exp_10_o_0_axb_0),.O(s_exp_10_o_0_0));
defparam s_exp_10_o_0_s_0_lut6_2_o6.INIT=4'h6;
  LUT4 s_exp_10_o_0_s_0_lut6_2_o5(.I0(N_48_0),.I1(N_1245),.I2(v_count[4:4]),.I3(s_opa_i[23:23]),.O(s_fracta_52_o_0_e[29:29]));
defparam s_exp_10_o_0_s_0_lut6_2_o5.INIT=16'h0A0C;
  LUT4 s_exp_10_o_6_ac0_5_lut6_2_o6(.I0(s_opb_i[25:25]),.I1(s_opb_i[26:26]),.I2(s_opb_i[24:24]),.I3(s_opb_i[23:23]),.O(s_exp_10_o_6_c4));
defparam s_exp_10_o_6_ac0_5_lut6_2_o6.INIT=16'h8000;
  LUT2 s_exp_10_o_6_ac0_5_lut6_2_o5(.I0(s_opb_i[30:30]),.I1(s_opb_i[25:25]),.O(un4_s_expb_in_2_i_o2_0));
defparam s_exp_10_o_6_ac0_5_lut6_2_o5.INIT=4'hE;
  LUT4 s_exp_10_o_axbxc7_lut6_2_o6(.I0(s_exp_10_o_0[7:7]),.I1(s_exp_10_o_0[5:5]),.I2(s_exp_10_o_0[6:6]),.I3(s_exp_10_o_c5),.O(s_exp_10_o[7:7]));
defparam s_exp_10_o_axbxc7_lut6_2_o6.INIT=16'h6AAA;
  LUT2 s_exp_10_o_axbxc7_lut6_2_o5(.I0(s_exp_10_o_0[5:5]),.I1(s_exp_10_o_c5),.O(s_exp_10_o[5:5]));
defparam s_exp_10_o_axbxc7_lut6_2_o5.INIT=4'h6;
  LUT5 s_exp_10_o_axbxc8_lut6_2_o6(.I0(s_exp_10_o_0[8:8]),.I1(s_exp_10_o_0[7:7]),.I2(s_exp_10_o_0[5:5]),.I3(s_exp_10_o_0[6:6]),.I4(s_exp_10_o_c5),.O(s_exp_10_o[8:8]));
defparam s_exp_10_o_axbxc8_lut6_2_o6.INIT=32'h6AAAAAAA;
  LUT3 s_exp_10_o_axbxc8_lut6_2_o5(.I0(s_exp_10_o_0[5:5]),.I1(s_exp_10_o_0[6:6]),.I2(s_exp_10_o_c5),.O(s_exp_10_o[6:6]));
defparam s_exp_10_o_axbxc8_lut6_2_o5.INIT=8'h6C;
endmodule
module mul_24_inj (s_fractb_i_11,s_fractb_i_8,s_fractb_i_20,s_fractb_i_10,s_fractb_i_9,s_fractb_i_22,s_fractb_i_21,s_fractb_i_7,s_fractb_i_6,s_fractb_i_19,s_fractb_i_18,s_fractb_i_5,s_fractb_i_4,s_fractb_i_17,s_fractb_i_16,s_fractb_i_3,s_fractb_i_15,s_fractb_i_2,s_fractb_i_14,s_fractb_i_1,s_fractb_i_13,s_fractb_i_0,s_fractb_i_12,s_fracta_i,s_opb_i_31,s_opb_i_11,s_opb_i_10,s_opb_i_22,s_opb_i_9,s_opb_i_21,s_opb_i_8,s_opb_i_20,s_opb_i_7,s_opb_i_19,s_opb_i_6,s_opb_i_18,s_opb_i_5,s_opb_i_17,s_opb_i_4,s_opb_i_16,s_opb_i_3,s_opb_i_15,s_opb_i_2,s_opb_i_14,s_opb_i_1,s_opb_i_13,s_opb_i_0,s_opb_i_12,s_opa_i_31,s_opa_i_11,s_opa_i_10,s_opa_i_22,s_opa_i_9,s_opa_i_21,s_opa_i_8,s_opa_i_20,s_opa_i_7,s_opa_i_19,s_opa_i_6,s_opa_i_18,s_opa_i_5,s_opa_i_17,s_opa_i_4,s_opa_i_16,s_opa_i_3,s_opa_i_15,s_opa_i_2,s_opa_i_14,s_opa_i_1,s_opa_i_13,s_opa_i_0,s_opa_i_12,mul_24_fract_48,opa_i,opb_i,clk_i,s_start_i,result_1_i_o3_0_e,s_signa_i,s_signb_i,result_i_o3_lut6_2_O6);
output s_fractb_i_11 ;
output s_fractb_i_8 ;
output s_fractb_i_20 ;
output s_fractb_i_10 ;
output s_fractb_i_9 ;
output s_fractb_i_22 ;
output s_fractb_i_21 ;
output s_fractb_i_7 ;
output s_fractb_i_6 ;
output s_fractb_i_19 ;
output s_fractb_i_18 ;
output s_fractb_i_5 ;
output s_fractb_i_4 ;
output s_fractb_i_17 ;
output s_fractb_i_16 ;
output s_fractb_i_3 ;
output s_fractb_i_15 ;
output s_fractb_i_2 ;
output s_fractb_i_14 ;
output s_fractb_i_1 ;
output s_fractb_i_13 ;
output s_fractb_i_0 ;
output s_fractb_i_12 ;
output [22:0] s_fracta_i ;
input s_opb_i_31 ;
input s_opb_i_11 ;
input s_opb_i_10 ;
input s_opb_i_22 ;
input s_opb_i_9 ;
input s_opb_i_21 ;
input s_opb_i_8 ;
input s_opb_i_20 ;
input s_opb_i_7 ;
input s_opb_i_19 ;
input s_opb_i_6 ;
input s_opb_i_18 ;
input s_opb_i_5 ;
input s_opb_i_17 ;
input s_opb_i_4 ;
input s_opb_i_16 ;
input s_opb_i_3 ;
input s_opb_i_15 ;
input s_opb_i_2 ;
input s_opb_i_14 ;
input s_opb_i_1 ;
input s_opb_i_13 ;
input s_opb_i_0 ;
input s_opb_i_12 ;
input s_opa_i_31 ;
input s_opa_i_11 ;
input s_opa_i_10 ;
input s_opa_i_22 ;
input s_opa_i_9 ;
input s_opa_i_21 ;
input s_opa_i_8 ;
input s_opa_i_20 ;
input s_opa_i_7 ;
input s_opa_i_19 ;
input s_opa_i_6 ;
input s_opa_i_18 ;
input s_opa_i_5 ;
input s_opa_i_17 ;
input s_opa_i_4 ;
input s_opa_i_16 ;
input s_opa_i_3 ;
input s_opa_i_15 ;
input s_opa_i_2 ;
input s_opa_i_14 ;
input s_opa_i_1 ;
input s_opa_i_13 ;
input s_opa_i_0 ;
input s_opa_i_12 ;
output [47:0] mul_24_fract_48 ;
input [17:12] opa_i ;
input [17:12] opb_i ;
input clk_i ;
input s_start_i ;
input result_1_i_o3_0_e ;
output s_signa_i ;
output s_signb_i ;
input result_i_o3_lut6_2_O6 ;
wire s_fractb_i_11 ;
wire s_fractb_i_8 ;
wire s_fractb_i_20 ;
wire s_fractb_i_10 ;
wire s_fractb_i_9 ;
wire s_fractb_i_22 ;
wire s_fractb_i_21 ;
wire s_fractb_i_7 ;
wire s_fractb_i_6 ;
wire s_fractb_i_19 ;
wire s_fractb_i_18 ;
wire s_fractb_i_5 ;
wire s_fractb_i_4 ;
wire s_fractb_i_17 ;
wire s_fractb_i_16 ;
wire s_fractb_i_3 ;
wire s_fractb_i_15 ;
wire s_fractb_i_2 ;
wire s_fractb_i_14 ;
wire s_fractb_i_1 ;
wire s_fractb_i_13 ;
wire s_fractb_i_0 ;
wire s_fractb_i_12 ;
wire s_opb_i_31 ;
wire s_opb_i_11 ;
wire s_opb_i_10 ;
wire s_opb_i_22 ;
wire s_opb_i_9 ;
wire s_opb_i_21 ;
wire s_opb_i_8 ;
wire s_opb_i_20 ;
wire s_opb_i_7 ;
wire s_opb_i_19 ;
wire s_opb_i_6 ;
wire s_opb_i_18 ;
wire s_opb_i_5 ;
wire s_opb_i_17 ;
wire s_opb_i_4 ;
wire s_opb_i_16 ;
wire s_opb_i_3 ;
wire s_opb_i_15 ;
wire s_opb_i_2 ;
wire s_opb_i_14 ;
wire s_opb_i_1 ;
wire s_opb_i_13 ;
wire s_opb_i_0 ;
wire s_opb_i_12 ;
wire s_opa_i_31 ;
wire s_opa_i_11 ;
wire s_opa_i_10 ;
wire s_opa_i_22 ;
wire s_opa_i_9 ;
wire s_opa_i_21 ;
wire s_opa_i_8 ;
wire s_opa_i_20 ;
wire s_opa_i_7 ;
wire s_opa_i_19 ;
wire s_opa_i_6 ;
wire s_opa_i_18 ;
wire s_opa_i_5 ;
wire s_opa_i_17 ;
wire s_opa_i_4 ;
wire s_opa_i_16 ;
wire s_opa_i_3 ;
wire s_opa_i_15 ;
wire s_opa_i_2 ;
wire s_opa_i_14 ;
wire s_opa_i_1 ;
wire s_opa_i_13 ;
wire s_opa_i_0 ;
wire s_opa_i_12 ;
wire clk_i ;
wire s_start_i ;
wire result_1_i_o3_0_e ;
wire s_signa_i ;
wire s_signb_i ;
wire result_i_o3_lut6_2_O6 ;
wire [2:0] count ;
wire s_state ;
wire [2:2] count_RNILIBD_O5 ;
wire [2:2] count_RNILIBD_2_O5 ;
wire [23:23] s_fractb_i ;
wire [47:30] un8_prod2 ;
wire [2:2] count_RNILIBD_0_O5 ;
wire [2:2] count_RNILIBD_1_O6 ;
wire [23:0] sum_0 ;
wire [670:653] un54_sum ;
wire [23:0] sum_1 ;
wire [23:0] sum_2 ;
wire [23:12] sum_3 ;
wire [23:12] prod2_2_0 ;
wire [11:0] un23_prod2 ;
wire [23:12] prod2_0_0 ;
wire [23:12] prod2_1_0 ;
wire [23:12] prod2_3_0 ;
wire [17:6] prod2_0_1 ;
wire [11:0] un92_prod2 ;
wire [17:6] prod2_1_1 ;
wire [17:6] prod2_2_1 ;
wire [17:6] prod2_3_1 ;
wire [17:6] prod2_0_2 ;
wire [11:0] un139_prod2 ;
wire [17:6] prod2_1_2 ;
wire [17:6] prod2_2_2 ;
wire [17:6] prod2_3_2 ;
wire [11:0] prod2_0_3 ;
wire [11:0] un184_prod2 ;
wire [11:0] prod2_1_3 ;
wire [11:0] prod2_2_3 ;
wire [11:0] prod2_3_3 ;
wire [29:0] ACOUT ;
wire [17:0] BCOUT ;
wire [3:0] CARRYOUT ;
wire [47:12] P_uc ;
wire [47:0] PCOUT ;
wire [29:0] ACOUT_0 ;
wire [17:0] BCOUT_0 ;
wire [3:0] CARRYOUT_0 ;
wire [47:12] P_uc_0 ;
wire [47:0] PCOUT_0 ;
wire [29:0] ACOUT_1 ;
wire [17:0] BCOUT_1 ;
wire [3:0] CARRYOUT_1 ;
wire [47:12] P_uc_1 ;
wire [47:0] PCOUT_1 ;
wire [29:0] ACOUT_2 ;
wire [17:0] BCOUT_2 ;
wire [3:0] CARRYOUT_2 ;
wire [47:12] P_uc_2 ;
wire [47:0] PCOUT_2 ;
wire VCC ;
wire N_246 ;
wire un2_i ;
wire GND ;
wire N_235_mux ;
wire N_2719 ;
wire N_124_0_i ;
wire prod2_3_0_1_sqmuxa ;
wire m39 ;
wire prod2_1_0_1_sqmuxa ;
wire N_2731_i_0_0 ;
wire N_1409 ;
wire prod2_2_0_1_sqmuxa ;
wire N_1411 ;
wire N_1410 ;
wire N_248 ;
wire N_1408 ;
wire N_85_0 ;
wire N_142_0 ;
wire N_145_0_i ;
wire N_3283 ;
wire un54_sum_axb_11 ;
wire N_103_0_i ;
wire N_100_0_i ;
wire N_97_0_i ;
wire N_94_0_i ;
wire N_91_0_i ;
wire N_88_0_i ;
wire un36_prod_a_b_axb_19 ;
wire un36_prod_a_b_axb_18 ;
wire un36_prod_a_b_axb_16 ;
wire un36_prod_a_b_axb_13 ;
wire un36_prod_a_b_axb_12 ;
wire un36_prod_a_b_axb_10 ;
wire un36_prod_a_b_axb_6 ;
wire un36_prod_a_b_axb_4 ;
wire un36_prod_a_b_axb_22 ;
wire un36_prod_a_b_axb_20 ;
wire un36_prod_a_b_axb_11 ;
wire un36_prod_a_b_axb_17 ;
wire un36_prod_a_b_axb_5 ;
wire un36_prod_a_b_axb_14 ;
wire N_136_0 ;
wire N_139_0 ;
wire N_3281 ;
wire N_3282 ;
wire N_3293 ;
wire N_3294 ;
wire un54_sum_axb_9 ;
wire N_130_0 ;
wire N_133_0 ;
wire N_3279 ;
wire N_3280 ;
wire N_3291 ;
wire N_3292 ;
wire un54_sum_axb_7 ;
wire un36_prod_a_b_axb_9 ;
wire un36_prod_a_b_axb_8 ;
wire N_127_0 ;
wire N_3278 ;
wire N_3290 ;
wire un54_sum_axb_6 ;
wire un54_sum_axb_8 ;
wire un54_sum_axb_10 ;
wire un36_prod_a_b_axb_21 ;
wire un36_prod_a_b_axb_15 ;
wire N_118_0 ;
wire N_121_0 ;
wire N_3276 ;
wire N_3277 ;
wire N_3288 ;
wire N_3289 ;
wire un54_sum_axb_4 ;
wire N_112_0 ;
wire N_115_0 ;
wire N_172_0 ;
wire N_3274 ;
wire N_3286 ;
wire N_3287 ;
wire un54_sum_axb_2 ;
wire un36_prod_a_b_axb_3 ;
wire un36_prod_a_b_axb_2 ;
wire un36_prod_a_b_axb_1 ;
wire N_106_0 ;
wire N_3272 ;
wire N_3284 ;
wire N_109_0 ;
wire N_3273 ;
wire N_3285 ;
wire un36_prod_a_b_axb_7 ;
wire un54_sum_axb_1 ;
wire un54_sum_axb_5 ;
wire un54_sum_axb_3 ;
wire un36_prod_a_b_axb_34 ;
wire un36_prod_a_b_axb_33 ;
wire un36_prod_a_b_axb_32 ;
wire un36_prod_a_b_axb_31 ;
wire un36_prod_a_b_axb_30 ;
wire un36_prod_a_b_axb_29 ;
wire un36_prod_a_b_axb_28 ;
wire un36_prod_a_b_axb_27 ;
wire un36_prod_a_b_axb_26 ;
wire un36_prod_a_b_axb_25 ;
wire un36_prod_a_b_axb_24 ;
wire un54_sum_axb_16 ;
wire un54_sum_axb_15 ;
wire un54_sum_axb_14 ;
wire un54_sum_axb_13 ;
wire un54_sum_axb_12 ;
wire un36_prod_a_b_axb_23 ;
wire un36_prod_a_b_cry_0_RNO ;
wire un36_prod_a_b_cry_1_RNO ;
wire un36_prod_a_b_cry_2_RNO ;
wire un36_prod_a_b_cry_3_RNO ;
wire un36_prod_a_b_cry_4_RNO ;
wire un36_prod_a_b_cry_5_RNO ;
wire un36_prod_a_b_cry_6_RNO ;
wire un36_prod_a_b_cry_7_RNO ;
wire un36_prod_a_b_cry_8_RNO ;
wire un36_prod_a_b_cry_9_RNO ;
wire un36_prod_a_b_cry_10_RNO ;
wire un36_prod_a_b_cry_11_RNO ;
wire un36_prod_a_b_cry_12_RNO ;
wire un36_prod_a_b_cry_13_RNO ;
wire un36_prod_a_b_cry_14_RNO ;
wire un36_prod_a_b_cry_15_RNO ;
wire un36_prod_a_b_cry_16_RNO ;
wire un36_prod_a_b_cry_17_RNO ;
wire un36_prod_a_b_cry_18_RNO ;
wire un36_prod_a_b_cry_19_RNO ;
wire un36_prod_a_b_cry_20_RNO ;
wire un36_prod_a_b_cry_21_RNO ;
wire un36_prod_a_b_cry_22_RNO ;
wire un54_sum_cry_0_RNO ;
wire un54_sum_cry_1_RNO ;
wire un54_sum_cry_2_RNO ;
wire un54_sum_cry_3_RNO ;
wire un54_sum_cry_4_RNO ;
wire un54_sum_cry_5_RNO ;
wire un54_sum_cry_6_RNO ;
wire un54_sum_cry_7_RNO ;
wire un54_sum_cry_8_RNO ;
wire un54_sum_cry_9_RNO ;
wire un54_sum_cry_10_RNO ;
wire un54_sum_cry_11_RNO ;
wire un54_sum_cry_15 ;
wire un54_sum_cry_14 ;
wire un54_sum_cry_13 ;
wire un54_sum_cry_12 ;
wire un54_sum_cry_11 ;
wire un54_sum_cry_10 ;
wire un54_sum_cry_9 ;
wire un54_sum_cry_8 ;
wire un54_sum_cry_7 ;
wire un54_sum_cry_6 ;
wire un54_sum_cry_5 ;
wire un54_sum_cry_4 ;
wire un54_sum_cry_3 ;
wire un54_sum_cry_2 ;
wire un54_sum_cry_1 ;
wire un54_sum_cry_0 ;
wire un36_prod_a_b_cry_33 ;
wire un36_prod_a_b_cry_32 ;
wire un36_prod_a_b_cry_31 ;
wire un36_prod_a_b_cry_30 ;
wire un36_prod_a_b_cry_29 ;
wire un36_prod_a_b_cry_28 ;
wire un36_prod_a_b_cry_27 ;
wire un36_prod_a_b_cry_26 ;
wire un36_prod_a_b_cry_25 ;
wire un36_prod_a_b_cry_24 ;
wire un36_prod_a_b_cry_23 ;
wire un36_prod_a_b_cry_22 ;
wire un36_prod_a_b_cry_21 ;
wire un36_prod_a_b_cry_20 ;
wire un36_prod_a_b_cry_19 ;
wire un36_prod_a_b_cry_18 ;
wire un36_prod_a_b_cry_17 ;
wire un36_prod_a_b_cry_16 ;
wire un36_prod_a_b_cry_15 ;
wire un36_prod_a_b_cry_14 ;
wire un36_prod_a_b_cry_13 ;
wire un36_prod_a_b_cry_12 ;
wire un36_prod_a_b_cry_11 ;
wire un36_prod_a_b_cry_10 ;
wire un36_prod_a_b_cry_9 ;
wire un36_prod_a_b_cry_8 ;
wire un36_prod_a_b_cry_7 ;
wire un36_prod_a_b_cry_6 ;
wire un36_prod_a_b_cry_5 ;
wire un36_prod_a_b_cry_4 ;
wire un36_prod_a_b_cry_3 ;
wire un36_prod_a_b_cry_2 ;
wire un36_prod_a_b_cry_1 ;
wire un36_prod_a_b_cry_0 ;
wire CARRYCASCOUT ;
wire MULTSIGNOUT ;
wire OVERFLOW ;
wire PATTERNBDETECT ;
wire PATTERNDETECT ;
wire UNDERFLOW ;
wire CARRYCASCOUT_0 ;
wire MULTSIGNOUT_0 ;
wire OVERFLOW_0 ;
wire PATTERNBDETECT_0 ;
wire PATTERNDETECT_0 ;
wire UNDERFLOW_0 ;
wire CARRYCASCOUT_1 ;
wire MULTSIGNOUT_1 ;
wire OVERFLOW_1 ;
wire PATTERNBDETECT_1 ;
wire PATTERNDETECT_1 ;
wire UNDERFLOW_1 ;
wire CARRYCASCOUT_2 ;
wire MULTSIGNOUT_2 ;
wire OVERFLOW_2 ;
wire PATTERNBDETECT_2 ;
wire PATTERNDETECT_2 ;
wire UNDERFLOW_2 ;
wire N_1 ;
// instances
  FDR desc605(.Q(count[2:2]),.D(m39),.C(clk_i),.R(s_start_i));
  FD desc606(.Q(s_fractb_i[23:23]),.D(result_1_i_o3_0_e),.C(clk_i));
  FDS desc607(.Q(s_state),.D(N_2731_i_0_0),.C(clk_i),.S(s_start_i));
  LUT4 desc608(.I0(N_85_0),.I1(N_142_0),.I2(N_145_0_i),.I3(N_3283),.O(un54_sum_axb_11));
defparam desc608.INIT=16'hE187;
  FD s_signa_i_Z(.Q(s_signa_i),.D(s_opa_i_31),.C(clk_i));
  FD s_signb_i_Z(.Q(s_signb_i),.D(s_opb_i_31),.C(clk_i));
  FDE desc609(.Q(sum_0[23:23]),.D(un54_sum[670:670]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc610(.Q(sum_1[23:23]),.D(un54_sum[670:670]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc611(.Q(sum_2[23:23]),.D(un54_sum[670:670]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc612(.Q(sum_3[23:23]),.D(un54_sum[670:670]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc613(.Q(sum_0[22:22]),.D(un54_sum[669:669]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc614(.Q(sum_1[22:22]),.D(un54_sum[669:669]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc615(.Q(sum_2[22:22]),.D(un54_sum[669:669]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc616(.Q(sum_3[22:22]),.D(un54_sum[669:669]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc617(.Q(sum_0[21:21]),.D(un54_sum[668:668]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc618(.Q(sum_1[21:21]),.D(un54_sum[668:668]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc619(.Q(sum_2[21:21]),.D(un54_sum[668:668]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc620(.Q(sum_3[21:21]),.D(un54_sum[668:668]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc621(.Q(sum_0[20:20]),.D(un54_sum[667:667]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc622(.Q(sum_1[20:20]),.D(un54_sum[667:667]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc623(.Q(sum_2[20:20]),.D(un54_sum[667:667]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc624(.Q(sum_3[20:20]),.D(un54_sum[667:667]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc625(.Q(sum_0[19:19]),.D(un54_sum[666:666]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc626(.Q(sum_1[19:19]),.D(un54_sum[666:666]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc627(.Q(sum_2[19:19]),.D(un54_sum[666:666]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc628(.Q(sum_3[19:19]),.D(un54_sum[666:666]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc629(.Q(sum_0[18:18]),.D(un54_sum[665:665]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc630(.Q(sum_1[18:18]),.D(un54_sum[665:665]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc631(.Q(sum_2[18:18]),.D(un54_sum[665:665]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc632(.Q(sum_3[18:18]),.D(un54_sum[665:665]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc633(.Q(sum_0[17:17]),.D(un54_sum[664:664]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc634(.Q(sum_1[17:17]),.D(un54_sum[664:664]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc635(.Q(sum_2[17:17]),.D(un54_sum[664:664]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc636(.Q(sum_3[17:17]),.D(un54_sum[664:664]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc637(.Q(sum_0[16:16]),.D(un54_sum[663:663]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc638(.Q(sum_1[16:16]),.D(un54_sum[663:663]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc639(.Q(sum_2[16:16]),.D(un54_sum[663:663]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc640(.Q(sum_3[16:16]),.D(un54_sum[663:663]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc641(.Q(sum_0[15:15]),.D(un54_sum[662:662]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc642(.Q(sum_1[15:15]),.D(un54_sum[662:662]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc643(.Q(sum_2[15:15]),.D(un54_sum[662:662]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc644(.Q(sum_3[15:15]),.D(un54_sum[662:662]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc645(.Q(sum_0[14:14]),.D(un54_sum[661:661]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc646(.Q(sum_1[14:14]),.D(un54_sum[661:661]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc647(.Q(sum_2[14:14]),.D(un54_sum[661:661]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc648(.Q(sum_3[14:14]),.D(un54_sum[661:661]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc649(.Q(sum_0[13:13]),.D(un54_sum[660:660]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc650(.Q(sum_1[13:13]),.D(un54_sum[660:660]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc651(.Q(sum_2[13:13]),.D(un54_sum[660:660]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc652(.Q(sum_3[13:13]),.D(un54_sum[660:660]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc653(.Q(sum_0[12:12]),.D(un54_sum[659:659]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc654(.Q(sum_1[12:12]),.D(un54_sum[659:659]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc655(.Q(sum_2[12:12]),.D(un54_sum[659:659]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc656(.Q(sum_3[12:12]),.D(un54_sum[659:659]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc657(.Q(sum_0[11:11]),.D(un54_sum[658:658]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc658(.Q(sum_1[11:11]),.D(un54_sum[658:658]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc659(.Q(sum_2[11:11]),.D(un54_sum[658:658]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc660(.Q(mul_24_fract_48[11:11]),.D(un54_sum[658:658]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc661(.Q(sum_0[10:10]),.D(un54_sum[657:657]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc662(.Q(sum_1[10:10]),.D(un54_sum[657:657]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc663(.Q(sum_2[10:10]),.D(un54_sum[657:657]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc664(.Q(mul_24_fract_48[10:10]),.D(un54_sum[657:657]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc665(.Q(sum_0[9:9]),.D(un54_sum[656:656]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc666(.Q(sum_1[9:9]),.D(un54_sum[656:656]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc667(.Q(sum_2[9:9]),.D(un54_sum[656:656]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc668(.Q(mul_24_fract_48[9:9]),.D(un54_sum[656:656]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc669(.Q(sum_0[8:8]),.D(un54_sum[655:655]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc670(.Q(sum_1[8:8]),.D(un54_sum[655:655]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc671(.Q(sum_2[8:8]),.D(un54_sum[655:655]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc672(.Q(mul_24_fract_48[8:8]),.D(un54_sum[655:655]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc673(.Q(sum_0[7:7]),.D(un54_sum[654:654]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc674(.Q(sum_1[7:7]),.D(un54_sum[654:654]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc675(.Q(sum_2[7:7]),.D(un54_sum[654:654]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc676(.Q(mul_24_fract_48[7:7]),.D(un54_sum[654:654]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc677(.Q(sum_0[6:6]),.D(un54_sum[653:653]),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc678(.Q(sum_1[6:6]),.D(un54_sum[653:653]),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc679(.Q(sum_2[6:6]),.D(un54_sum[653:653]),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc680(.Q(mul_24_fract_48[6:6]),.D(un54_sum[653:653]),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc681(.Q(sum_0[5:5]),.D(N_103_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc682(.Q(sum_1[5:5]),.D(N_103_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc683(.Q(sum_2[5:5]),.D(N_103_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc684(.Q(mul_24_fract_48[5:5]),.D(N_103_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc685(.Q(sum_0[4:4]),.D(N_100_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc686(.Q(sum_1[4:4]),.D(N_100_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc687(.Q(sum_2[4:4]),.D(N_100_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc688(.Q(mul_24_fract_48[4:4]),.D(N_100_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc689(.Q(sum_0[3:3]),.D(N_97_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc690(.Q(sum_1[3:3]),.D(N_97_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc691(.Q(sum_2[3:3]),.D(N_97_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc692(.Q(mul_24_fract_48[3:3]),.D(N_97_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc693(.Q(sum_0[2:2]),.D(N_94_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc694(.Q(sum_1[2:2]),.D(N_94_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc695(.Q(sum_2[2:2]),.D(N_94_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc696(.Q(mul_24_fract_48[2:2]),.D(N_94_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc697(.Q(sum_0[1:1]),.D(N_91_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc698(.Q(sum_1[1:1]),.D(N_91_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc699(.Q(sum_2[1:1]),.D(N_91_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc700(.Q(mul_24_fract_48[1:1]),.D(N_91_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FDE desc701(.Q(sum_0[0:0]),.D(N_88_0_i),.C(clk_i),.CE(count_RNILIBD_2_O5[2:2]));
  FDE desc702(.Q(sum_1[0:0]),.D(N_88_0_i),.C(clk_i),.CE(count_RNILIBD_0_O5[2:2]));
  FDE desc703(.Q(sum_2[0:0]),.D(N_88_0_i),.C(clk_i),.CE(count_RNILIBD_O5[2:2]));
  FDE desc704(.Q(mul_24_fract_48[0:0]),.D(N_88_0_i),.C(clk_i),.CE(count_RNILIBD_1_O6[2:2]));
  FD desc705(.Q(s_fractb_i_11),.D(s_opb_i_11),.C(clk_i));
  FDE desc706(.Q(prod2_2_0[23:23]),.D(un23_prod2[11:11]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc707(.Q(prod2_0_0[23:23]),.D(un23_prod2[11:11]),.C(clk_i),.CE(un2_i));
  FDE desc708(.Q(prod2_1_0[23:23]),.D(un23_prod2[11:11]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc709(.Q(prod2_3_0[23:23]),.D(un23_prod2[11:11]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc710(.Q(prod2_2_0[22:22]),.D(un23_prod2[10:10]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc711(.Q(prod2_0_0[22:22]),.D(un23_prod2[10:10]),.C(clk_i),.CE(un2_i));
  FDE desc712(.Q(prod2_1_0[22:22]),.D(un23_prod2[10:10]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc713(.Q(prod2_3_0[22:22]),.D(un23_prod2[10:10]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc714(.Q(prod2_2_0[21:21]),.D(un23_prod2[9:9]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc715(.Q(prod2_0_0[21:21]),.D(un23_prod2[9:9]),.C(clk_i),.CE(un2_i));
  FDE desc716(.Q(prod2_1_0[21:21]),.D(un23_prod2[9:9]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc717(.Q(prod2_3_0[21:21]),.D(un23_prod2[9:9]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc718(.Q(prod2_2_0[20:20]),.D(un23_prod2[8:8]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc719(.Q(prod2_0_0[20:20]),.D(un23_prod2[8:8]),.C(clk_i),.CE(un2_i));
  FDE desc720(.Q(prod2_1_0[20:20]),.D(un23_prod2[8:8]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc721(.Q(prod2_3_0[20:20]),.D(un23_prod2[8:8]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc722(.Q(prod2_2_0[19:19]),.D(un23_prod2[7:7]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc723(.Q(prod2_0_0[19:19]),.D(un23_prod2[7:7]),.C(clk_i),.CE(un2_i));
  FDE desc724(.Q(prod2_1_0[19:19]),.D(un23_prod2[7:7]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc725(.Q(prod2_3_0[19:19]),.D(un23_prod2[7:7]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc726(.Q(prod2_2_0[18:18]),.D(un23_prod2[6:6]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc727(.Q(prod2_0_0[18:18]),.D(un23_prod2[6:6]),.C(clk_i),.CE(un2_i));
  FDE desc728(.Q(prod2_1_0[18:18]),.D(un23_prod2[6:6]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc729(.Q(prod2_3_0[18:18]),.D(un23_prod2[6:6]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc730(.Q(prod2_2_0[17:17]),.D(un23_prod2[5:5]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc731(.Q(prod2_0_0[17:17]),.D(un23_prod2[5:5]),.C(clk_i),.CE(un2_i));
  FDE desc732(.Q(prod2_1_0[17:17]),.D(un23_prod2[5:5]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc733(.Q(prod2_3_0[17:17]),.D(un23_prod2[5:5]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc734(.Q(prod2_2_0[16:16]),.D(un23_prod2[4:4]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc735(.Q(prod2_0_0[16:16]),.D(un23_prod2[4:4]),.C(clk_i),.CE(un2_i));
  FDE desc736(.Q(prod2_1_0[16:16]),.D(un23_prod2[4:4]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc737(.Q(prod2_3_0[16:16]),.D(un23_prod2[4:4]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc738(.Q(prod2_2_0[15:15]),.D(un23_prod2[3:3]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc739(.Q(prod2_0_0[15:15]),.D(un23_prod2[3:3]),.C(clk_i),.CE(un2_i));
  FDE desc740(.Q(prod2_1_0[15:15]),.D(un23_prod2[3:3]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc741(.Q(prod2_3_0[15:15]),.D(un23_prod2[3:3]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc742(.Q(prod2_2_0[14:14]),.D(un23_prod2[2:2]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc743(.Q(prod2_0_0[14:14]),.D(un23_prod2[2:2]),.C(clk_i),.CE(un2_i));
  FDE desc744(.Q(prod2_1_0[14:14]),.D(un23_prod2[2:2]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc745(.Q(prod2_3_0[14:14]),.D(un23_prod2[2:2]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc746(.Q(prod2_2_0[13:13]),.D(un23_prod2[1:1]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc747(.Q(prod2_0_0[13:13]),.D(un23_prod2[1:1]),.C(clk_i),.CE(un2_i));
  FDE desc748(.Q(prod2_1_0[13:13]),.D(un23_prod2[1:1]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc749(.Q(prod2_3_0[13:13]),.D(un23_prod2[1:1]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc750(.Q(prod2_2_0[12:12]),.D(un23_prod2[0:0]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc751(.Q(prod2_0_0[12:12]),.D(un23_prod2[0:0]),.C(clk_i),.CE(un2_i));
  FDE desc752(.Q(prod2_1_0[12:12]),.D(un23_prod2[0:0]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc753(.Q(prod2_3_0[12:12]),.D(un23_prod2[0:0]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FD desc754(.Q(s_fracta_i[11:11]),.D(s_opa_i_11),.C(clk_i));
  FD desc755(.Q(s_fracta_i[10:10]),.D(s_opa_i_10),.C(clk_i));
  FD desc756(.Q(s_fracta_i[22:22]),.D(s_opa_i_22),.C(clk_i));
  FD desc757(.Q(s_fracta_i[9:9]),.D(s_opa_i_9),.C(clk_i));
  FD desc758(.Q(s_fracta_i[21:21]),.D(s_opa_i_21),.C(clk_i));
  FD desc759(.Q(s_fracta_i[8:8]),.D(s_opa_i_8),.C(clk_i));
  FD desc760(.Q(s_fracta_i[20:20]),.D(s_opa_i_20),.C(clk_i));
  FD desc761(.Q(s_fracta_i[7:7]),.D(s_opa_i_7),.C(clk_i));
  FD desc762(.Q(s_fracta_i[19:19]),.D(s_opa_i_19),.C(clk_i));
  FD desc763(.Q(s_fracta_i[6:6]),.D(s_opa_i_6),.C(clk_i));
  FD desc764(.Q(s_fracta_i[18:18]),.D(s_opa_i_18),.C(clk_i));
  FD desc765(.Q(s_fractb_i_10),.D(s_opb_i_10),.C(clk_i));
  FD desc766(.Q(s_fractb_i_22),.D(s_opb_i_22),.C(clk_i));
  FD desc767(.Q(s_fractb_i_9),.D(s_opb_i_9),.C(clk_i));
  FD desc768(.Q(s_fractb_i_21),.D(s_opb_i_21),.C(clk_i));
  FD desc769(.Q(s_fractb_i_8),.D(s_opb_i_8),.C(clk_i));
  FD desc770(.Q(s_fractb_i_20),.D(s_opb_i_20),.C(clk_i));
  FD desc771(.Q(s_fractb_i_7),.D(s_opb_i_7),.C(clk_i));
  FD desc772(.Q(s_fractb_i_19),.D(s_opb_i_19),.C(clk_i));
  FD desc773(.Q(s_fractb_i_6),.D(s_opb_i_6),.C(clk_i));
  FD desc774(.Q(s_fractb_i_18),.D(s_opb_i_18),.C(clk_i));
  FDE desc775(.Q(prod2_0_1[17:17]),.D(un92_prod2[11:11]),.C(clk_i),.CE(un2_i));
  FDE desc776(.Q(prod2_1_1[17:17]),.D(un92_prod2[11:11]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc777(.Q(prod2_2_1[17:17]),.D(un92_prod2[11:11]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc778(.Q(prod2_3_1[17:17]),.D(un92_prod2[11:11]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc779(.Q(prod2_0_1[16:16]),.D(un92_prod2[10:10]),.C(clk_i),.CE(un2_i));
  FDE desc780(.Q(prod2_1_1[16:16]),.D(un92_prod2[10:10]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc781(.Q(prod2_2_1[16:16]),.D(un92_prod2[10:10]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc782(.Q(prod2_3_1[16:16]),.D(un92_prod2[10:10]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc783(.Q(prod2_0_1[15:15]),.D(un92_prod2[9:9]),.C(clk_i),.CE(un2_i));
  FDE desc784(.Q(prod2_1_1[15:15]),.D(un92_prod2[9:9]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc785(.Q(prod2_2_1[15:15]),.D(un92_prod2[9:9]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc786(.Q(prod2_3_1[15:15]),.D(un92_prod2[9:9]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc787(.Q(prod2_0_1[14:14]),.D(un92_prod2[8:8]),.C(clk_i),.CE(un2_i));
  FDE desc788(.Q(prod2_1_1[14:14]),.D(un92_prod2[8:8]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc789(.Q(prod2_2_1[14:14]),.D(un92_prod2[8:8]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc790(.Q(prod2_3_1[14:14]),.D(un92_prod2[8:8]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc791(.Q(prod2_0_1[13:13]),.D(un92_prod2[7:7]),.C(clk_i),.CE(un2_i));
  FDE desc792(.Q(prod2_1_1[13:13]),.D(un92_prod2[7:7]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc793(.Q(prod2_2_1[13:13]),.D(un92_prod2[7:7]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc794(.Q(prod2_3_1[13:13]),.D(un92_prod2[7:7]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc795(.Q(prod2_0_1[12:12]),.D(un92_prod2[6:6]),.C(clk_i),.CE(un2_i));
  FDE desc796(.Q(prod2_1_1[12:12]),.D(un92_prod2[6:6]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc797(.Q(prod2_2_1[12:12]),.D(un92_prod2[6:6]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc798(.Q(prod2_3_1[12:12]),.D(un92_prod2[6:6]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc799(.Q(prod2_0_1[11:11]),.D(un92_prod2[5:5]),.C(clk_i),.CE(un2_i));
  FDE desc800(.Q(prod2_1_1[11:11]),.D(un92_prod2[5:5]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc801(.Q(prod2_2_1[11:11]),.D(un92_prod2[5:5]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc802(.Q(prod2_3_1[11:11]),.D(un92_prod2[5:5]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc803(.Q(prod2_0_1[10:10]),.D(un92_prod2[4:4]),.C(clk_i),.CE(un2_i));
  FDE desc804(.Q(prod2_1_1[10:10]),.D(un92_prod2[4:4]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc805(.Q(prod2_2_1[10:10]),.D(un92_prod2[4:4]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc806(.Q(prod2_3_1[10:10]),.D(un92_prod2[4:4]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc807(.Q(prod2_0_1[9:9]),.D(un92_prod2[3:3]),.C(clk_i),.CE(un2_i));
  FDE desc808(.Q(prod2_1_1[9:9]),.D(un92_prod2[3:3]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc809(.Q(prod2_2_1[9:9]),.D(un92_prod2[3:3]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc810(.Q(prod2_3_1[9:9]),.D(un92_prod2[3:3]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc811(.Q(prod2_0_1[8:8]),.D(un92_prod2[2:2]),.C(clk_i),.CE(un2_i));
  FDE desc812(.Q(prod2_1_1[8:8]),.D(un92_prod2[2:2]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc813(.Q(prod2_2_1[8:8]),.D(un92_prod2[2:2]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc814(.Q(prod2_3_1[8:8]),.D(un92_prod2[2:2]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc815(.Q(prod2_0_1[7:7]),.D(un92_prod2[1:1]),.C(clk_i),.CE(un2_i));
  FDE desc816(.Q(prod2_1_1[7:7]),.D(un92_prod2[1:1]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc817(.Q(prod2_2_1[7:7]),.D(un92_prod2[1:1]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc818(.Q(prod2_3_1[7:7]),.D(un92_prod2[1:1]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc819(.Q(prod2_0_1[6:6]),.D(un92_prod2[0:0]),.C(clk_i),.CE(un2_i));
  FDE desc820(.Q(prod2_1_1[6:6]),.D(un92_prod2[0:0]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc821(.Q(prod2_2_1[6:6]),.D(un92_prod2[0:0]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc822(.Q(prod2_3_1[6:6]),.D(un92_prod2[0:0]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc823(.Q(prod2_0_2[17:17]),.D(un139_prod2[11:11]),.C(clk_i),.CE(un2_i));
  FDE desc824(.Q(prod2_1_2[17:17]),.D(un139_prod2[11:11]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc825(.Q(prod2_2_2[17:17]),.D(un139_prod2[11:11]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc826(.Q(prod2_3_2[17:17]),.D(un139_prod2[11:11]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc827(.Q(prod2_0_2[16:16]),.D(un139_prod2[10:10]),.C(clk_i),.CE(un2_i));
  FDE desc828(.Q(prod2_1_2[16:16]),.D(un139_prod2[10:10]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc829(.Q(prod2_2_2[16:16]),.D(un139_prod2[10:10]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc830(.Q(prod2_3_2[16:16]),.D(un139_prod2[10:10]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc831(.Q(prod2_0_2[15:15]),.D(un139_prod2[9:9]),.C(clk_i),.CE(un2_i));
  FDE desc832(.Q(prod2_1_2[15:15]),.D(un139_prod2[9:9]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc833(.Q(prod2_2_2[15:15]),.D(un139_prod2[9:9]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc834(.Q(prod2_3_2[15:15]),.D(un139_prod2[9:9]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc835(.Q(prod2_0_2[14:14]),.D(un139_prod2[8:8]),.C(clk_i),.CE(un2_i));
  FDE desc836(.Q(prod2_1_2[14:14]),.D(un139_prod2[8:8]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc837(.Q(prod2_2_2[14:14]),.D(un139_prod2[8:8]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc838(.Q(prod2_3_2[14:14]),.D(un139_prod2[8:8]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc839(.Q(prod2_0_2[13:13]),.D(un139_prod2[7:7]),.C(clk_i),.CE(un2_i));
  FDE desc840(.Q(prod2_1_2[13:13]),.D(un139_prod2[7:7]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc841(.Q(prod2_2_2[13:13]),.D(un139_prod2[7:7]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc842(.Q(prod2_3_2[13:13]),.D(un139_prod2[7:7]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc843(.Q(prod2_0_2[12:12]),.D(un139_prod2[6:6]),.C(clk_i),.CE(un2_i));
  FDE desc844(.Q(prod2_1_2[12:12]),.D(un139_prod2[6:6]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc845(.Q(prod2_2_2[12:12]),.D(un139_prod2[6:6]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc846(.Q(prod2_3_2[12:12]),.D(un139_prod2[6:6]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc847(.Q(prod2_0_2[11:11]),.D(un139_prod2[5:5]),.C(clk_i),.CE(un2_i));
  FDE desc848(.Q(prod2_1_2[11:11]),.D(un139_prod2[5:5]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc849(.Q(prod2_2_2[11:11]),.D(un139_prod2[5:5]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc850(.Q(prod2_3_2[11:11]),.D(un139_prod2[5:5]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc851(.Q(prod2_0_2[10:10]),.D(un139_prod2[4:4]),.C(clk_i),.CE(un2_i));
  FDE desc852(.Q(prod2_1_2[10:10]),.D(un139_prod2[4:4]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc853(.Q(prod2_2_2[10:10]),.D(un139_prod2[4:4]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc854(.Q(prod2_3_2[10:10]),.D(un139_prod2[4:4]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc855(.Q(prod2_0_2[9:9]),.D(un139_prod2[3:3]),.C(clk_i),.CE(un2_i));
  FDE desc856(.Q(prod2_1_2[9:9]),.D(un139_prod2[3:3]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc857(.Q(prod2_2_2[9:9]),.D(un139_prod2[3:3]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc858(.Q(prod2_3_2[9:9]),.D(un139_prod2[3:3]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc859(.Q(prod2_0_2[8:8]),.D(un139_prod2[2:2]),.C(clk_i),.CE(un2_i));
  FDE desc860(.Q(prod2_1_2[8:8]),.D(un139_prod2[2:2]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc861(.Q(prod2_2_2[8:8]),.D(un139_prod2[2:2]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc862(.Q(prod2_3_2[8:8]),.D(un139_prod2[2:2]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc863(.Q(prod2_0_2[7:7]),.D(un139_prod2[1:1]),.C(clk_i),.CE(un2_i));
  FDE desc864(.Q(prod2_1_2[7:7]),.D(un139_prod2[1:1]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc865(.Q(prod2_2_2[7:7]),.D(un139_prod2[1:1]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc866(.Q(prod2_3_2[7:7]),.D(un139_prod2[1:1]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc867(.Q(prod2_0_2[6:6]),.D(un139_prod2[0:0]),.C(clk_i),.CE(un2_i));
  FDE desc868(.Q(prod2_1_2[6:6]),.D(un139_prod2[0:0]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc869(.Q(prod2_2_2[6:6]),.D(un139_prod2[0:0]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc870(.Q(prod2_3_2[6:6]),.D(un139_prod2[0:0]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FD desc871(.Q(s_fractb_i_5),.D(s_opb_i_5),.C(clk_i));
  FD desc872(.Q(s_fractb_i_17),.D(s_opb_i_17),.C(clk_i));
  FD desc873(.Q(s_fractb_i_4),.D(s_opb_i_4),.C(clk_i));
  FD desc874(.Q(s_fractb_i_16),.D(s_opb_i_16),.C(clk_i));
  FD desc875(.Q(s_fractb_i_3),.D(s_opb_i_3),.C(clk_i));
  FD desc876(.Q(s_fractb_i_15),.D(s_opb_i_15),.C(clk_i));
  FD desc877(.Q(s_fractb_i_2),.D(s_opb_i_2),.C(clk_i));
  FD desc878(.Q(s_fractb_i_14),.D(s_opb_i_14),.C(clk_i));
  FD desc879(.Q(s_fractb_i_1),.D(s_opb_i_1),.C(clk_i));
  FD desc880(.Q(s_fractb_i_13),.D(s_opb_i_13),.C(clk_i));
  FD desc881(.Q(s_fractb_i_0),.D(s_opb_i_0),.C(clk_i));
  FD desc882(.Q(s_fractb_i_12),.D(s_opb_i_12),.C(clk_i));
  FD desc883(.Q(s_fracta_i[5:5]),.D(s_opa_i_5),.C(clk_i));
  FD desc884(.Q(s_fracta_i[17:17]),.D(s_opa_i_17),.C(clk_i));
  FD desc885(.Q(s_fracta_i[4:4]),.D(s_opa_i_4),.C(clk_i));
  FD desc886(.Q(s_fracta_i[16:16]),.D(s_opa_i_16),.C(clk_i));
  FD desc887(.Q(s_fracta_i[3:3]),.D(s_opa_i_3),.C(clk_i));
  FD desc888(.Q(s_fracta_i[15:15]),.D(s_opa_i_15),.C(clk_i));
  FD desc889(.Q(s_fracta_i[2:2]),.D(s_opa_i_2),.C(clk_i));
  FD desc890(.Q(s_fracta_i[14:14]),.D(s_opa_i_14),.C(clk_i));
  FD desc891(.Q(s_fracta_i[1:1]),.D(s_opa_i_1),.C(clk_i));
  FD desc892(.Q(s_fracta_i[13:13]),.D(s_opa_i_13),.C(clk_i));
  FD desc893(.Q(s_fracta_i[0:0]),.D(s_opa_i_0),.C(clk_i));
  FD desc894(.Q(s_fracta_i[12:12]),.D(s_opa_i_12),.C(clk_i));
  FDE desc895(.Q(prod2_0_3[11:11]),.D(un184_prod2[11:11]),.C(clk_i),.CE(un2_i));
  FDE desc896(.Q(prod2_1_3[11:11]),.D(un184_prod2[11:11]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc897(.Q(prod2_2_3[11:11]),.D(un184_prod2[11:11]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc898(.Q(prod2_3_3[11:11]),.D(un184_prod2[11:11]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc899(.Q(prod2_0_3[10:10]),.D(un184_prod2[10:10]),.C(clk_i),.CE(un2_i));
  FDE desc900(.Q(prod2_1_3[10:10]),.D(un184_prod2[10:10]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc901(.Q(prod2_2_3[10:10]),.D(un184_prod2[10:10]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc902(.Q(prod2_3_3[10:10]),.D(un184_prod2[10:10]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc903(.Q(prod2_0_3[9:9]),.D(un184_prod2[9:9]),.C(clk_i),.CE(un2_i));
  FDE desc904(.Q(prod2_1_3[9:9]),.D(un184_prod2[9:9]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc905(.Q(prod2_2_3[9:9]),.D(un184_prod2[9:9]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc906(.Q(prod2_3_3[9:9]),.D(un184_prod2[9:9]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc907(.Q(prod2_0_3[8:8]),.D(un184_prod2[8:8]),.C(clk_i),.CE(un2_i));
  FDE desc908(.Q(prod2_1_3[8:8]),.D(un184_prod2[8:8]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc909(.Q(prod2_2_3[8:8]),.D(un184_prod2[8:8]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc910(.Q(prod2_3_3[8:8]),.D(un184_prod2[8:8]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc911(.Q(prod2_0_3[7:7]),.D(un184_prod2[7:7]),.C(clk_i),.CE(un2_i));
  FDE desc912(.Q(prod2_1_3[7:7]),.D(un184_prod2[7:7]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc913(.Q(prod2_2_3[7:7]),.D(un184_prod2[7:7]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc914(.Q(prod2_3_3[7:7]),.D(un184_prod2[7:7]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc915(.Q(prod2_0_3[6:6]),.D(un184_prod2[6:6]),.C(clk_i),.CE(un2_i));
  FDE desc916(.Q(prod2_1_3[6:6]),.D(un184_prod2[6:6]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc917(.Q(prod2_2_3[6:6]),.D(un184_prod2[6:6]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc918(.Q(prod2_3_3[6:6]),.D(un184_prod2[6:6]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc919(.Q(prod2_0_3[5:5]),.D(un184_prod2[5:5]),.C(clk_i),.CE(un2_i));
  FDE desc920(.Q(prod2_1_3[5:5]),.D(un184_prod2[5:5]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc921(.Q(prod2_2_3[5:5]),.D(un184_prod2[5:5]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc922(.Q(prod2_3_3[5:5]),.D(un184_prod2[5:5]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc923(.Q(prod2_0_3[4:4]),.D(un184_prod2[4:4]),.C(clk_i),.CE(un2_i));
  FDE desc924(.Q(prod2_1_3[4:4]),.D(un184_prod2[4:4]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc925(.Q(prod2_2_3[4:4]),.D(un184_prod2[4:4]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc926(.Q(prod2_3_3[4:4]),.D(un184_prod2[4:4]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc927(.Q(prod2_0_3[3:3]),.D(un184_prod2[3:3]),.C(clk_i),.CE(un2_i));
  FDE desc928(.Q(prod2_1_3[3:3]),.D(un184_prod2[3:3]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc929(.Q(prod2_2_3[3:3]),.D(un184_prod2[3:3]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc930(.Q(prod2_3_3[3:3]),.D(un184_prod2[3:3]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc931(.Q(prod2_0_3[2:2]),.D(un184_prod2[2:2]),.C(clk_i),.CE(un2_i));
  FDE desc932(.Q(prod2_1_3[2:2]),.D(un184_prod2[2:2]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc933(.Q(prod2_2_3[2:2]),.D(un184_prod2[2:2]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc934(.Q(prod2_3_3[2:2]),.D(un184_prod2[2:2]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc935(.Q(prod2_0_3[1:1]),.D(un184_prod2[1:1]),.C(clk_i),.CE(un2_i));
  FDE desc936(.Q(prod2_1_3[1:1]),.D(un184_prod2[1:1]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc937(.Q(prod2_2_3[1:1]),.D(un184_prod2[1:1]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc938(.Q(prod2_3_3[1:1]),.D(un184_prod2[1:1]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  FDE desc939(.Q(prod2_0_3[0:0]),.D(un184_prod2[0:0]),.C(clk_i),.CE(un2_i));
  FDE desc940(.Q(prod2_1_3[0:0]),.D(un184_prod2[0:0]),.C(clk_i),.CE(prod2_1_0_1_sqmuxa));
  FDE desc941(.Q(prod2_2_3[0:0]),.D(un184_prod2[0:0]),.C(clk_i),.CE(prod2_2_0_1_sqmuxa));
  FDE desc942(.Q(prod2_3_3[0:0]),.D(un184_prod2[0:0]),.C(clk_i),.CE(prod2_3_0_1_sqmuxa));
  LUT6_L desc943(.I0(sum_0[7:7]),.I1(sum_0[8:8]),.I2(sum_1[19:19]),.I3(sum_1[20:20]),.I4(sum_2[19:19]),.I5(sum_2[20:20]),.LO(un36_prod_a_b_axb_19));
defparam desc943.INIT=64'h36C96C93C936936C;
  LUT6_L desc944(.I0(sum_0[6:6]),.I1(sum_0[7:7]),.I2(sum_1[18:18]),.I3(sum_1[19:19]),.I4(sum_2[18:18]),.I5(sum_2[19:19]),.LO(un36_prod_a_b_axb_18));
defparam desc944.INIT=64'h36C96C93C936936C;
  LUT6_L desc945(.I0(sum_0[4:4]),.I1(sum_0[5:5]),.I2(sum_1[16:16]),.I3(sum_1[17:17]),.I4(sum_2[16:16]),.I5(sum_2[17:17]),.LO(un36_prod_a_b_axb_16));
defparam desc945.INIT=64'h36C96C93C936936C;
  LUT6_L desc946(.I0(sum_0[1:1]),.I1(sum_0[2:2]),.I2(sum_1[13:13]),.I3(sum_1[14:14]),.I4(sum_2[13:13]),.I5(sum_2[14:14]),.LO(un36_prod_a_b_axb_13));
defparam desc946.INIT=64'h36C96C93C936936C;
  LUT6_L desc947(.I0(sum_0[0:0]),.I1(sum_0[1:1]),.I2(sum_1[12:12]),.I3(sum_1[13:13]),.I4(sum_2[12:12]),.I5(sum_2[13:13]),.LO(un36_prod_a_b_axb_12));
defparam desc947.INIT=64'h36C96C93C936936C;
  LUT6_L desc948(.I0(sum_1[10:10]),.I1(sum_1[11:11]),.I2(sum_2[10:10]),.I3(sum_2[11:11]),.I4(sum_3[22:22]),.I5(sum_3[23:23]),.LO(un36_prod_a_b_axb_10));
defparam desc948.INIT=64'h36C96C93C936936C;
  LUT6_L desc949(.I0(sum_1[6:6]),.I1(sum_1[7:7]),.I2(sum_2[6:6]),.I3(sum_2[7:7]),.I4(sum_3[18:18]),.I5(sum_3[19:19]),.LO(un36_prod_a_b_axb_6));
defparam desc949.INIT=64'h36C96C93C936936C;
  LUT6_L desc950(.I0(sum_1[4:4]),.I1(sum_1[5:5]),.I2(sum_2[4:4]),.I3(sum_2[5:5]),.I4(sum_3[16:16]),.I5(sum_3[17:17]),.LO(un36_prod_a_b_axb_4));
defparam desc950.INIT=64'h36C96C93C936936C;
  LUT6_L desc951(.I0(sum_0[10:10]),.I1(sum_0[11:11]),.I2(sum_1[22:22]),.I3(sum_1[23:23]),.I4(sum_2[22:22]),.I5(sum_2[23:23]),.LO(un36_prod_a_b_axb_22));
defparam desc951.INIT=64'h36C96C93C936936C;
  LUT6_L desc952(.I0(sum_0[8:8]),.I1(sum_0[9:9]),.I2(sum_1[20:20]),.I3(sum_1[21:21]),.I4(sum_2[20:20]),.I5(sum_2[21:21]),.LO(un36_prod_a_b_axb_20));
defparam desc952.INIT=64'h36C96C93C936936C;
  LUT6_L desc953(.I0(sum_0[0:0]),.I1(sum_1[11:11]),.I2(sum_1[12:12]),.I3(sum_2[11:11]),.I4(sum_2[12:12]),.I5(sum_3[23:23]),.LO(un36_prod_a_b_axb_11));
defparam desc953.INIT=64'h5A69A59669A5965A;
  LUT6_L desc954(.I0(sum_0[5:5]),.I1(sum_0[6:6]),.I2(sum_1[17:17]),.I3(sum_1[18:18]),.I4(sum_2[17:17]),.I5(sum_2[18:18]),.LO(un36_prod_a_b_axb_17));
defparam desc954.INIT=64'h36C96C93C936936C;
  LUT6_L desc955(.I0(sum_1[5:5]),.I1(sum_1[6:6]),.I2(sum_2[5:5]),.I3(sum_2[6:6]),.I4(sum_3[17:17]),.I5(sum_3[18:18]),.LO(un36_prod_a_b_axb_5));
defparam desc955.INIT=64'h36C96C93C936936C;
  LUT6_L desc956(.I0(sum_0[2:2]),.I1(sum_0[3:3]),.I2(sum_1[14:14]),.I3(sum_1[15:15]),.I4(sum_2[14:14]),.I5(sum_2[15:15]),.LO(un36_prod_a_b_axb_14));
defparam desc956.INIT=64'h36C96C93C936936C;
  LUT6 desc957(.I0(N_136_0),.I1(N_139_0),.I2(N_3281),.I3(N_3282),.I4(N_3293),.I5(N_3294),.O(un54_sum_axb_9));
defparam desc957.INIT=64'h36C96C93C936936C;
  LUT6 desc958(.I0(N_130_0),.I1(N_133_0),.I2(N_3279),.I3(N_3280),.I4(N_3291),.I5(N_3292),.O(un54_sum_axb_7));
defparam desc958.INIT=64'h36C96C93C936936C;
  LUT6_L desc959(.I0(sum_1[9:9]),.I1(sum_1[10:10]),.I2(sum_2[9:9]),.I3(sum_2[10:10]),.I4(sum_3[21:21]),.I5(sum_3[22:22]),.LO(un36_prod_a_b_axb_9));
defparam desc959.INIT=64'h36C96C93C936936C;
  LUT6_L desc960(.I0(sum_1[8:8]),.I1(sum_1[9:9]),.I2(sum_2[8:8]),.I3(sum_2[9:9]),.I4(sum_3[20:20]),.I5(sum_3[21:21]),.LO(un36_prod_a_b_axb_8));
defparam desc960.INIT=64'h36C96C93C936936C;
  LUT6 desc961(.I0(N_127_0),.I1(N_130_0),.I2(N_3278),.I3(N_3279),.I4(N_3290),.I5(N_3291),.O(un54_sum_axb_6));
defparam desc961.INIT=64'h36C96C93C936936C;
  LUT6 desc962(.I0(N_133_0),.I1(N_136_0),.I2(N_3280),.I3(N_3281),.I4(N_3292),.I5(N_3293),.O(un54_sum_axb_8));
defparam desc962.INIT=64'h36C96C93C936936C;
  LUT6 desc963(.I0(N_139_0),.I1(N_3282),.I2(N_3294),.I3(N_85_0),.I4(N_142_0),.I5(N_3283),.O(un54_sum_axb_10));
defparam desc963.INIT=64'h17E8E817E81717E8;
  LUT6_L desc964(.I0(sum_0[9:9]),.I1(sum_0[10:10]),.I2(sum_1[21:21]),.I3(sum_1[22:22]),.I4(sum_2[21:21]),.I5(sum_2[22:22]),.LO(un36_prod_a_b_axb_21));
defparam desc964.INIT=64'h36C96C93C936936C;
  LUT6_L desc965(.I0(sum_0[3:3]),.I1(sum_0[4:4]),.I2(sum_1[15:15]),.I3(sum_1[16:16]),.I4(sum_2[15:15]),.I5(sum_2[16:16]),.LO(un36_prod_a_b_axb_15));
defparam desc965.INIT=64'h36C96C93C936936C;
  LUT6 desc966(.I0(N_118_0),.I1(N_121_0),.I2(N_3276),.I3(N_3277),.I4(N_3288),.I5(N_3289),.O(un54_sum_axb_4));
defparam desc966.INIT=64'h36C96C93C936936C;
  LUT6 desc967(.I0(N_112_0),.I1(N_115_0),.I2(N_172_0),.I3(N_3274),.I4(N_3286),.I5(N_3287),.O(un54_sum_axb_2));
defparam desc967.INIT=64'h3C6969C3C396963C;
  LUT6_L desc968(.I0(sum_1[3:3]),.I1(sum_1[4:4]),.I2(sum_2[3:3]),.I3(sum_2[4:4]),.I4(sum_3[15:15]),.I5(sum_3[16:16]),.LO(un36_prod_a_b_axb_3));
defparam desc968.INIT=64'h36C96C93C936936C;
  LUT6_L desc969(.I0(sum_1[2:2]),.I1(sum_1[3:3]),.I2(sum_2[2:2]),.I3(sum_2[3:3]),.I4(sum_3[14:14]),.I5(sum_3[15:15]),.LO(un36_prod_a_b_axb_2));
defparam desc969.INIT=64'h36C96C93C936936C;
  LUT6_L desc970(.I0(sum_1[1:1]),.I1(sum_1[2:2]),.I2(sum_2[1:1]),.I3(sum_2[2:2]),.I4(sum_3[13:13]),.I5(sum_3[14:14]),.LO(un36_prod_a_b_axb_1));
defparam desc970.INIT=64'h36C96C93C936936C;
  LUT6 desc971(.I0(sum_1[0:0]),.I1(sum_2[0:0]),.I2(sum_3[12:12]),.I3(sum_1[1:1]),.I4(sum_2[1:1]),.I5(sum_3[13:13]),.O(mul_24_fract_48[13:13]));
defparam desc971.INIT=64'h17E8E817E81717E8;
  LUT6 desc972(.I0(N_106_0),.I1(N_3272),.I2(N_3284),.I3(N_109_0),.I4(N_3273),.I5(N_3285),.O(un54_sum[654:654]));
defparam desc972.INIT=64'h17E8E817E81717E8;
  LUT6_L desc973(.I0(sum_1[7:7]),.I1(sum_1[8:8]),.I2(sum_2[7:7]),.I3(sum_2[8:8]),.I4(sum_3[19:19]),.I5(sum_3[20:20]),.LO(un36_prod_a_b_axb_7));
defparam desc973.INIT=64'h36C96C93C936936C;
  LUT6 desc974(.I0(N_109_0),.I1(N_112_0),.I2(N_3273),.I3(N_3274),.I4(N_3285),.I5(N_3286),.O(un54_sum_axb_1));
defparam desc974.INIT=64'h36C96C93C936936C;
  LUT6 desc975(.I0(N_121_0),.I1(N_127_0),.I2(N_3277),.I3(N_3278),.I4(N_3289),.I5(N_3290),.O(un54_sum_axb_5));
defparam desc975.INIT=64'h36C96C93C936936C;
  LUT6 desc976(.I0(N_115_0),.I1(N_118_0),.I2(N_172_0),.I3(N_3276),.I4(N_3287),.I5(N_3288),.O(un54_sum_axb_3));
defparam desc976.INIT=64'h36C96C93C936936C;
  LUT1_L un36_prod_a_b_axb_34_cZ(.I0(sum_0[23:23]),.LO(un36_prod_a_b_axb_34));
defparam un36_prod_a_b_axb_34_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_33_cZ(.I0(sum_0[22:22]),.LO(un36_prod_a_b_axb_33));
defparam un36_prod_a_b_axb_33_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_32_cZ(.I0(sum_0[21:21]),.LO(un36_prod_a_b_axb_32));
defparam un36_prod_a_b_axb_32_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_31_cZ(.I0(sum_0[20:20]),.LO(un36_prod_a_b_axb_31));
defparam un36_prod_a_b_axb_31_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_30_cZ(.I0(sum_0[19:19]),.LO(un36_prod_a_b_axb_30));
defparam un36_prod_a_b_axb_30_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_29_cZ(.I0(sum_0[18:18]),.LO(un36_prod_a_b_axb_29));
defparam un36_prod_a_b_axb_29_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_28_cZ(.I0(sum_0[17:17]),.LO(un36_prod_a_b_axb_28));
defparam un36_prod_a_b_axb_28_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_27_cZ(.I0(sum_0[16:16]),.LO(un36_prod_a_b_axb_27));
defparam un36_prod_a_b_axb_27_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_26_cZ(.I0(sum_0[15:15]),.LO(un36_prod_a_b_axb_26));
defparam un36_prod_a_b_axb_26_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_25_cZ(.I0(sum_0[14:14]),.LO(un36_prod_a_b_axb_25));
defparam un36_prod_a_b_axb_25_cZ.INIT=2'h2;
  LUT1_L un36_prod_a_b_axb_24_cZ(.I0(sum_0[13:13]),.LO(un36_prod_a_b_axb_24));
defparam un36_prod_a_b_axb_24_cZ.INIT=2'h2;
  LUT3_L un36_prod_a_b(.I0(sum_1[0:0]),.I1(sum_2[0:0]),.I2(sum_3[12:12]),.LO(mul_24_fract_48[12:12]));
defparam un36_prod_a_b.INIT=8'h96;
  LUT6 desc977(.I0(prod2_0_2[17:17]),.I1(prod2_1_2[17:17]),.I2(prod2_2_2[17:17]),.I3(prod2_3_2[17:17]),.I4(count[1:1]),.I5(count[0:0]),.O(N_85_0));
defparam desc977.INIT=64'h0F0F5555333300FF;
  LUT6 desc978(.I0(prod2_0_3[6:6]),.I1(prod2_1_3[6:6]),.I2(prod2_2_3[6:6]),.I3(prod2_3_3[6:6]),.I4(count[1:1]),.I5(count[0:0]),.O(N_106_0));
defparam desc978.INIT=64'h0F0F5555333300FF;
  LUT6 desc979(.I0(prod2_0_3[7:7]),.I1(prod2_1_3[7:7]),.I2(prod2_2_3[7:7]),.I3(prod2_3_3[7:7]),.I4(count[1:1]),.I5(count[0:0]),.O(N_109_0));
defparam desc979.INIT=64'h0F0F5555333300FF;
  LUT6 desc980(.I0(prod2_0_3[8:8]),.I1(prod2_1_3[8:8]),.I2(prod2_2_3[8:8]),.I3(prod2_3_3[8:8]),.I4(count[1:1]),.I5(count[0:0]),.O(N_112_0));
defparam desc980.INIT=64'h0F0F5555333300FF;
  LUT6 desc981(.I0(prod2_0_3[9:9]),.I1(prod2_1_3[9:9]),.I2(prod2_2_3[9:9]),.I3(prod2_3_3[9:9]),.I4(count[1:1]),.I5(count[0:0]),.O(N_115_0));
defparam desc981.INIT=64'h0F0F5555333300FF;
  LUT6 desc982(.I0(prod2_0_3[10:10]),.I1(prod2_1_3[10:10]),.I2(prod2_2_3[10:10]),.I3(prod2_3_3[10:10]),.I4(count[1:1]),.I5(count[0:0]),.O(N_118_0));
defparam desc982.INIT=64'h0F0F5555333300FF;
  LUT6 desc983(.I0(prod2_0_3[11:11]),.I1(prod2_1_3[11:11]),.I2(prod2_2_3[11:11]),.I3(prod2_3_3[11:11]),.I4(count[1:1]),.I5(count[0:0]),.O(N_121_0));
defparam desc983.INIT=64'h0F0F5555333300FF;
  LUT6 desc984(.I0(prod2_0_0[12:12]),.I1(prod2_1_0[12:12]),.I2(prod2_2_0[12:12]),.I3(prod2_3_0[12:12]),.I4(count[1:1]),.I5(count[0:0]),.O(N_127_0));
defparam desc984.INIT=64'h0F0F5555333300FF;
  LUT6 desc985(.I0(prod2_0_0[13:13]),.I1(prod2_1_0[13:13]),.I2(prod2_2_0[13:13]),.I3(prod2_3_0[13:13]),.I4(count[1:1]),.I5(count[0:0]),.O(N_130_0));
defparam desc985.INIT=64'h0F0F5555333300FF;
  LUT6 desc986(.I0(prod2_0_0[14:14]),.I1(prod2_1_0[14:14]),.I2(prod2_2_0[14:14]),.I3(prod2_3_0[14:14]),.I4(count[1:1]),.I5(count[0:0]),.O(N_133_0));
defparam desc986.INIT=64'h0F0F5555333300FF;
  LUT6 desc987(.I0(prod2_0_0[15:15]),.I1(prod2_1_0[15:15]),.I2(prod2_2_0[15:15]),.I3(prod2_3_0[15:15]),.I4(count[1:1]),.I5(count[0:0]),.O(N_136_0));
defparam desc987.INIT=64'h0F0F5555333300FF;
  LUT6 desc988(.I0(prod2_0_0[16:16]),.I1(prod2_1_0[16:16]),.I2(prod2_2_0[16:16]),.I3(prod2_3_0[16:16]),.I4(count[1:1]),.I5(count[0:0]),.O(N_139_0));
defparam desc988.INIT=64'h0F0F5555333300FF;
  LUT6 desc989(.I0(prod2_0_0[17:17]),.I1(prod2_1_0[17:17]),.I2(prod2_2_0[17:17]),.I3(prod2_3_0[17:17]),.I4(count[1:1]),.I5(count[0:0]),.O(N_142_0));
defparam desc989.INIT=64'h0F0F5555333300FF;
  LUT6 desc990(.I0(prod2_0_1[6:6]),.I1(prod2_1_1[6:6]),.I2(prod2_2_1[6:6]),.I3(prod2_3_1[6:6]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3272));
defparam desc990.INIT=64'h0F0F5555333300FF;
  LUT6 desc991(.I0(prod2_0_1[7:7]),.I1(prod2_1_1[7:7]),.I2(prod2_2_1[7:7]),.I3(prod2_3_1[7:7]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3273));
defparam desc991.INIT=64'h0F0F5555333300FF;
  LUT6 desc992(.I0(prod2_0_1[8:8]),.I1(prod2_1_1[8:8]),.I2(prod2_2_1[8:8]),.I3(prod2_3_1[8:8]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3274));
defparam desc992.INIT=64'h0F0F5555333300FF;
  LUT6 desc993(.I0(prod2_0_1[9:9]),.I1(prod2_1_1[9:9]),.I2(prod2_2_1[9:9]),.I3(prod2_3_1[9:9]),.I4(count[1:1]),.I5(count[0:0]),.O(N_172_0));
defparam desc993.INIT=64'h0F0F5555333300FF;
  LUT6 desc994(.I0(prod2_0_1[10:10]),.I1(prod2_1_1[10:10]),.I2(prod2_2_1[10:10]),.I3(prod2_3_1[10:10]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3276));
defparam desc994.INIT=64'h0F0F5555333300FF;
  LUT6 desc995(.I0(prod2_0_1[11:11]),.I1(prod2_1_1[11:11]),.I2(prod2_2_1[11:11]),.I3(prod2_3_1[11:11]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3277));
defparam desc995.INIT=64'h0F0F5555333300FF;
  LUT6 desc996(.I0(prod2_0_1[12:12]),.I1(prod2_1_1[12:12]),.I2(prod2_2_1[12:12]),.I3(prod2_3_1[12:12]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3278));
defparam desc996.INIT=64'h0F0F5555333300FF;
  LUT6 desc997(.I0(prod2_0_1[13:13]),.I1(prod2_1_1[13:13]),.I2(prod2_2_1[13:13]),.I3(prod2_3_1[13:13]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3279));
defparam desc997.INIT=64'h0F0F5555333300FF;
  LUT6 desc998(.I0(prod2_0_1[14:14]),.I1(prod2_1_1[14:14]),.I2(prod2_2_1[14:14]),.I3(prod2_3_1[14:14]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3280));
defparam desc998.INIT=64'h0F0F5555333300FF;
  LUT6 desc999(.I0(prod2_0_1[15:15]),.I1(prod2_1_1[15:15]),.I2(prod2_2_1[15:15]),.I3(prod2_3_1[15:15]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3281));
defparam desc999.INIT=64'h0F0F5555333300FF;
  LUT6 desc1000(.I0(prod2_0_1[16:16]),.I1(prod2_1_1[16:16]),.I2(prod2_2_1[16:16]),.I3(prod2_3_1[16:16]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3282));
defparam desc1000.INIT=64'h0F0F5555333300FF;
  LUT6 desc1001(.I0(prod2_0_1[17:17]),.I1(prod2_1_1[17:17]),.I2(prod2_2_1[17:17]),.I3(prod2_3_1[17:17]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3283));
defparam desc1001.INIT=64'h0F0F5555333300FF;
  LUT6 desc1002(.I0(prod2_0_2[6:6]),.I1(prod2_1_2[6:6]),.I2(prod2_2_2[6:6]),.I3(prod2_3_2[6:6]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3284));
defparam desc1002.INIT=64'h0F0F5555333300FF;
  LUT6 desc1003(.I0(prod2_0_2[7:7]),.I1(prod2_1_2[7:7]),.I2(prod2_2_2[7:7]),.I3(prod2_3_2[7:7]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3285));
defparam desc1003.INIT=64'h0F0F5555333300FF;
  LUT6 desc1004(.I0(prod2_0_2[8:8]),.I1(prod2_1_2[8:8]),.I2(prod2_2_2[8:8]),.I3(prod2_3_2[8:8]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3286));
defparam desc1004.INIT=64'h0F0F5555333300FF;
  LUT6 desc1005(.I0(prod2_0_2[9:9]),.I1(prod2_1_2[9:9]),.I2(prod2_2_2[9:9]),.I3(prod2_3_2[9:9]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3287));
defparam desc1005.INIT=64'h0F0F5555333300FF;
  LUT6 desc1006(.I0(prod2_0_2[10:10]),.I1(prod2_1_2[10:10]),.I2(prod2_2_2[10:10]),.I3(prod2_3_2[10:10]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3288));
defparam desc1006.INIT=64'h0F0F5555333300FF;
  LUT6 desc1007(.I0(prod2_0_2[11:11]),.I1(prod2_1_2[11:11]),.I2(prod2_2_2[11:11]),.I3(prod2_3_2[11:11]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3289));
defparam desc1007.INIT=64'h0F0F5555333300FF;
  LUT6 desc1008(.I0(prod2_0_2[12:12]),.I1(prod2_1_2[12:12]),.I2(prod2_2_2[12:12]),.I3(prod2_3_2[12:12]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3290));
defparam desc1008.INIT=64'h0F0F5555333300FF;
  LUT6 desc1009(.I0(prod2_0_2[13:13]),.I1(prod2_1_2[13:13]),.I2(prod2_2_2[13:13]),.I3(prod2_3_2[13:13]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3291));
defparam desc1009.INIT=64'h0F0F5555333300FF;
  LUT6 desc1010(.I0(prod2_0_2[14:14]),.I1(prod2_1_2[14:14]),.I2(prod2_2_2[14:14]),.I3(prod2_3_2[14:14]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3292));
defparam desc1010.INIT=64'h0F0F5555333300FF;
  LUT6 desc1011(.I0(prod2_0_2[15:15]),.I1(prod2_1_2[15:15]),.I2(prod2_2_2[15:15]),.I3(prod2_3_2[15:15]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3293));
defparam desc1011.INIT=64'h0F0F5555333300FF;
  LUT6 desc1012(.I0(prod2_0_2[16:16]),.I1(prod2_1_2[16:16]),.I2(prod2_2_2[16:16]),.I3(prod2_3_2[16:16]),.I4(count[1:1]),.I5(count[0:0]),.O(N_3294));
defparam desc1012.INIT=64'h0F0F5555333300FF;
  LUT6 un54_sum_axb_16_cZ(.I0(prod2_0_0[23:23]),.I1(prod2_1_0[23:23]),.I2(prod2_2_0[23:23]),.I3(prod2_3_0[23:23]),.I4(count[1:1]),.I5(count[0:0]),.O(un54_sum_axb_16));
defparam un54_sum_axb_16_cZ.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 un54_sum_axb_15_cZ(.I0(prod2_0_0[22:22]),.I1(prod2_1_0[22:22]),.I2(prod2_2_0[22:22]),.I3(prod2_3_0[22:22]),.I4(count[1:1]),.I5(count[0:0]),.O(un54_sum_axb_15));
defparam un54_sum_axb_15_cZ.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 un54_sum_axb_14_cZ(.I0(prod2_0_0[21:21]),.I1(prod2_1_0[21:21]),.I2(prod2_2_0[21:21]),.I3(prod2_3_0[21:21]),.I4(count[1:1]),.I5(count[0:0]),.O(un54_sum_axb_14));
defparam un54_sum_axb_14_cZ.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 un54_sum_axb_13_cZ(.I0(prod2_0_0[20:20]),.I1(prod2_1_0[20:20]),.I2(prod2_2_0[20:20]),.I3(prod2_3_0[20:20]),.I4(count[1:1]),.I5(count[0:0]),.O(un54_sum_axb_13));
defparam un54_sum_axb_13_cZ.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 un54_sum_axb_12_cZ(.I0(prod2_0_0[19:19]),.I1(prod2_1_0[19:19]),.I2(prod2_2_0[19:19]),.I3(prod2_3_0[19:19]),.I4(count[1:1]),.I5(count[0:0]),.O(un54_sum_axb_12));
defparam un54_sum_axb_12_cZ.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1013(.I0(prod2_0_0[18:18]),.I1(prod2_1_0[18:18]),.I2(prod2_2_0[18:18]),.I3(prod2_3_0[18:18]),.I4(count[1:1]),.I5(count[0:0]),.O(N_145_0_i));
defparam desc1013.INIT=64'hF0F0AAAACCCCFF00;
  LUT4_L un36_prod_a_b_axb_23_cZ(.I0(sum_0[12:12]),.I1(sum_0[11:11]),.I2(sum_1[23:23]),.I3(sum_2[23:23]),.LO(un36_prod_a_b_axb_23));
defparam un36_prod_a_b_axb_23_cZ.INIT=16'h566A;
  LUT6 desc1014(.I0(prod2_0_3[0:0]),.I1(prod2_1_3[0:0]),.I2(prod2_2_3[0:0]),.I3(prod2_3_3[0:0]),.I4(count[1:1]),.I5(count[0:0]),.O(N_88_0_i));
defparam desc1014.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1015(.I0(prod2_0_3[1:1]),.I1(prod2_1_3[1:1]),.I2(prod2_2_3[1:1]),.I3(prod2_3_3[1:1]),.I4(count[1:1]),.I5(count[0:0]),.O(N_91_0_i));
defparam desc1015.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1016(.I0(prod2_0_3[2:2]),.I1(prod2_1_3[2:2]),.I2(prod2_2_3[2:2]),.I3(prod2_3_3[2:2]),.I4(count[1:1]),.I5(count[0:0]),.O(N_94_0_i));
defparam desc1016.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1017(.I0(prod2_0_3[3:3]),.I1(prod2_1_3[3:3]),.I2(prod2_2_3[3:3]),.I3(prod2_3_3[3:3]),.I4(count[1:1]),.I5(count[0:0]),.O(N_97_0_i));
defparam desc1017.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1018(.I0(prod2_0_3[4:4]),.I1(prod2_1_3[4:4]),.I2(prod2_2_3[4:4]),.I3(prod2_3_3[4:4]),.I4(count[1:1]),.I5(count[0:0]),.O(N_100_0_i));
defparam desc1018.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1019(.I0(prod2_0_3[5:5]),.I1(prod2_1_3[5:5]),.I2(prod2_2_3[5:5]),.I3(prod2_3_3[5:5]),.I4(count[1:1]),.I5(count[0:0]),.O(N_103_0_i));
defparam desc1019.INIT=64'hF0F0AAAACCCCFF00;
  LUT3 un54_sum_cZ(.I0(N_106_0),.I1(N_3272),.I2(N_3284),.O(un54_sum[653:653]));
defparam un54_sum_cZ.INIT=8'h69;
  LUT3 un36_prod_a_b_cry_0_RNO_cZ(.I0(sum_1[1:1]),.I1(sum_2[1:1]),.I2(sum_3[13:13]),.O(un36_prod_a_b_cry_0_RNO));
defparam un36_prod_a_b_cry_0_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_1_RNO_cZ(.I0(sum_1[2:2]),.I1(sum_2[2:2]),.I2(sum_3[14:14]),.O(un36_prod_a_b_cry_1_RNO));
defparam un36_prod_a_b_cry_1_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_2_RNO_cZ(.I0(sum_1[3:3]),.I1(sum_2[3:3]),.I2(sum_3[15:15]),.O(un36_prod_a_b_cry_2_RNO));
defparam un36_prod_a_b_cry_2_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_3_RNO_cZ(.I0(sum_1[4:4]),.I1(sum_2[4:4]),.I2(sum_3[16:16]),.O(un36_prod_a_b_cry_3_RNO));
defparam un36_prod_a_b_cry_3_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_4_RNO_cZ(.I0(sum_1[5:5]),.I1(sum_2[5:5]),.I2(sum_3[17:17]),.O(un36_prod_a_b_cry_4_RNO));
defparam un36_prod_a_b_cry_4_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_5_RNO_cZ(.I0(sum_1[6:6]),.I1(sum_2[6:6]),.I2(sum_3[18:18]),.O(un36_prod_a_b_cry_5_RNO));
defparam un36_prod_a_b_cry_5_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_6_RNO_cZ(.I0(sum_1[7:7]),.I1(sum_2[7:7]),.I2(sum_3[19:19]),.O(un36_prod_a_b_cry_6_RNO));
defparam un36_prod_a_b_cry_6_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_7_RNO_cZ(.I0(sum_1[8:8]),.I1(sum_2[8:8]),.I2(sum_3[20:20]),.O(un36_prod_a_b_cry_7_RNO));
defparam un36_prod_a_b_cry_7_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_8_RNO_cZ(.I0(sum_1[9:9]),.I1(sum_2[9:9]),.I2(sum_3[21:21]),.O(un36_prod_a_b_cry_8_RNO));
defparam un36_prod_a_b_cry_8_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_9_RNO_cZ(.I0(sum_1[10:10]),.I1(sum_2[10:10]),.I2(sum_3[22:22]),.O(un36_prod_a_b_cry_9_RNO));
defparam un36_prod_a_b_cry_9_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_10_RNO_cZ(.I0(sum_1[11:11]),.I1(sum_2[11:11]),.I2(sum_3[23:23]),.O(un36_prod_a_b_cry_10_RNO));
defparam un36_prod_a_b_cry_10_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_11_RNO_cZ(.I0(sum_0[0:0]),.I1(sum_1[12:12]),.I2(sum_2[12:12]),.O(un36_prod_a_b_cry_11_RNO));
defparam un36_prod_a_b_cry_11_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_12_RNO_cZ(.I0(sum_0[1:1]),.I1(sum_1[13:13]),.I2(sum_2[13:13]),.O(un36_prod_a_b_cry_12_RNO));
defparam un36_prod_a_b_cry_12_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_13_RNO_cZ(.I0(sum_0[2:2]),.I1(sum_1[14:14]),.I2(sum_2[14:14]),.O(un36_prod_a_b_cry_13_RNO));
defparam un36_prod_a_b_cry_13_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_14_RNO_cZ(.I0(sum_0[3:3]),.I1(sum_1[15:15]),.I2(sum_2[15:15]),.O(un36_prod_a_b_cry_14_RNO));
defparam un36_prod_a_b_cry_14_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_15_RNO_cZ(.I0(sum_0[4:4]),.I1(sum_1[16:16]),.I2(sum_2[16:16]),.O(un36_prod_a_b_cry_15_RNO));
defparam un36_prod_a_b_cry_15_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_16_RNO_cZ(.I0(sum_0[5:5]),.I1(sum_1[17:17]),.I2(sum_2[17:17]),.O(un36_prod_a_b_cry_16_RNO));
defparam un36_prod_a_b_cry_16_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_17_RNO_cZ(.I0(sum_0[6:6]),.I1(sum_1[18:18]),.I2(sum_2[18:18]),.O(un36_prod_a_b_cry_17_RNO));
defparam un36_prod_a_b_cry_17_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_18_RNO_cZ(.I0(sum_0[7:7]),.I1(sum_1[19:19]),.I2(sum_2[19:19]),.O(un36_prod_a_b_cry_18_RNO));
defparam un36_prod_a_b_cry_18_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_19_RNO_cZ(.I0(sum_0[8:8]),.I1(sum_1[20:20]),.I2(sum_2[20:20]),.O(un36_prod_a_b_cry_19_RNO));
defparam un36_prod_a_b_cry_19_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_20_RNO_cZ(.I0(sum_0[9:9]),.I1(sum_1[21:21]),.I2(sum_2[21:21]),.O(un36_prod_a_b_cry_20_RNO));
defparam un36_prod_a_b_cry_20_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_21_RNO_cZ(.I0(sum_0[10:10]),.I1(sum_1[22:22]),.I2(sum_2[22:22]),.O(un36_prod_a_b_cry_21_RNO));
defparam un36_prod_a_b_cry_21_RNO_cZ.INIT=8'h96;
  LUT3 un36_prod_a_b_cry_22_RNO_cZ(.I0(sum_0[11:11]),.I1(sum_1[23:23]),.I2(sum_2[23:23]),.O(un36_prod_a_b_cry_22_RNO));
defparam un36_prod_a_b_cry_22_RNO_cZ.INIT=8'h96;
  LUT3 un54_sum_cry_0_RNO_cZ(.I0(N_109_0),.I1(N_3273),.I2(N_3285),.O(un54_sum_cry_0_RNO));
defparam un54_sum_cry_0_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_1_RNO_cZ(.I0(N_112_0),.I1(N_3274),.I2(N_3286),.O(un54_sum_cry_1_RNO));
defparam un54_sum_cry_1_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_2_RNO_cZ(.I0(N_115_0),.I1(N_172_0),.I2(N_3287),.O(un54_sum_cry_2_RNO));
defparam un54_sum_cry_2_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_3_RNO_cZ(.I0(N_118_0),.I1(N_3276),.I2(N_3288),.O(un54_sum_cry_3_RNO));
defparam un54_sum_cry_3_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_4_RNO_cZ(.I0(N_121_0),.I1(N_3277),.I2(N_3289),.O(un54_sum_cry_4_RNO));
defparam un54_sum_cry_4_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_5_RNO_cZ(.I0(N_127_0),.I1(N_3278),.I2(N_3290),.O(un54_sum_cry_5_RNO));
defparam un54_sum_cry_5_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_6_RNO_cZ(.I0(N_130_0),.I1(N_3279),.I2(N_3291),.O(un54_sum_cry_6_RNO));
defparam un54_sum_cry_6_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_7_RNO_cZ(.I0(N_133_0),.I1(N_3280),.I2(N_3292),.O(un54_sum_cry_7_RNO));
defparam un54_sum_cry_7_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_8_RNO_cZ(.I0(N_136_0),.I1(N_3281),.I2(N_3293),.O(un54_sum_cry_8_RNO));
defparam un54_sum_cry_8_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_9_RNO_cZ(.I0(N_139_0),.I1(N_3282),.I2(N_3294),.O(un54_sum_cry_9_RNO));
defparam un54_sum_cry_9_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_10_RNO_cZ(.I0(N_85_0),.I1(N_142_0),.I2(N_3283),.O(un54_sum_cry_10_RNO));
defparam un54_sum_cry_10_RNO_cZ.INIT=8'h69;
  LUT3 un54_sum_cry_11_RNO_cZ(.I0(N_85_0),.I1(N_142_0),.I2(N_3283),.O(un54_sum_cry_11_RNO));
defparam un54_sum_cry_11_RNO_cZ.INIT=8'h17;
  XORCY un54_sum_s_16(.LI(un54_sum_axb_16),.CI(un54_sum_cry_15),.O(un54_sum[670:670]));
  XORCY un54_sum_s_15(.LI(un54_sum_axb_15),.CI(un54_sum_cry_14),.O(un54_sum[669:669]));
  MUXCY_L un54_sum_cry_15_cZ(.DI(GND),.CI(un54_sum_cry_14),.S(un54_sum_axb_15),.LO(un54_sum_cry_15));
  XORCY un54_sum_s_14(.LI(un54_sum_axb_14),.CI(un54_sum_cry_13),.O(un54_sum[668:668]));
  MUXCY_L un54_sum_cry_14_cZ(.DI(GND),.CI(un54_sum_cry_13),.S(un54_sum_axb_14),.LO(un54_sum_cry_14));
  XORCY un54_sum_s_13(.LI(un54_sum_axb_13),.CI(un54_sum_cry_12),.O(un54_sum[667:667]));
  MUXCY_L un54_sum_cry_13_cZ(.DI(GND),.CI(un54_sum_cry_12),.S(un54_sum_axb_13),.LO(un54_sum_cry_13));
  XORCY un54_sum_s_12(.LI(un54_sum_axb_12),.CI(un54_sum_cry_11),.O(un54_sum[666:666]));
  MUXCY_L un54_sum_cry_12_cZ(.DI(GND),.CI(un54_sum_cry_11),.S(un54_sum_axb_12),.LO(un54_sum_cry_12));
  XORCY un54_sum_s_11(.LI(un54_sum_axb_11),.CI(un54_sum_cry_10),.O(un54_sum[665:665]));
  MUXCY_L un54_sum_cry_11_cZ(.DI(un54_sum_cry_11_RNO),.CI(un54_sum_cry_10),.S(un54_sum_axb_11),.LO(un54_sum_cry_11));
  XORCY un54_sum_s_10(.LI(un54_sum_axb_10),.CI(un54_sum_cry_9),.O(un54_sum[664:664]));
  MUXCY_L un54_sum_cry_10_cZ(.DI(un54_sum_cry_10_RNO),.CI(un54_sum_cry_9),.S(un54_sum_axb_10),.LO(un54_sum_cry_10));
  XORCY un54_sum_s_9(.LI(un54_sum_axb_9),.CI(un54_sum_cry_8),.O(un54_sum[663:663]));
  MUXCY_L un54_sum_cry_9_cZ(.DI(un54_sum_cry_9_RNO),.CI(un54_sum_cry_8),.S(un54_sum_axb_9),.LO(un54_sum_cry_9));
  XORCY un54_sum_s_8(.LI(un54_sum_axb_8),.CI(un54_sum_cry_7),.O(un54_sum[662:662]));
  MUXCY_L un54_sum_cry_8_cZ(.DI(un54_sum_cry_8_RNO),.CI(un54_sum_cry_7),.S(un54_sum_axb_8),.LO(un54_sum_cry_8));
  XORCY un54_sum_s_7(.LI(un54_sum_axb_7),.CI(un54_sum_cry_6),.O(un54_sum[661:661]));
  MUXCY_L un54_sum_cry_7_cZ(.DI(un54_sum_cry_7_RNO),.CI(un54_sum_cry_6),.S(un54_sum_axb_7),.LO(un54_sum_cry_7));
  XORCY un54_sum_s_6(.LI(un54_sum_axb_6),.CI(un54_sum_cry_5),.O(un54_sum[660:660]));
  MUXCY_L un54_sum_cry_6_cZ(.DI(un54_sum_cry_6_RNO),.CI(un54_sum_cry_5),.S(un54_sum_axb_6),.LO(un54_sum_cry_6));
  XORCY un54_sum_s_5(.LI(un54_sum_axb_5),.CI(un54_sum_cry_4),.O(un54_sum[659:659]));
  MUXCY_L un54_sum_cry_5_cZ(.DI(un54_sum_cry_5_RNO),.CI(un54_sum_cry_4),.S(un54_sum_axb_5),.LO(un54_sum_cry_5));
  XORCY un54_sum_s_4(.LI(un54_sum_axb_4),.CI(un54_sum_cry_3),.O(un54_sum[658:658]));
  MUXCY_L un54_sum_cry_4_cZ(.DI(un54_sum_cry_4_RNO),.CI(un54_sum_cry_3),.S(un54_sum_axb_4),.LO(un54_sum_cry_4));
  XORCY un54_sum_s_3(.LI(un54_sum_axb_3),.CI(un54_sum_cry_2),.O(un54_sum[657:657]));
  MUXCY_L un54_sum_cry_3_cZ(.DI(un54_sum_cry_3_RNO),.CI(un54_sum_cry_2),.S(un54_sum_axb_3),.LO(un54_sum_cry_3));
  XORCY un54_sum_s_2(.LI(un54_sum_axb_2),.CI(un54_sum_cry_1),.O(un54_sum[656:656]));
  MUXCY_L un54_sum_cry_2_cZ(.DI(un54_sum_cry_2_RNO),.CI(un54_sum_cry_1),.S(un54_sum_axb_2),.LO(un54_sum_cry_2));
  XORCY un54_sum_s_1(.LI(un54_sum_axb_1),.CI(un54_sum_cry_0),.O(un54_sum[655:655]));
  MUXCY_L un54_sum_cry_1_cZ(.DI(un54_sum_cry_1_RNO),.CI(un54_sum_cry_0),.S(un54_sum_axb_1),.LO(un54_sum_cry_1));
  MUXCY_L un54_sum_cry_0_cZ(.DI(un54_sum_cry_0_RNO),.CI(GND),.S(un54_sum[654:654]),.LO(un54_sum_cry_0));
  XORCY un36_prod_a_b_s_34(.LI(un36_prod_a_b_axb_34),.CI(un36_prod_a_b_cry_33),.O(mul_24_fract_48[47:47]));
  XORCY un36_prod_a_b_s_33(.LI(un36_prod_a_b_axb_33),.CI(un36_prod_a_b_cry_32),.O(mul_24_fract_48[46:46]));
  MUXCY_L un36_prod_a_b_cry_33_cZ(.DI(GND),.CI(un36_prod_a_b_cry_32),.S(un36_prod_a_b_axb_33),.LO(un36_prod_a_b_cry_33));
  XORCY un36_prod_a_b_s_32(.LI(un36_prod_a_b_axb_32),.CI(un36_prod_a_b_cry_31),.O(mul_24_fract_48[45:45]));
  MUXCY_L un36_prod_a_b_cry_32_cZ(.DI(GND),.CI(un36_prod_a_b_cry_31),.S(un36_prod_a_b_axb_32),.LO(un36_prod_a_b_cry_32));
  XORCY un36_prod_a_b_s_31(.LI(un36_prod_a_b_axb_31),.CI(un36_prod_a_b_cry_30),.O(mul_24_fract_48[44:44]));
  MUXCY_L un36_prod_a_b_cry_31_cZ(.DI(GND),.CI(un36_prod_a_b_cry_30),.S(un36_prod_a_b_axb_31),.LO(un36_prod_a_b_cry_31));
  XORCY un36_prod_a_b_s_30(.LI(un36_prod_a_b_axb_30),.CI(un36_prod_a_b_cry_29),.O(mul_24_fract_48[43:43]));
  MUXCY_L un36_prod_a_b_cry_30_cZ(.DI(GND),.CI(un36_prod_a_b_cry_29),.S(un36_prod_a_b_axb_30),.LO(un36_prod_a_b_cry_30));
  XORCY un36_prod_a_b_s_29(.LI(un36_prod_a_b_axb_29),.CI(un36_prod_a_b_cry_28),.O(mul_24_fract_48[42:42]));
  MUXCY_L un36_prod_a_b_cry_29_cZ(.DI(GND),.CI(un36_prod_a_b_cry_28),.S(un36_prod_a_b_axb_29),.LO(un36_prod_a_b_cry_29));
  XORCY un36_prod_a_b_s_28(.LI(un36_prod_a_b_axb_28),.CI(un36_prod_a_b_cry_27),.O(mul_24_fract_48[41:41]));
  MUXCY_L un36_prod_a_b_cry_28_cZ(.DI(GND),.CI(un36_prod_a_b_cry_27),.S(un36_prod_a_b_axb_28),.LO(un36_prod_a_b_cry_28));
  XORCY un36_prod_a_b_s_27(.LI(un36_prod_a_b_axb_27),.CI(un36_prod_a_b_cry_26),.O(mul_24_fract_48[40:40]));
  MUXCY_L un36_prod_a_b_cry_27_cZ(.DI(GND),.CI(un36_prod_a_b_cry_26),.S(un36_prod_a_b_axb_27),.LO(un36_prod_a_b_cry_27));
  XORCY un36_prod_a_b_s_26(.LI(un36_prod_a_b_axb_26),.CI(un36_prod_a_b_cry_25),.O(mul_24_fract_48[39:39]));
  MUXCY_L un36_prod_a_b_cry_26_cZ(.DI(GND),.CI(un36_prod_a_b_cry_25),.S(un36_prod_a_b_axb_26),.LO(un36_prod_a_b_cry_26));
  XORCY un36_prod_a_b_s_25(.LI(un36_prod_a_b_axb_25),.CI(un36_prod_a_b_cry_24),.O(mul_24_fract_48[38:38]));
  MUXCY_L un36_prod_a_b_cry_25_cZ(.DI(GND),.CI(un36_prod_a_b_cry_24),.S(un36_prod_a_b_axb_25),.LO(un36_prod_a_b_cry_25));
  XORCY un36_prod_a_b_s_24(.LI(un36_prod_a_b_axb_24),.CI(un36_prod_a_b_cry_23),.O(mul_24_fract_48[37:37]));
  MUXCY_L un36_prod_a_b_cry_24_cZ(.DI(GND),.CI(un36_prod_a_b_cry_23),.S(un36_prod_a_b_axb_24),.LO(un36_prod_a_b_cry_24));
  XORCY un36_prod_a_b_s_23(.LI(un36_prod_a_b_axb_23),.CI(un36_prod_a_b_cry_22),.O(mul_24_fract_48[36:36]));
  MUXCY_L un36_prod_a_b_cry_23_cZ(.DI(sum_0[12:12]),.CI(un36_prod_a_b_cry_22),.S(un36_prod_a_b_axb_23),.LO(un36_prod_a_b_cry_23));
  XORCY un36_prod_a_b_s_22(.LI(un36_prod_a_b_axb_22),.CI(un36_prod_a_b_cry_21),.O(mul_24_fract_48[35:35]));
  MUXCY_L un36_prod_a_b_cry_22_cZ(.DI(un36_prod_a_b_cry_22_RNO),.CI(un36_prod_a_b_cry_21),.S(un36_prod_a_b_axb_22),.LO(un36_prod_a_b_cry_22));
  XORCY un36_prod_a_b_s_21(.LI(un36_prod_a_b_axb_21),.CI(un36_prod_a_b_cry_20),.O(mul_24_fract_48[34:34]));
  MUXCY_L un36_prod_a_b_cry_21_cZ(.DI(un36_prod_a_b_cry_21_RNO),.CI(un36_prod_a_b_cry_20),.S(un36_prod_a_b_axb_21),.LO(un36_prod_a_b_cry_21));
  XORCY un36_prod_a_b_s_20(.LI(un36_prod_a_b_axb_20),.CI(un36_prod_a_b_cry_19),.O(mul_24_fract_48[33:33]));
  MUXCY_L un36_prod_a_b_cry_20_cZ(.DI(un36_prod_a_b_cry_20_RNO),.CI(un36_prod_a_b_cry_19),.S(un36_prod_a_b_axb_20),.LO(un36_prod_a_b_cry_20));
  XORCY un36_prod_a_b_s_19(.LI(un36_prod_a_b_axb_19),.CI(un36_prod_a_b_cry_18),.O(mul_24_fract_48[32:32]));
  MUXCY_L un36_prod_a_b_cry_19_cZ(.DI(un36_prod_a_b_cry_19_RNO),.CI(un36_prod_a_b_cry_18),.S(un36_prod_a_b_axb_19),.LO(un36_prod_a_b_cry_19));
  XORCY un36_prod_a_b_s_18(.LI(un36_prod_a_b_axb_18),.CI(un36_prod_a_b_cry_17),.O(mul_24_fract_48[31:31]));
  MUXCY_L un36_prod_a_b_cry_18_cZ(.DI(un36_prod_a_b_cry_18_RNO),.CI(un36_prod_a_b_cry_17),.S(un36_prod_a_b_axb_18),.LO(un36_prod_a_b_cry_18));
  XORCY un36_prod_a_b_s_17(.LI(un36_prod_a_b_axb_17),.CI(un36_prod_a_b_cry_16),.O(mul_24_fract_48[30:30]));
  MUXCY_L un36_prod_a_b_cry_17_cZ(.DI(un36_prod_a_b_cry_17_RNO),.CI(un36_prod_a_b_cry_16),.S(un36_prod_a_b_axb_17),.LO(un36_prod_a_b_cry_17));
  XORCY un36_prod_a_b_s_16(.LI(un36_prod_a_b_axb_16),.CI(un36_prod_a_b_cry_15),.O(mul_24_fract_48[29:29]));
  MUXCY_L un36_prod_a_b_cry_16_cZ(.DI(un36_prod_a_b_cry_16_RNO),.CI(un36_prod_a_b_cry_15),.S(un36_prod_a_b_axb_16),.LO(un36_prod_a_b_cry_16));
  XORCY un36_prod_a_b_s_15(.LI(un36_prod_a_b_axb_15),.CI(un36_prod_a_b_cry_14),.O(mul_24_fract_48[28:28]));
  MUXCY_L un36_prod_a_b_cry_15_cZ(.DI(un36_prod_a_b_cry_15_RNO),.CI(un36_prod_a_b_cry_14),.S(un36_prod_a_b_axb_15),.LO(un36_prod_a_b_cry_15));
  XORCY un36_prod_a_b_s_14(.LI(un36_prod_a_b_axb_14),.CI(un36_prod_a_b_cry_13),.O(mul_24_fract_48[27:27]));
  MUXCY_L un36_prod_a_b_cry_14_cZ(.DI(un36_prod_a_b_cry_14_RNO),.CI(un36_prod_a_b_cry_13),.S(un36_prod_a_b_axb_14),.LO(un36_prod_a_b_cry_14));
  XORCY un36_prod_a_b_s_13(.LI(un36_prod_a_b_axb_13),.CI(un36_prod_a_b_cry_12),.O(mul_24_fract_48[26:26]));
  MUXCY_L un36_prod_a_b_cry_13_cZ(.DI(un36_prod_a_b_cry_13_RNO),.CI(un36_prod_a_b_cry_12),.S(un36_prod_a_b_axb_13),.LO(un36_prod_a_b_cry_13));
  XORCY un36_prod_a_b_s_12(.LI(un36_prod_a_b_axb_12),.CI(un36_prod_a_b_cry_11),.O(mul_24_fract_48[25:25]));
  MUXCY_L un36_prod_a_b_cry_12_cZ(.DI(un36_prod_a_b_cry_12_RNO),.CI(un36_prod_a_b_cry_11),.S(un36_prod_a_b_axb_12),.LO(un36_prod_a_b_cry_12));
  XORCY un36_prod_a_b_s_11(.LI(un36_prod_a_b_axb_11),.CI(un36_prod_a_b_cry_10),.O(mul_24_fract_48[24:24]));
  MUXCY_L un36_prod_a_b_cry_11_cZ(.DI(un36_prod_a_b_cry_11_RNO),.CI(un36_prod_a_b_cry_10),.S(un36_prod_a_b_axb_11),.LO(un36_prod_a_b_cry_11));
  XORCY un36_prod_a_b_s_10(.LI(un36_prod_a_b_axb_10),.CI(un36_prod_a_b_cry_9),.O(mul_24_fract_48[23:23]));
  MUXCY_L un36_prod_a_b_cry_10_cZ(.DI(un36_prod_a_b_cry_10_RNO),.CI(un36_prod_a_b_cry_9),.S(un36_prod_a_b_axb_10),.LO(un36_prod_a_b_cry_10));
  XORCY un36_prod_a_b_s_9(.LI(un36_prod_a_b_axb_9),.CI(un36_prod_a_b_cry_8),.O(mul_24_fract_48[22:22]));
  MUXCY_L un36_prod_a_b_cry_9_cZ(.DI(un36_prod_a_b_cry_9_RNO),.CI(un36_prod_a_b_cry_8),.S(un36_prod_a_b_axb_9),.LO(un36_prod_a_b_cry_9));
  XORCY un36_prod_a_b_s_8(.LI(un36_prod_a_b_axb_8),.CI(un36_prod_a_b_cry_7),.O(mul_24_fract_48[21:21]));
  MUXCY_L un36_prod_a_b_cry_8_cZ(.DI(un36_prod_a_b_cry_8_RNO),.CI(un36_prod_a_b_cry_7),.S(un36_prod_a_b_axb_8),.LO(un36_prod_a_b_cry_8));
  XORCY un36_prod_a_b_s_7(.LI(un36_prod_a_b_axb_7),.CI(un36_prod_a_b_cry_6),.O(mul_24_fract_48[20:20]));
  MUXCY_L un36_prod_a_b_cry_7_cZ(.DI(un36_prod_a_b_cry_7_RNO),.CI(un36_prod_a_b_cry_6),.S(un36_prod_a_b_axb_7),.LO(un36_prod_a_b_cry_7));
  XORCY un36_prod_a_b_s_6(.LI(un36_prod_a_b_axb_6),.CI(un36_prod_a_b_cry_5),.O(mul_24_fract_48[19:19]));
  MUXCY_L un36_prod_a_b_cry_6_cZ(.DI(un36_prod_a_b_cry_6_RNO),.CI(un36_prod_a_b_cry_5),.S(un36_prod_a_b_axb_6),.LO(un36_prod_a_b_cry_6));
  XORCY un36_prod_a_b_s_5(.LI(un36_prod_a_b_axb_5),.CI(un36_prod_a_b_cry_4),.O(mul_24_fract_48[18:18]));
  MUXCY_L un36_prod_a_b_cry_5_cZ(.DI(un36_prod_a_b_cry_5_RNO),.CI(un36_prod_a_b_cry_4),.S(un36_prod_a_b_axb_5),.LO(un36_prod_a_b_cry_5));
  XORCY un36_prod_a_b_s_4(.LI(un36_prod_a_b_axb_4),.CI(un36_prod_a_b_cry_3),.O(mul_24_fract_48[17:17]));
  MUXCY_L un36_prod_a_b_cry_4_cZ(.DI(un36_prod_a_b_cry_4_RNO),.CI(un36_prod_a_b_cry_3),.S(un36_prod_a_b_axb_4),.LO(un36_prod_a_b_cry_4));
  XORCY un36_prod_a_b_s_3(.LI(un36_prod_a_b_axb_3),.CI(un36_prod_a_b_cry_2),.O(mul_24_fract_48[16:16]));
  MUXCY_L un36_prod_a_b_cry_3_cZ(.DI(un36_prod_a_b_cry_3_RNO),.CI(un36_prod_a_b_cry_2),.S(un36_prod_a_b_axb_3),.LO(un36_prod_a_b_cry_3));
  XORCY un36_prod_a_b_s_2(.LI(un36_prod_a_b_axb_2),.CI(un36_prod_a_b_cry_1),.O(mul_24_fract_48[15:15]));
  MUXCY_L un36_prod_a_b_cry_2_cZ(.DI(un36_prod_a_b_cry_2_RNO),.CI(un36_prod_a_b_cry_1),.S(un36_prod_a_b_axb_2),.LO(un36_prod_a_b_cry_2));
  XORCY un36_prod_a_b_s_1(.LI(un36_prod_a_b_axb_1),.CI(un36_prod_a_b_cry_0),.O(mul_24_fract_48[14:14]));
  MUXCY_L un36_prod_a_b_cry_1_cZ(.DI(un36_prod_a_b_cry_1_RNO),.CI(un36_prod_a_b_cry_0),.S(un36_prod_a_b_axb_1),.LO(un36_prod_a_b_cry_1));
  MUXCY_L un36_prod_a_b_cry_0_cZ(.DI(un36_prod_a_b_cry_0_RNO),.CI(GND),.S(mul_24_fract_48[13:13]),.LO(un36_prod_a_b_cry_0));
  DSP48E1 desc1020(.ACOUT(ACOUT[29:0]),.BCOUT(BCOUT[17:0]),.CARRYCASCOUT(CARRYCASCOUT),.CARRYOUT(CARRYOUT[3:0]),.MULTSIGNOUT(MULTSIGNOUT),.OVERFLOW(OVERFLOW),.P({P_uc[47:12],un139_prod2[11:0]}),.PATTERNBDETECT(PATTERNBDETECT),.PATTERNDETECT(PATTERNDETECT),.PCOUT(PCOUT[47:0]),.UNDERFLOW(UNDERFLOW),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,opa_i[17:12]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,N_124_0_i,un8_prod2[34:30]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(s_state),.CEM(GND),.CEP(GND),.CLK(clk_i),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,s_opa_i_5,s_opa_i_4,s_opa_i_3,s_opa_i_2,s_opa_i_1,s_opa_i_0}),.INMODE({GND,GND,N_2719,N_2719,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(s_start_i),.RSTM(GND),.RSTP(GND));
defparam desc1020.ACASCREG=2;
defparam desc1020.ADREG=0;
defparam desc1020.ALUMODEREG=0;
defparam desc1020.AREG=2;
defparam desc1020.AUTORESET_PATDET="NO_RESET";
defparam desc1020.A_INPUT="DIRECT";
defparam desc1020.BCASCREG=0;
defparam desc1020.BREG=0;
defparam desc1020.B_INPUT="DIRECT";
defparam desc1020.CARRYINREG=0;
defparam desc1020.CARRYINSELREG=0;
defparam desc1020.CREG=1;
defparam desc1020.DREG=1;
defparam desc1020.INMODEREG=1;
defparam desc1020.MREG=0;
defparam desc1020.OPMODEREG=0;
defparam desc1020.PREG=0;
defparam desc1020.USE_DPORT="TRUE";
defparam desc1020.USE_MULT="MULTIPLY";
defparam desc1020.USE_SIMD="ONE48";
  DSP48E1 desc1021(.ACOUT(ACOUT_0[29:0]),.BCOUT(BCOUT_0[17:0]),.CARRYCASCOUT(CARRYCASCOUT_0),.CARRYOUT(CARRYOUT_0[3:0]),.MULTSIGNOUT(MULTSIGNOUT_0),.OVERFLOW(OVERFLOW_0),.P({P_uc_0[47:12],un184_prod2[11:0]}),.PATTERNBDETECT(PATTERNBDETECT_0),.PATTERNDETECT(PATTERNDETECT_0),.PCOUT(PCOUT_0[47:0]),.UNDERFLOW(UNDERFLOW_0),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,opb_i[17:12]}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,N_1411,N_1410,N_1409,N_248,N_1408,N_246}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(VCC),.CEM(GND),.CEP(GND),.CLK(clk_i),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,s_opb_i_5,s_opb_i_4,s_opb_i_3,s_opb_i_2,s_opb_i_1,s_opb_i_0}),.INMODE({GND,GND,N_235_mux,N_235_mux,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(s_start_i),.RSTM(GND),.RSTP(GND));
defparam desc1021.ACASCREG=2;
defparam desc1021.ADREG=0;
defparam desc1021.ALUMODEREG=0;
defparam desc1021.AREG=2;
defparam desc1021.AUTORESET_PATDET="NO_RESET";
defparam desc1021.A_INPUT="DIRECT";
defparam desc1021.BCASCREG=0;
defparam desc1021.BREG=0;
defparam desc1021.B_INPUT="DIRECT";
defparam desc1021.CARRYINREG=0;
defparam desc1021.CARRYINSELREG=0;
defparam desc1021.CREG=1;
defparam desc1021.DREG=1;
defparam desc1021.INMODEREG=1;
defparam desc1021.MREG=0;
defparam desc1021.OPMODEREG=0;
defparam desc1021.PREG=0;
defparam desc1021.USE_DPORT="TRUE";
defparam desc1021.USE_MULT="MULTIPLY";
defparam desc1021.USE_SIMD="ONE48";
  DSP48E1 desc1022(.ACOUT(ACOUT_1[29:0]),.BCOUT(BCOUT_1[17:0]),.CARRYCASCOUT(CARRYCASCOUT_1),.CARRYOUT(CARRYOUT_1[3:0]),.MULTSIGNOUT(MULTSIGNOUT_1),.OVERFLOW(OVERFLOW_1),.P({P_uc_1[47:12],un23_prod2[11:0]}),.PATTERNBDETECT(PATTERNBDETECT_1),.PATTERNDETECT(PATTERNDETECT_1),.PCOUT(PCOUT_1[47:0]),.UNDERFLOW(UNDERFLOW_1),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,result_i_o3_lut6_2_O6,s_opa_i_22,s_opa_i_21,s_opa_i_20,s_opa_i_19,s_opa_i_18}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,N_124_0_i,un8_prod2[34:30]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(s_state),.CEM(GND),.CEP(GND),.CLK(clk_i),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,s_opa_i_11,s_opa_i_10,s_opa_i_9,s_opa_i_8,s_opa_i_7,s_opa_i_6}),.INMODE({GND,GND,N_2719,N_2719,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(s_start_i),.RSTM(GND),.RSTP(GND));
defparam desc1022.ACASCREG=1;
defparam desc1022.ADREG=0;
defparam desc1022.ALUMODEREG=0;
defparam desc1022.AREG=1;
defparam desc1022.AUTORESET_PATDET="NO_RESET";
defparam desc1022.A_INPUT="DIRECT";
defparam desc1022.BCASCREG=0;
defparam desc1022.BREG=0;
defparam desc1022.B_INPUT="DIRECT";
defparam desc1022.CARRYINREG=0;
defparam desc1022.CARRYINSELREG=0;
defparam desc1022.CREG=1;
defparam desc1022.DREG=1;
defparam desc1022.INMODEREG=1;
defparam desc1022.MREG=0;
defparam desc1022.OPMODEREG=0;
defparam desc1022.PREG=0;
defparam desc1022.USE_DPORT="TRUE";
defparam desc1022.USE_MULT="MULTIPLY";
defparam desc1022.USE_SIMD="ONE48";
  DSP48E1 desc1023(.ACOUT(ACOUT_2[29:0]),.BCOUT(BCOUT_2[17:0]),.CARRYCASCOUT(CARRYCASCOUT_2),.CARRYOUT(CARRYOUT_2[3:0]),.MULTSIGNOUT(MULTSIGNOUT_2),.OVERFLOW(OVERFLOW_2),.P({P_uc_2[47:12],un92_prod2[11:0]}),.PATTERNBDETECT(PATTERNBDETECT_2),.PATTERNDETECT(PATTERNDETECT_2),.PCOUT(PCOUT_2[47:0]),.UNDERFLOW(UNDERFLOW_2),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,result_i_o3_lut6_2_O6,s_opa_i_22,s_opa_i_21,s_opa_i_20,s_opa_i_19,s_opa_i_18}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,un8_prod2[47:42]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(GND),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(VCC),.CEINMODE(s_state),.CEM(GND),.CEP(GND),.CLK(clk_i),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,s_opa_i_11,s_opa_i_10,s_opa_i_9,s_opa_i_8,s_opa_i_7,s_opa_i_6}),.INMODE({GND,GND,N_2719,N_2719,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(s_start_i),.RSTM(GND),.RSTP(GND));
defparam desc1023.ACASCREG=1;
defparam desc1023.ADREG=0;
defparam desc1023.ALUMODEREG=0;
defparam desc1023.AREG=1;
defparam desc1023.AUTORESET_PATDET="NO_RESET";
defparam desc1023.A_INPUT="DIRECT";
defparam desc1023.BCASCREG=0;
defparam desc1023.BREG=0;
defparam desc1023.B_INPUT="DIRECT";
defparam desc1023.CARRYINREG=0;
defparam desc1023.CARRYINSELREG=0;
defparam desc1023.CREG=1;
defparam desc1023.DREG=1;
defparam desc1023.INMODEREG=1;
defparam desc1023.MREG=0;
defparam desc1023.OPMODEREG=0;
defparam desc1023.PREG=0;
defparam desc1023.USE_DPORT="TRUE";
defparam desc1023.USE_MULT="MULTIPLY";
defparam desc1023.USE_SIMD="ONE48";
  FDRE desc1024(.Q(count[1:1]),.D(N_2719),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDR desc1025(.Q(count[0:0]),.D(N_235_mux),.C(clk_i),.R(s_start_i));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT3 desc1026(.I0(s_fracta_i[2:2]),.I1(s_fracta_i[14:14]),.I2(count[1:1]),.O(N_248));
defparam desc1026.INIT=8'hAC;
  LUT3 desc1027(.I0(s_fracta_i[1:1]),.I1(s_fracta_i[13:13]),.I2(count[1:1]),.O(N_1408));
defparam desc1027.INIT=8'hAC;
  LUT3 desc1028(.I0(s_fracta_i[5:5]),.I1(s_fracta_i[17:17]),.I2(count[1:1]),.O(N_1411));
defparam desc1028.INIT=8'hAC;
  LUT3 desc1029(.I0(s_fracta_i[4:4]),.I1(s_fracta_i[16:16]),.I2(count[1:1]),.O(N_1410));
defparam desc1029.INIT=8'hAC;
  LUT3 desc1030(.I0(s_fractb_i_1),.I1(s_fractb_i_13),.I2(count[0:0]),.O(un8_prod2[43:43]));
defparam desc1030.INIT=8'hAC;
  LUT3 desc1031(.I0(s_fractb_i_0),.I1(s_fractb_i_12),.I2(count[0:0]),.O(un8_prod2[42:42]));
defparam desc1031.INIT=8'hAC;
  LUT3 desc1032(.I0(s_fractb_i_3),.I1(s_fractb_i_15),.I2(count[0:0]),.O(un8_prod2[45:45]));
defparam desc1032.INIT=8'hAC;
  LUT3 desc1033(.I0(s_fractb_i_2),.I1(s_fractb_i_14),.I2(count[0:0]),.O(un8_prod2[44:44]));
defparam desc1033.INIT=8'hAC;
  LUT3 desc1034(.I0(s_fractb_i_5),.I1(s_fractb_i_17),.I2(count[0:0]),.O(un8_prod2[47:47]));
defparam desc1034.INIT=8'hAC;
  LUT3 desc1035(.I0(s_fractb_i_4),.I1(s_fractb_i_16),.I2(count[0:0]),.O(un8_prod2[46:46]));
defparam desc1035.INIT=8'hAC;
  LUT3 desc1036(.I0(s_fractb_i_7),.I1(s_fractb_i_19),.I2(count[0:0]),.O(un8_prod2[31:31]));
defparam desc1036.INIT=8'hAC;
  LUT3 desc1037(.I0(s_fractb_i_6),.I1(s_fractb_i_18),.I2(count[0:0]),.O(un8_prod2[30:30]));
defparam desc1037.INIT=8'hAC;
  LUT3 desc1038(.I0(s_fractb_i_10),.I1(s_fractb_i_22),.I2(count[0:0]),.O(un8_prod2[34:34]));
defparam desc1038.INIT=8'hAC;
  LUT3 desc1039(.I0(s_fractb_i_9),.I1(s_fractb_i_21),.I2(count[0:0]),.O(un8_prod2[33:33]));
defparam desc1039.INIT=8'hAC;
  LUT3 desc1040(.I0(s_fracta_i[3:3]),.I1(s_fracta_i[15:15]),.I2(count[1:1]),.O(N_1409));
defparam desc1040.INIT=8'hAC;
  LUT3 desc1041(.I0(count[2:2]),.I1(count[1:1]),.I2(count[0:0]),.O(prod2_2_0_1_sqmuxa));
defparam desc1041.INIT=8'h04;
  LUT3 desc1042(.I0(count[2:2]),.I1(count[1:1]),.I2(count[0:0]),.O(prod2_1_0_1_sqmuxa));
defparam desc1042.INIT=8'h10;
  LUT3 desc1043(.I0(s_state),.I1(count[2:2]),.I2(count[1:1]),.O(N_2731_i_0_0));
defparam desc1043.INIT=8'hA2;
  LUT3 desc1044(.I0(s_state),.I1(count[2:2]),.I2(count[1:1]),.O(count_RNILIBD_1_O6[2:2]));
defparam desc1044.INIT=8'h08;
  LUT4 desc1045(.I0(s_state),.I1(count[2:2]),.I2(count[1:1]),.I3(count[0:0]),.O(m39));
defparam desc1045.INIT=16'h64C4;
  LUT3 desc1046(.I0(count[2:2]),.I1(count[1:1]),.I2(count[0:0]),.O(prod2_3_0_1_sqmuxa));
defparam desc1046.INIT=8'h40;
  LUT3 desc1047(.I0(s_state),.I1(count[1:1]),.I2(count[0:0]),.O(count_RNILIBD_0_O5[2:2]));
defparam desc1047.INIT=8'h08;
  LUT3 desc1048(.I0(s_fractb_i[23:23]),.I1(s_fractb_i_11),.I2(count[0:0]),.O(N_124_0_i));
defparam desc1048.INIT=8'hCA;
  LUT3 desc1049(.I0(s_fractb_i_8),.I1(s_fractb_i_20),.I2(count[0:0]),.O(un8_prod2[32:32]));
defparam desc1049.INIT=8'hAC;
  LUT3 desc1050(.I0(count[2:2]),.I1(count[1:1]),.I2(count[0:0]),.O(N_2719));
defparam desc1050.INIT=8'h1C;
  LUT3 desc1051(.I0(s_state),.I1(count[1:1]),.I2(count[0:0]),.O(count_RNILIBD_2_O5[2:2]));
defparam desc1051.INIT=8'h20;
  LUT4 desc1052(.I0(s_state),.I1(count[2:2]),.I2(count[1:1]),.I3(count[0:0]),.O(N_235_mux));
defparam desc1052.INIT=16'h55A2;
  LUT3 desc1053(.I0(s_state),.I1(count[1:1]),.I2(count[0:0]),.O(count_RNILIBD_O5[2:2]));
defparam desc1053.INIT=8'h80;
  LUT3 desc1054(.I0(s_fracta_i[0:0]),.I1(s_fracta_i[12:12]),.I2(count[1:1]),.O(N_246));
defparam desc1054.INIT=8'hAC;
  LUT3 desc1055(.I0(count[2:2]),.I1(count[1:1]),.I2(count[0:0]),.O(un2_i));
defparam desc1055.INIT=8'h01;
endmodule
module post_norm_mul_inj (pre_norm_mul_exp_10,mul_24_fract_48,s_fracta_i_20,s_fracta_i_21,s_fracta_i_0,s_fracta_i_1,s_fracta_i_2,s_fracta_i_3,s_fracta_i_4,s_fracta_i_5,s_fracta_i_6,s_fracta_i_7,s_fracta_i_8,s_fracta_i_9,s_fracta_i_10,s_fracta_i_11,s_fracta_i_12,s_fracta_i_13,s_fracta_i_14,s_fracta_i_15,s_rmode_i,post_norm_mul_output,clk_i,N_6_i,post_norm_mul_ine,s_infb,un1_s_infa,result_5,un1_s_nan_b,result_4,un1_s_nan_a,un3_s_op_0,result_11,result_3_21_1,result_3_21_3,p_desc1070_p_O_FD,p_desc1071_p_O_FD,p_desc1072_p_O_FD,p_desc1073_p_O_FD,p_desc1074_p_O_FD,p_desc1075_p_O_FD,p_desc1076_p_O_FD,p_desc1077_p_O_FD,p_desc1078_p_O_FD,p_desc1079_p_O_FD,p_desc1080_p_O_FD,p_desc1081_p_O_FD,p_desc1082_p_O_FD,p_desc1083_p_O_FD,p_desc1084_p_O_FD,p_desc1085_p_O_FD,p_desc1086_p_O_FD,p_desc1087_p_O_FD,p_desc1088_p_O_FD,p_desc1089_p_O_FD,p_desc1090_p_O_FD,p_desc1091_p_O_FD,p_desc1092_p_O_FD,p_desc1163_p_O_FD,p_desc1164_p_O_FD,p_desc1165_p_O_FD,p_desc1166_p_O_FD,p_desc1167_p_O_FD,p_desc1168_p_O_FD,p_desc1169_p_O_FD,p_desc1170_p_O_FD,p_desc1171_p_O_FD,p_desc1172_p_O_FD,p_desc1173_p_O_FD,p_desc1174_p_O_FD,p_desc1175_p_O_FD,p_desc1176_p_O_FD,p_desc1177_p_O_FD,p_desc1178_p_O_FD,p_desc1179_p_O_FD,p_desc1180_p_O_FD,p_desc1181_p_O_FD,p_desc1182_p_O_FD,p_desc1183_p_O_FD,p_desc1184_p_O_FD,p_desc1185_p_O_FD,p_desc1186_p_O_FD,p_desc1187_p_O_FD,p_desc1188_p_O_FD,p_desc1189_p_O_FD,p_desc1190_p_O_FD,p_desc1191_p_O_FD,p_desc1192_p_O_FD,p_desc1193_p_O_FD,p_desc1194_p_O_FD,p_desc1195_p_O_FD,p_desc1196_p_O_FD,p_desc1197_p_O_FD,p_desc1198_p_O_FD,p_desc1199_p_O_FD,p_desc1200_p_O_FD,p_desc1201_p_O_FD,p_desc1202_p_O_FD,p_desc1203_p_O_FD,p_desc1204_p_O_FD,p_desc1205_p_O_FD,p_desc1206_p_O_FD,p_desc1207_p_O_FD,p_desc1208_p_O_FD,p_desc1209_p_O_FD,p_desc1210_p_O_FD,p_desc1211_p_O_FD,p_desc1212_p_O_FD,p_desc1213_p_O_FD,p_desc1214_p_O_FD,p_desc1215_p_O_FD,p_desc1216_p_O_FD,p_desc1217_p_O_FD,p_desc1218_p_O_FD,p_desc1219_p_O_FD,p_desc1220_p_O_FD,p_desc1221_p_O_FD,p_s_sign_i_Z_p_O_FD,p_ine_o_Z_p_O_FD,p_desc1244_p_O_FD,p_desc1245_p_O_FD,p_desc1246_p_O_FD,p_desc1247_p_O_FD,p_desc1248_p_O_FD,p_desc1249_p_O_FD,p_desc1250_p_O_FD,p_desc1251_p_O_FD,p_desc1252_p_O_FD,p_desc1253_p_O_FD,p_desc1254_p_O_FD,p_desc1255_p_O_FD,p_desc1256_p_O_FD,p_desc1257_p_O_FD,p_desc1258_p_O_FD,p_desc1259_p_O_FD,p_desc1260_p_O_FD,p_desc1261_p_O_FD,p_desc1262_p_O_FD,p_desc1263_p_O_FD,p_desc1264_p_O_FD,p_desc1265_p_O_FD,p_desc1266_p_O_FD,p_desc1267_p_O_FD,p_desc1268_p_O_FD,p_desc1269_p_O_FD,p_desc1270_p_O_FD,p_desc1271_p_O_FD,p_desc1272_p_O_FD,p_desc1273_p_O_FD,p_desc1274_p_O_FD,p_desc1275_p_O_FD,p_desc1276_p_O_FD,p_desc1277_p_O_FD,p_desc1278_p_O_FD,p_desc1279_p_O_FD,p_desc1280_p_O_FD,p_desc1281_p_O_FD,p_desc1282_p_O_FD,p_desc1283_p_O_FD,p_desc1284_p_O_FD,p_desc1285_p_O_FD,p_desc1286_p_O_FD,p_desc1287_p_O_FD,p_desc1288_p_O_FD,p_desc1289_p_O_FD,p_desc1290_p_O_FD,p_desc1291_p_O_FD);
input [9:0] pre_norm_mul_exp_10 ;
input [47:0] mul_24_fract_48 ;
input s_fracta_i_20 ;
input s_fracta_i_21 ;
input s_fracta_i_0 ;
input s_fracta_i_1 ;
input s_fracta_i_2 ;
input s_fracta_i_3 ;
input s_fracta_i_4 ;
input s_fracta_i_5 ;
input s_fracta_i_6 ;
input s_fracta_i_7 ;
input s_fracta_i_8 ;
input s_fracta_i_9 ;
input s_fracta_i_10 ;
input s_fracta_i_11 ;
input s_fracta_i_12 ;
input s_fracta_i_13 ;
input s_fracta_i_14 ;
input s_fracta_i_15 ;
input [1:0] s_rmode_i ;
output [31:0] post_norm_mul_output ;
input clk_i ;
input N_6_i ;
output post_norm_mul_ine ;
input s_infb ;
input un1_s_infa ;
input result_5 ;
input un1_s_nan_b ;
input result_4 ;
input un1_s_nan_a ;
input un3_s_op_0 ;
output result_11 ;
output result_3_21_1 ;
output result_3_21_3 ;
wire s_fracta_i_20 ;
wire s_fracta_i_21 ;
wire s_fracta_i_0 ;
wire s_fracta_i_1 ;
wire s_fracta_i_2 ;
wire s_fracta_i_3 ;
wire s_fracta_i_4 ;
wire s_fracta_i_5 ;
wire s_fracta_i_6 ;
wire s_fracta_i_7 ;
wire s_fracta_i_8 ;
wire s_fracta_i_9 ;
wire s_fracta_i_10 ;
wire s_fracta_i_11 ;
wire s_fracta_i_12 ;
wire s_fracta_i_13 ;
wire s_fracta_i_14 ;
wire s_fracta_i_15 ;
wire clk_i ;
wire N_6_i ;
wire post_norm_mul_ine ;
wire s_infb ;
wire un1_s_infa ;
wire result_5 ;
wire un1_s_nan_b ;
wire result_4 ;
wire un1_s_nan_a ;
wire un3_s_op_0 ;
wire result_11 ;
wire result_3_21_1 ;
wire result_3_21_3 ;
wire [5:0] s_zeros ;
wire [9:0] s_exp_10_i ;
wire [47:0] s_fract_48_i ;
wire s_exp_10b_i ;
wire s_zeros_RNI0TNS_O5 ;
wire [47:0] s_frac2a ;
wire [24:0] s_frac_rnd_3 ;
wire [5:0] s_shr2 ;
wire [15:0] s_frac2a_3 ;
wire [6:6] v_shr1_4 ;
wire [5:1] v_shr1_4_e ;
wire [9:1] s_exp_10b ;
wire [7:1] s_expo1_5 ;
wire [5:0] s_shl2 ;
wire [24:0] s_frac_rnd ;
wire s_zeros_2_0_i_a2_3_lut6_2_O5 ;
wire [46:46] s_fract_48_i_RNI21942_O6 ;
wire [3:3] s_fract_48_i_RNIEUJ9_O5 ;
wire [3:3] v_count_49_i_o3_i_a2_lut6_2_O5 ;
wire [1:1] v_count_49_i_a2_0_lut6_2_O6 ;
wire [3:3] v_count_49_i_o3_i_a2_lut6_2_O6 ;
wire [2:2] v_count_49_i_o2_1_i_a2_lut6_2_O6 ;
wire [2:2] v_count_49_i_o2_0_i_a2_lut6_2_O6 ;
wire s_zeros_2_0_i_a2_1_2_lut6_2_O5 ;
wire [1:1] v_count_49_i_0 ;
wire [5:0] s_r_zeros ;
wire [21:0] s_output_o_0 ;
wire [7:0] s_expo1 ;
wire s_expo1_5_e ;
wire s_shr2_0_e ;
wire [2:2] s_exp_10_i_RNIE6AQ1 ;
wire [2:2] s_exp_10_i_RNI5I152 ;
wire [2:2] s_zeros_2_2 ;
wire [3:2] s_zeros_2_0 ;
wire [22:22] s_output_o ;
wire [30:23] s_output_o_m0 ;
wire [7:0] s_expo2b ;
wire [7:7] s_expo3 ;
wire [4:4] v_count_49_0_o2 ;
wire [1:1] v_count_49_i_o3_1 ;
wire [4:4] v_count_49_0_o2_9 ;
wire [4:4] v_count_49_0_o2_6 ;
wire [2:2] s_exp_10_i_RNIORIF1 ;
wire v_count_49_1_3 ;
wire [4:0] v_count_49 ;
wire [3:3] v_count_49_i_i ;
wire v_count_49_0_4 ;
wire v_count_49_0 ;
wire [2:2] s_r_zeros_RNO_0 ;
wire v_count_49_1_1 ;
wire N_1247_i ;
wire N_1247 ;
wire N_903_i ;
wire N_903 ;
wire N_16_0_i ;
wire N_16_0 ;
wire GND ;
wire VCC ;
wire s_frac_rnd_3_0_s_1 ;
wire s_roundup ;
wire s_frac_rnd_3_0_s_2 ;
wire s_frac_rnd_3_0_s_3 ;
wire s_frac_rnd_3_0_s_4 ;
wire s_frac_rnd_3_0_s_5 ;
wire s_frac_rnd_3_0_s_6 ;
wire s_frac_rnd_3_0_s_7 ;
wire s_frac_rnd_3_0_s_8 ;
wire s_frac_rnd_3_0_s_9 ;
wire s_frac_rnd_3_0_s_10 ;
wire s_frac_rnd_3_0_s_11 ;
wire s_frac_rnd_3_0_s_12 ;
wire s_frac_rnd_3_0_s_13 ;
wire s_frac_rnd_3_0_s_14 ;
wire s_frac_rnd_3_0_s_15 ;
wire s_frac_rnd_3_0_s_17 ;
wire s_frac_rnd_3_0_s_18 ;
wire s_frac_rnd_3_0_s_19 ;
wire s_frac_rnd_3_0_s_20 ;
wire s_frac_rnd_3_0_s_21 ;
wire s_frac_rnd_3_0_s_22 ;
wire s_frac_rnd_3_0_s_23 ;
wire s_frac_rnd_3_0_s_24 ;
wire N_82_0 ;
wire N_80_0 ;
wire N_79_0 ;
wire N_459_i ;
wire un6_s_exp_10a ;
wire un1_s_exp_10a_3_1 ;
wire un1_s_exp_10a_3_lut6_2_O6 ;
wire s_exp_10b_s_1_RNI0PGD1_O6 ;
wire N_368 ;
wire N_1078 ;
wire m368_lut6_2_O6 ;
wire N_1081 ;
wire N_1120 ;
wire N_240 ;
wire N_242 ;
wire N_1114 ;
wire N_1121 ;
wire N_243 ;
wire N_67 ;
wire N_71 ;
wire N_111 ;
wire N_1103 ;
wire N_1102 ;
wire N_69 ;
wire N_65 ;
wire N_109 ;
wire N_219 ;
wire N_218 ;
wire N_126 ;
wire N_134 ;
wire s_frac2a_1_132 ;
wire s_frac2a_1_124 ;
wire s_frac2a_1_124_RNIEJB51_O6 ;
wire N_355 ;
wire N_85 ;
wire N_905 ;
wire N_904 ;
wire N_223 ;
wire N_1165 ;
wire un1_s_shr2_1_4 ;
wire N_138 ;
wire N_1156 ;
wire N_337 ;
wire N_396 ;
wire N_72 ;
wire N_80 ;
wire N_76 ;
wire N_25_0 ;
wire N_297 ;
wire N_68 ;
wire N_52 ;
wire N_1084 ;
wire N_265 ;
wire N_64 ;
wire N_60 ;
wire N_1085 ;
wire N_289 ;
wire N_56 ;
wire N_1086 ;
wire N_280 ;
wire N_62 ;
wire N_66 ;
wire N_58 ;
wire N_1094 ;
wire N_360 ;
wire N_50 ;
wire N_54 ;
wire N_1096 ;
wire N_361 ;
wire N_78 ;
wire N_74 ;
wire N_70 ;
wire N_1140 ;
wire N_370 ;
wire N_139 ;
wire N_228 ;
wire N_245 ;
wire N_196 ;
wire N_371 ;
wire N_1158 ;
wire N_1160 ;
wire N_357 ;
wire N_51 ;
wire N_55 ;
wire N_214 ;
wire N_99 ;
wire N_71_0 ;
wire N_67_0 ;
wire N_79 ;
wire N_75 ;
wire N_977 ;
wire N_115_i ;
wire N_73 ;
wire N_106 ;
wire N_121 ;
wire N_81 ;
wire N_77 ;
wire N_110 ;
wire N_129 ;
wire N_63 ;
wire N_59 ;
wire s_frac2a_2_115_lut6_2_O6 ;
wire N_61 ;
wire N_57 ;
wire N_115 ;
wire N_85_0 ;
wire N_86 ;
wire s_frac2a_2_91 ;
wire N_49 ;
wire N_137 ;
wire N_1157 ;
wire un2_s_lost_c4 ;
wire un2_s_lost_ac0_5_lut6_2_O5 ;
wire N_55_0 ;
wire un2_s_exp_10a_c3 ;
wire un5_v_shr1_c3 ;
wire un2_s_exp_10a_c2 ;
wire v_shl1_5_0_0_c2 ;
wire N_654 ;
wire N_1255 ;
wire N_1317 ;
wire N_35_0 ;
wire v_count_0_sqmuxa_47_4_4 ;
wire m107_i_a2_7_0 ;
wire v_count_0_sqmuxa_47_1_4 ;
wire N_425 ;
wire N_641_1 ;
wire N_314_1 ;
wire N_320_0_3 ;
wire N_173 ;
wire N_40 ;
wire N_20_0 ;
wire N_88 ;
wire N_92 ;
wire N_269 ;
wire N_1254 ;
wire N_1076 ;
wire N_1124 ;
wire N_1289 ;
wire N_1077 ;
wire N_1288 ;
wire N_36 ;
wire N_1252 ;
wire N_3 ;
wire N_653 ;
wire N_326_2 ;
wire v_count_0_sqmuxa_47_2_4 ;
wire N_624 ;
wire N_588 ;
wire N_668_3 ;
wire N_614 ;
wire v_count_0_sqmuxa_47_3_3 ;
wire N_592 ;
wire N_1353 ;
wire N_707 ;
wire N_1361 ;
wire N_447 ;
wire N_449 ;
wire N_1264 ;
wire N_426 ;
wire N_1350 ;
wire N_582 ;
wire N_597 ;
wire N_672 ;
wire N_673 ;
wire N_677 ;
wire N_37 ;
wire N_446 ;
wire N_1251 ;
wire N_434_i_0 ;
wire N_610 ;
wire N_1371 ;
wire N_1367 ;
wire N_1260 ;
wire N_591 ;
wire N_1249 ;
wire N_1245 ;
wire N_464_1 ;
wire N_1246 ;
wire N_638 ;
wire N_326_1 ;
wire N_1253 ;
wire N_704 ;
wire N_687 ;
wire N_1259 ;
wire N_689 ;
wire N_239 ;
wire N_301 ;
wire N_663_3 ;
wire N_708 ;
wire N_320_2 ;
wire N_1308 ;
wire un1_s_expo3 ;
wire s_output_o25_sn ;
wire N_530_1 ;
wire N_505_1_2 ;
wire v_count_0_sqmuxa_47_3_4 ;
wire N_331_1 ;
wire N_481 ;
wire N_1261 ;
wire N_326_0_3 ;
wire N_599 ;
wire N_543 ;
wire m80_0_e ;
wire m97_0_e ;
wire m37_0_0_e ;
wire m102_0_e ;
wire m108_0_0_e ;
wire m113_0_e ;
wire m119_0_0_e ;
wire m169_0_e ;
wire m224_0_e ;
wire m231_0_e ;
wire m237_0_e ;
wire m293_0_e ;
wire m365_0_e ;
wire m374_0_e ;
wire m378_0_e ;
wire m435_0_e ;
wire N_1168 ;
wire N_169 ;
wire N_284 ;
wire N_286 ;
wire N_376 ;
wire N_372 ;
wire N_333 ;
wire N_363 ;
wire N_271 ;
wire N_275 ;
wire N_291 ;
wire N_211 ;
wire N_235 ;
wire N_194 ;
wire N_229 ;
wire N_217 ;
wire N_221 ;
wire N_1137 ;
wire N_1142 ;
wire N_1112 ;
wire N_69_0 ;
wire N_71_0_0 ;
wire N_1109 ;
wire N_52_0 ;
wire N_56_0 ;
wire N_1104 ;
wire N_60_0 ;
wire N_64_0 ;
wire N_1098 ;
wire N_1083 ;
wire N_1087 ;
wire N_1090 ;
wire s_frac2a_1_141_RNIA10R ;
wire N_78_0 ;
wire N_382 ;
wire N_161 ;
wire un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91 ;
wire N_503_1 ;
wire s_output_o_sm0 ;
wire N_247 ;
wire N_1277 ;
wire N_1372 ;
wire N_315 ;
wire N_414_i_0 ;
wire v_count_0_sqmuxa_47_0 ;
wire v_count_0_sqmuxa_47_1_0 ;
wire v_count_0_sqmuxa_47_1 ;
wire N_23_0_3 ;
wire N_23_0_4 ;
wire N_23_4 ;
wire N_23_i_0 ;
wire N_62_1 ;
wire N_62_i_0 ;
wire s_expo2b_axb_1 ;
wire s_expo2b_axb_2 ;
wire s_expo2b_axb_3 ;
wire s_expo2b_axb_4 ;
wire s_expo2b_axb_5 ;
wire s_expo2b_axb_6 ;
wire s_exp_10b_axb_1 ;
wire s_frac_rnd_3_0_axb_1 ;
wire s_frac_rnd_3_0_axb_2 ;
wire s_frac_rnd_3_0_axb_3 ;
wire s_frac_rnd_3_0_axb_4 ;
wire s_frac_rnd_3_0_axb_5 ;
wire s_frac_rnd_3_0_axb_6 ;
wire s_frac_rnd_3_0_axb_7 ;
wire s_frac_rnd_3_0_axb_8 ;
wire s_frac_rnd_3_0_axb_9 ;
wire s_frac_rnd_3_0_axb_10 ;
wire s_frac_rnd_3_0_axb_11 ;
wire s_frac_rnd_3_0_axb_12 ;
wire s_frac_rnd_3_0_axb_13 ;
wire s_frac_rnd_3_0_axb_14 ;
wire s_frac_rnd_3_0_axb_15 ;
wire s_frac_rnd_3_0_axb_16 ;
wire s_frac_rnd_3_0_axb_17 ;
wire s_frac_rnd_3_0_axb_18 ;
wire s_frac_rnd_3_0_axb_19 ;
wire s_frac_rnd_3_0_axb_20 ;
wire s_frac_rnd_3_0_axb_21 ;
wire s_frac_rnd_3_0_axb_22 ;
wire s_frac_rnd_3_0_axb_23 ;
wire s_sign_i ;
wire un1_s_ine_o ;
wire N_715 ;
wire N_716 ;
wire N_717 ;
wire N_718 ;
wire N_719 ;
wire N_406 ;
wire N_411 ;
wire N_1117 ;
wire N_1148 ;
wire N_441 ;
wire N_308 ;
wire N_256 ;
wire N_184 ;
wire N_1123 ;
wire N_1131 ;
wire N_389 ;
wire N_401 ;
wire N_300 ;
wire N_714 ;
wire N_709 ;
wire N_331_0_4 ;
wire N_1328 ;
wire N_535 ;
wire N_693 ;
wire N_700_1 ;
wire N_320_0 ;
wire un7_s_expo3_c4 ;
wire N_307 ;
wire N_299 ;
wire N_1147 ;
wire N_410 ;
wire N_679 ;
wire N_1364 ;
wire N_611 ;
wire N_637 ;
wire un1_s_overflow_2 ;
wire N_1358 ;
wire N_1365 ;
wire N_1370 ;
wire N_1267 ;
wire N_626 ;
wire N_253 ;
wire N_404 ;
wire N_234 ;
wire N_260 ;
wire N_84 ;
wire N_66_0 ;
wire N_74_0 ;
wire N_72_0 ;
wire N_1141 ;
wire s_exp_10b_axb_3 ;
wire N_80_1 ;
wire N_76_0 ;
wire N_70_0 ;
wire N_64_1 ;
wire N_68_0 ;
wire m40 ;
wire N_47 ;
wire N_304 ;
wire N_327 ;
wire N_31_0 ;
wire N_87 ;
wire N_83 ;
wire N_103 ;
wire N_77_0 ;
wire N_131 ;
wire N_1337 ;
wire N_60_1 ;
wire N_62_0 ;
wire N_322 ;
wire N_101 ;
wire N_206 ;
wire N_1273 ;
wire N_192 ;
wire s_output_o_sn_N_5_mux ;
wire un1_s_overflow_0 ;
wire N_1129 ;
wire N_354 ;
wire N_12_0 ;
wire s_frac2a_1_134 ;
wire un3_s_ine_o ;
wire N_443 ;
wire s_frac_rnd_3_0_axb_24 ;
wire s_expo2b_axb_7 ;
wire N_30 ;
wire N_273 ;
wire N_279 ;
wire un4_s_exp_10b_0_2 ;
wire un3_s_ine_o_0_0 ;
wire un3_s_ine_o_0_1 ;
wire un3_s_ine_o_0_2 ;
wire result_3_21_0 ;
wire N_49_0 ;
wire N_53 ;
wire N_55_1 ;
wire N_53_0 ;
wire s_frac2a_1_58 ;
wire N_58_0 ;
wire N_59_0 ;
wire s_frac2a_1_62 ;
wire N_63_0 ;
wire N_65_0 ;
wire N_69_1 ;
wire N_75_0 ;
wire N_84_0 ;
wire N_60_0_0 ;
wire N_81_0 ;
wire N_82 ;
wire N_79_1 ;
wire N_87_0 ;
wire N_83_0 ;
wire N_77_1 ;
wire N_73_0 ;
wire un5_v_shr1_axb1 ;
wire un5_s_exp_10a_1 ;
wire un2_s_lost_axbxc3 ;
wire un2_s_exp_10a_c4 ;
wire N_1305 ;
wire N_318 ;
wire N_250 ;
wire N_1150 ;
wire N_1125 ;
wire s_frac2a_2_111 ;
wire N_105 ;
wire s_frac2a_1_109 ;
wire N_23_0_2 ;
wire un4_s_lost_c2 ;
wire N_686 ;
wire N_1093 ;
wire v_count_0_sqmuxa_46_0 ;
wire N_331_0 ;
wire N_669_0 ;
wire N_662 ;
wire N_650 ;
wire un3_s_ine_o_0 ;
wire N_263 ;
wire N_161_0 ;
wire N_153 ;
wire N_423 ;
wire N_1154 ;
wire N_349 ;
wire N_342 ;
wire N_325 ;
wire N_296 ;
wire N_278 ;
wire N_201 ;
wire N_1152 ;
wire N_1128 ;
wire N_85_0_0 ;
wire N_74_0_0 ;
wire N_64_0_0 ;
wire N_44_1 ;
wire N_938 ;
wire N_7_0 ;
wire N_158 ;
wire v_count_0_sqmuxa_46 ;
wire N_1281_2 ;
wire N_1167 ;
wire N_190 ;
wire N_116 ;
wire i40_mux ;
wire N_399 ;
wire N_254 ;
wire N_1153 ;
wire N_1115 ;
wire N_921 ;
wire N_195 ;
wire N_1340 ;
wire v_shl1_5_0_0_c4 ;
wire un2_s_exp_10a_c8 ;
wire N_688 ;
wire N_658 ;
wire N_330 ;
wire N_268 ;
wire i104_mux ;
wire un4_s_lost_c4 ;
wire N_344 ;
wire N_67_0_0 ;
wire N_49_0_0 ;
wire N_57_0 ;
wire N_1163 ;
wire N_283 ;
wire N_208 ;
wire N_1134 ;
wire N_87_0_0 ;
wire N_6484_i ;
wire N_622 ;
wire N_6485_i ;
wire N_6482_i ;
wire N_6483_i ;
wire N_326_2_0 ;
wire un4_s_lost_c6 ;
wire N_1271 ;
wire un16_s_roundup ;
wire N_663_2 ;
wire N_314 ;
wire N_641 ;
wire N_566_i ;
wire s_frac_rnd_3_0_s_16 ;
wire N_564_i ;
wire s_exp_10b_axb_2 ;
wire s_exp_10b_axb_4 ;
wire s_exp_10b_axb_5 ;
wire s_exp_10b_cry_6_RNO ;
wire s_exp_10b_cry_7_RNO ;
wire s_frac_rnd_3_0_cry_23 ;
wire s_frac_rnd_3_0_cry_22 ;
wire s_frac_rnd_3_0_cry_21 ;
wire s_frac_rnd_3_0_cry_20 ;
wire s_frac_rnd_3_0_cry_19 ;
wire s_frac_rnd_3_0_cry_18 ;
wire s_frac_rnd_3_0_cry_17 ;
wire s_frac_rnd_3_0_cry_16 ;
wire s_frac_rnd_3_0_cry_15 ;
wire s_frac_rnd_3_0_cry_14 ;
wire s_frac_rnd_3_0_cry_13 ;
wire s_frac_rnd_3_0_cry_12 ;
wire s_frac_rnd_3_0_cry_11 ;
wire s_frac_rnd_3_0_cry_10 ;
wire s_frac_rnd_3_0_cry_9 ;
wire s_frac_rnd_3_0_cry_8 ;
wire s_frac_rnd_3_0_cry_7 ;
wire s_frac_rnd_3_0_cry_6 ;
wire s_frac_rnd_3_0_cry_5 ;
wire s_frac_rnd_3_0_cry_4 ;
wire s_frac_rnd_3_0_cry_3 ;
wire s_frac_rnd_3_0_cry_2 ;
wire s_frac_rnd_3_0_cry_1 ;
wire s_exp_10b_cry_8 ;
wire s_exp_10b_cry_7 ;
wire s_exp_10b_cry_6 ;
wire s_exp_10b_cry_5 ;
wire s_exp_10b_cry_4 ;
wire s_exp_10b_cry_3 ;
wire s_exp_10b_cry_2 ;
wire s_exp_10b_cry_1 ;
wire s_exp_10b_cry_0 ;
wire s_expo2b_cry_6 ;
wire s_expo2b_cry_5 ;
wire s_expo2b_cry_4 ;
wire s_expo2b_cry_3 ;
wire s_expo2b_cry_2 ;
wire s_expo2b_cry_1 ;
wire s_expo2b_cry_0 ;
input p_desc1070_p_O_FD ;
input p_desc1071_p_O_FD ;
input p_desc1072_p_O_FD ;
input p_desc1073_p_O_FD ;
input p_desc1074_p_O_FD ;
input p_desc1075_p_O_FD ;
input p_desc1076_p_O_FD ;
input p_desc1077_p_O_FD ;
input p_desc1078_p_O_FD ;
input p_desc1079_p_O_FD ;
input p_desc1080_p_O_FD ;
input p_desc1081_p_O_FD ;
input p_desc1082_p_O_FD ;
input p_desc1083_p_O_FD ;
input p_desc1084_p_O_FD ;
input p_desc1085_p_O_FD ;
input p_desc1086_p_O_FD ;
input p_desc1087_p_O_FD ;
input p_desc1088_p_O_FD ;
input p_desc1089_p_O_FD ;
input p_desc1090_p_O_FD ;
input p_desc1091_p_O_FD ;
input p_desc1092_p_O_FD ;
input p_desc1163_p_O_FD ;
input p_desc1164_p_O_FD ;
input p_desc1165_p_O_FD ;
input p_desc1166_p_O_FD ;
input p_desc1167_p_O_FD ;
input p_desc1168_p_O_FD ;
input p_desc1169_p_O_FD ;
input p_desc1170_p_O_FD ;
input p_desc1171_p_O_FD ;
input p_desc1172_p_O_FD ;
input p_desc1173_p_O_FD ;
input p_desc1174_p_O_FD ;
input p_desc1175_p_O_FD ;
input p_desc1176_p_O_FD ;
input p_desc1177_p_O_FD ;
input p_desc1178_p_O_FD ;
input p_desc1179_p_O_FD ;
input p_desc1180_p_O_FD ;
input p_desc1181_p_O_FD ;
input p_desc1182_p_O_FD ;
input p_desc1183_p_O_FD ;
input p_desc1184_p_O_FD ;
input p_desc1185_p_O_FD ;
input p_desc1186_p_O_FD ;
input p_desc1187_p_O_FD ;
input p_desc1188_p_O_FD ;
input p_desc1189_p_O_FD ;
input p_desc1190_p_O_FD ;
input p_desc1191_p_O_FD ;
input p_desc1192_p_O_FD ;
input p_desc1193_p_O_FD ;
input p_desc1194_p_O_FD ;
input p_desc1195_p_O_FD ;
input p_desc1196_p_O_FD ;
input p_desc1197_p_O_FD ;
input p_desc1198_p_O_FD ;
input p_desc1199_p_O_FD ;
input p_desc1200_p_O_FD ;
input p_desc1201_p_O_FD ;
input p_desc1202_p_O_FD ;
input p_desc1203_p_O_FD ;
input p_desc1204_p_O_FD ;
input p_desc1205_p_O_FD ;
input p_desc1206_p_O_FD ;
input p_desc1207_p_O_FD ;
input p_desc1208_p_O_FD ;
input p_desc1209_p_O_FD ;
input p_desc1210_p_O_FD ;
input p_desc1211_p_O_FD ;
input p_desc1212_p_O_FD ;
input p_desc1213_p_O_FD ;
input p_desc1214_p_O_FD ;
input p_desc1215_p_O_FD ;
input p_desc1216_p_O_FD ;
input p_desc1217_p_O_FD ;
input p_desc1218_p_O_FD ;
input p_desc1219_p_O_FD ;
input p_desc1220_p_O_FD ;
input p_desc1221_p_O_FD ;
input p_s_sign_i_Z_p_O_FD ;
input p_ine_o_Z_p_O_FD ;
input p_desc1244_p_O_FD ;
input p_desc1245_p_O_FD ;
input p_desc1246_p_O_FD ;
input p_desc1247_p_O_FD ;
input p_desc1248_p_O_FD ;
input p_desc1249_p_O_FD ;
input p_desc1250_p_O_FD ;
input p_desc1251_p_O_FD ;
input p_desc1252_p_O_FD ;
input p_desc1253_p_O_FD ;
input p_desc1254_p_O_FD ;
input p_desc1255_p_O_FD ;
input p_desc1256_p_O_FD ;
input p_desc1257_p_O_FD ;
input p_desc1258_p_O_FD ;
input p_desc1259_p_O_FD ;
input p_desc1260_p_O_FD ;
input p_desc1261_p_O_FD ;
input p_desc1262_p_O_FD ;
input p_desc1263_p_O_FD ;
input p_desc1264_p_O_FD ;
input p_desc1265_p_O_FD ;
input p_desc1266_p_O_FD ;
input p_desc1267_p_O_FD ;
input p_desc1268_p_O_FD ;
input p_desc1269_p_O_FD ;
input p_desc1270_p_O_FD ;
input p_desc1271_p_O_FD ;
input p_desc1272_p_O_FD ;
input p_desc1273_p_O_FD ;
input p_desc1274_p_O_FD ;
input p_desc1275_p_O_FD ;
input p_desc1276_p_O_FD ;
input p_desc1277_p_O_FD ;
input p_desc1278_p_O_FD ;
input p_desc1279_p_O_FD ;
input p_desc1280_p_O_FD ;
input p_desc1281_p_O_FD ;
input p_desc1282_p_O_FD ;
input p_desc1283_p_O_FD ;
input p_desc1284_p_O_FD ;
input p_desc1285_p_O_FD ;
input p_desc1286_p_O_FD ;
input p_desc1287_p_O_FD ;
input p_desc1288_p_O_FD ;
input p_desc1289_p_O_FD ;
input p_desc1290_p_O_FD ;
input p_desc1291_p_O_FD ;
// instances
  INV desc1056(.I(N_1247_i),.O(N_1247));
  INV desc1057(.I(N_903_i),.O(N_903));
  INV desc1058(.I(N_16_0_i),.O(N_16_0));
  LUT6_2 desc1059(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_67),.I3(N_71),.I4(N_111),.I5(s_shl2[3:3]),.O6(N_1103),.O5(N_1102));
defparam desc1059.INIT=64'h3333000031203120;
  LUT6_2 desc1060(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_69),.I3(N_65),.I4(N_109),.I5(s_shl2[3:3]),.O6(N_219),.O5(N_218));
defparam desc1060.INIT=64'h3333000032103210;
  LUT6_2 desc1061(.I0(s_shl2[4:4]),.I1(s_shr2[3:3]),.I2(N_139),.I3(N_243),.I4(N_228),.I5(un1_s_shr2_1_4),.O6(N_245),.O5(N_196));
defparam desc1061.INIT=64'hFFAA550030303030;
  LUT6_2 desc1062(.I0(s_shl2[4:4]),.I1(s_shr2[3:3]),.I2(N_138),.I3(N_371),.I4(N_1158),.I5(un1_s_shr2_1_4),.O6(N_1160),.O5(N_357));
defparam desc1062.INIT=64'hAA00FF5530303030;
  LUT6_2 desc1063(.I0(s_shr2[2:2]),.I1(N_71_0),.I2(N_67_0),.I3(N_79),.I4(N_75),.I5(s_shr2[3:3]),.O6(N_977),.O5(N_115_i));
defparam desc1063.INIT=64'h00AA55FF27272727;
  LUT6_2 desc1064(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[47:47]),.I2(s_shr2[2:2]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.I5(s_shr2[3:3]),.O6(N_82_0),.O5(N_55_0));
defparam desc1064.INIT=64'h00000000000C000A;
  LUT6_2 desc1065(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[39:39]),.I2(s_fract_48_i[41:41]),.I3(s_fract_48_i[42:42]),.I4(s_shr2[0:0]),.I5(s_shr2[1:1]),.O6(N_88),.O5(N_16_0_i));
defparam desc1065.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_2 desc1066(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[43:43]),.I4(s_shr2[0:0]),.I5(s_shr2[1:1]),.O6(N_92),.O5(N_903_i));
defparam desc1066.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6_2 desc1067(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[41:41]),.I2(s_fract_48_i[42:42]),.I3(s_fract_48_i[43:43]),.I4(s_shl2[0:0]),.I5(s_shl2[1:1]),.O6(N_1124),.O5(N_1289));
defparam desc1067.INIT=64'hAAAACCCCF0F0FF00;
  LUT6_2 desc1068(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[41:41]),.I2(s_fract_48_i[39:39]),.I3(s_fract_48_i[42:42]),.I4(s_shl2[0:0]),.I5(s_shl2[1:1]),.O6(N_1077),.O5(N_1288));
defparam desc1068.INIT=64'hF0F0AAAACCCCFF00;
  LUT6_2 desc1069(.I0(s_fract_48_i[41:41]),.I1(s_fract_48_i[45:45]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[42:42]),.I4(N_1254),.I5(s_fract_48_i[33:33]),.O6(N_326_1),.O5(N_1247_i));
defparam desc1069.INIT=64'h1111111011111111;
  p_O_FD desc1070(.Q(s_expo1[0:0]),.D(s_expo1_5_e),.C(clk_i),.E(p_desc1070_p_O_FD));
  p_O_FD desc1071(.Q(s_shr2[0:0]),.D(s_shr2_0_e),.C(clk_i),.E(p_desc1071_p_O_FD));
  p_O_FD desc1072(.Q(s_shr2[5:5]),.D(v_shr1_4_e[5:5]),.C(clk_i),.E(p_desc1072_p_O_FD));
  p_O_FD desc1073(.Q(s_shr2[4:4]),.D(v_shr1_4_e[4:4]),.C(clk_i),.E(p_desc1073_p_O_FD));
  p_O_FD desc1074(.Q(s_shr2[3:3]),.D(v_shr1_4_e[3:3]),.C(clk_i),.E(p_desc1074_p_O_FD));
  p_O_FD desc1075(.Q(s_shr2[2:2]),.D(v_shr1_4_e[2:2]),.C(clk_i),.E(p_desc1075_p_O_FD));
  p_O_FD desc1076(.Q(s_shr2[1:1]),.D(v_shr1_4_e[1:1]),.C(clk_i),.E(p_desc1076_p_O_FD));
  p_O_FD desc1077(.Q(s_frac2a[16:16]),.D(m80_0_e),.C(clk_i),.E(p_desc1077_p_O_FD));
  p_O_FD desc1078(.Q(s_frac2a[18:18]),.D(m97_0_e),.C(clk_i),.E(p_desc1078_p_O_FD));
  p_O_FD desc1079(.Q(s_frac2a[31:31]),.D(m37_0_0_e),.C(clk_i),.E(p_desc1079_p_O_FD));
  p_O_FD desc1080(.Q(s_frac2a[21:21]),.D(m102_0_e),.C(clk_i),.E(p_desc1080_p_O_FD));
  p_O_FD desc1081(.Q(s_frac2a[22:22]),.D(m108_0_0_e),.C(clk_i),.E(p_desc1081_p_O_FD));
  p_O_FD desc1082(.Q(s_frac2a[23:23]),.D(m113_0_e),.C(clk_i),.E(p_desc1082_p_O_FD));
  p_O_FD desc1083(.Q(s_frac2a[30:30]),.D(m119_0_0_e),.C(clk_i),.E(p_desc1083_p_O_FD));
  p_O_FD desc1084(.Q(s_frac2a[29:29]),.D(m169_0_e),.C(clk_i),.E(p_desc1084_p_O_FD));
  p_O_FD desc1085(.Q(s_frac2a[20:20]),.D(m224_0_e),.C(clk_i),.E(p_desc1085_p_O_FD));
  p_O_FD desc1086(.Q(s_frac2a[26:26]),.D(m231_0_e),.C(clk_i),.E(p_desc1086_p_O_FD));
  p_O_FD desc1087(.Q(s_frac2a[28:28]),.D(m237_0_e),.C(clk_i),.E(p_desc1087_p_O_FD));
  p_O_FD desc1088(.Q(s_frac2a[19:19]),.D(m293_0_e),.C(clk_i),.E(p_desc1088_p_O_FD));
  p_O_FD desc1089(.Q(s_frac2a[17:17]),.D(m365_0_e),.C(clk_i),.E(p_desc1089_p_O_FD));
  p_O_FD desc1090(.Q(s_frac2a[25:25]),.D(m374_0_e),.C(clk_i),.E(p_desc1090_p_O_FD));
  p_O_FD desc1091(.Q(s_frac2a[27:27]),.D(m378_0_e),.C(clk_i),.E(p_desc1091_p_O_FD));
  p_O_FD desc1092(.Q(s_frac2a[24:24]),.D(m435_0_e),.C(clk_i),.E(p_desc1092_p_O_FD));
  LUT6 desc1093(.I0(N_1165),.I1(N_1168),.I2(N_169),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m435_0_e));
defparam desc1093.INIT=64'h00000000AACCAAF0;
  LUT6 desc1094(.I0(N_284),.I1(N_286),.I2(N_376),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m378_0_e));
defparam desc1094.INIT=64'h00000000CCF0CC55;
  LUT6 desc1095(.I0(N_355),.I1(N_357),.I2(N_372),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m374_0_e));
defparam desc1095.INIT=64'h00000000CCF0CCAA;
  LUT6 desc1096(.I0(N_333),.I1(N_337),.I2(N_363),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m365_0_e));
defparam desc1096.INIT=64'h00000000CCF0CCAA;
  LUT6 desc1097(.I0(N_271),.I1(N_275),.I2(N_291),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m293_0_e));
defparam desc1097.INIT=64'h0000000033F03355;
  LUT6 desc1098(.I0(N_211),.I1(N_214),.I2(N_235),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m237_0_e));
defparam desc1098.INIT=64'h00000000CCF0CC55;
  LUT6 desc1099(.I0(N_194),.I1(N_196),.I2(N_229),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m231_0_e));
defparam desc1099.INIT=64'h00000000CCF0CC55;
  LUT6 desc1100(.I0(N_217),.I1(N_221),.I2(N_223),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m224_0_e));
defparam desc1100.INIT=64'h00000000F0CCF055;
  LUT6 desc1101(.I0(s_frac2a_1_124_RNIEJB51_O6),.I1(N_1137),.I2(N_1142),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m169_0_e));
defparam desc1101.INIT=64'h00000000CCF0CC55;
  LUT6 desc1102(.I0(N_80_0),.I1(N_82_0),.I2(N_1112),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m119_0_0_e));
defparam desc1102.INIT=64'h00000000CCF0CC55;
  LUT6 desc1103(.I0(N_69_0),.I1(N_71_0_0),.I2(N_1109),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m113_0_e));
defparam desc1103.INIT=64'h00000000CCF0CC55;
  LUT6 desc1104(.I0(N_52_0),.I1(N_56_0),.I2(N_1104),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m108_0_0_e));
defparam desc1104.INIT=64'h00000000CCF0CC55;
  LUT6 desc1105(.I0(N_60_0),.I1(N_64_0),.I2(N_1098),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m102_0_e));
defparam desc1105.INIT=64'h0000000033F03355;
  LUT6 desc1106(.I0(N_1083),.I1(N_1087),.I2(N_1090),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m37_0_0_e));
defparam desc1106.INIT=64'h00000000F0CCF055;
  LUT6 desc1107(.I0(m368_lut6_2_O6),.I1(N_977),.I2(s_frac2a_1_141_RNIA10R),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m97_0_e));
defparam desc1107.INIT=64'h000000000FAA0F33;
  LUT6 desc1108(.I0(N_78_0),.I1(N_382),.I2(N_161),.I3(s_shr2[4:4]),.I4(un1_s_shr2_1_4),.I5(s_shr2[5:5]),.O(m80_0_e));
defparam desc1108.INIT=64'h0000000033AA33F0;
  LUT5 desc1109(.I0(s_zeros[0:0]),.I1(s_exp_10_i[0:0]),.I2(s_fract_48_i[47:47]),.I3(s_exp_10b[8:8]),.I4(un1_s_exp_10a_3_lut6_2_O6),.O(s_expo1_5_e));
defparam desc1109.INIT=32'hFFFFFF96;
  LUT5 desc1110(.I0(un5_v_shr1_c3),.I1(s_exp_10_i_RNIE6AQ1[2:2]),.I2(s_exp_10_i_RNI5I152[2:2]),.I3(un6_s_exp_10a),.I4(v_shr1_4[6:6]),.O(v_shr1_4_e[4:4]));
defparam desc1110.INIT=32'hFFFF2D00;
  LUT6 desc1111(.I0(un5_v_shr1_c3),.I1(s_exp_10_i_RNIE6AQ1[2:2]),.I2(s_exp_10_i_RNI5I152[2:2]),.I3(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91),.I4(un6_s_exp_10a),.I5(v_shr1_4[6:6]),.O(v_shr1_4_e[5:5]));
defparam desc1111.INIT=64'hFFFFFFFF02FD0000;
  LUT6 desc1112(.I0(s_exp_10_i[0:0]),.I1(s_fract_48_i[47:47]),.I2(un6_s_exp_10a),.I3(s_exp_10b[8:8]),.I4(un1_s_exp_10a_3_1),.I5(v_shr1_4[6:6]),.O(s_shr2_0_e));
defparam desc1112.INIT=64'hFFFFFFFF505050DC;
  LUT6 desc1113(.I0(N_173),.I1(N_481),.I2(N_503_1),.I3(N_505_1_2),.I4(N_543),.I5(s_zeros_2_2[2:2]),.O(s_zeros_2_0[2:2]));
defparam desc1113.INIT=64'hFFFFFFFFECCC0000;
  FDR desc1114(.Q(post_norm_mul_output[12:12]),.D(s_output_o_0[12:12]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1115(.I0(s_frac_rnd[12:12]),.I1(s_frac_rnd[13:13]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[12:12]));
defparam desc1115.INIT=32'h0CCC0AAA;
  FDR desc1116(.Q(post_norm_mul_output[0:0]),.D(s_output_o_0[0:0]),.C(clk_i),.R(s_output_o_sm0));
  FDR desc1117(.Q(post_norm_mul_output[1:1]),.D(s_output_o_0[1:1]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1118(.I0(s_frac_rnd[1:1]),.I1(s_frac_rnd[2:2]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[1:1]));
defparam desc1118.INIT=32'h0CCC0AAA;
  FDR desc1119(.Q(post_norm_mul_output[10:10]),.D(s_output_o_0[10:10]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1120(.I0(s_frac_rnd[10:10]),.I1(s_frac_rnd[11:11]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[10:10]));
defparam desc1120.INIT=32'h0CCC0AAA;
  FDR desc1121(.Q(post_norm_mul_output[5:5]),.D(s_output_o_0[5:5]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1122(.I0(s_frac_rnd[5:5]),.I1(s_frac_rnd[6:6]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[5:5]));
defparam desc1122.INIT=32'h0CCC0AAA;
  FDR desc1123(.Q(post_norm_mul_output[4:4]),.D(s_output_o_0[4:4]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1124(.I0(s_frac_rnd[4:4]),.I1(s_frac_rnd[5:5]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[4:4]));
defparam desc1124.INIT=32'h0CCC0AAA;
  FDR desc1125(.Q(post_norm_mul_output[19:19]),.D(s_output_o_0[19:19]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1126(.I0(s_frac_rnd[19:19]),.I1(s_frac_rnd[20:20]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[19:19]));
defparam desc1126.INIT=32'h0CCC0AAA;
  FDR desc1127(.Q(post_norm_mul_output[15:15]),.D(s_output_o_0[15:15]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1128(.I0(s_frac_rnd[15:15]),.I1(s_frac_rnd[16:16]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[15:15]));
defparam desc1128.INIT=32'h0CCC0AAA;
  FDR desc1129(.Q(post_norm_mul_output[2:2]),.D(s_output_o_0[2:2]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1130(.I0(s_frac_rnd[2:2]),.I1(s_frac_rnd[3:3]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[2:2]));
defparam desc1130.INIT=32'h0CCC0AAA;
  FDR desc1131(.Q(post_norm_mul_output[7:7]),.D(s_output_o_0[7:7]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1132(.I0(s_frac_rnd[7:7]),.I1(s_frac_rnd[8:8]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[7:7]));
defparam desc1132.INIT=32'h0CCC0AAA;
  FDR desc1133(.Q(post_norm_mul_output[20:20]),.D(s_output_o_0[20:20]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1134(.I0(s_frac_rnd[20:20]),.I1(s_frac_rnd[21:21]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[20:20]));
defparam desc1134.INIT=32'h0CCC0AAA;
  FDR desc1135(.Q(post_norm_mul_output[3:3]),.D(s_output_o_0[3:3]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1136(.I0(s_frac_rnd[3:3]),.I1(s_frac_rnd[4:4]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[3:3]));
defparam desc1136.INIT=32'h0CCC0AAA;
  FDR desc1137(.Q(post_norm_mul_output[13:13]),.D(s_output_o_0[13:13]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1138(.I0(s_frac_rnd[13:13]),.I1(s_frac_rnd[14:14]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[13:13]));
defparam desc1138.INIT=32'h0CCC0AAA;
  FDR desc1139(.Q(post_norm_mul_output[14:14]),.D(s_output_o_0[14:14]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1140(.I0(s_frac_rnd[14:14]),.I1(s_frac_rnd[15:15]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[14:14]));
defparam desc1140.INIT=32'h0CCC0AAA;
  FDR desc1141(.Q(post_norm_mul_output[8:8]),.D(s_output_o_0[8:8]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1142(.I0(s_frac_rnd[8:8]),.I1(s_frac_rnd[9:9]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[8:8]));
defparam desc1142.INIT=32'h0CCC0AAA;
  FDR desc1143(.Q(post_norm_mul_output[17:17]),.D(s_output_o_0[17:17]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1144(.I0(s_frac_rnd[17:17]),.I1(s_frac_rnd[18:18]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[17:17]));
defparam desc1144.INIT=32'h0CCC0AAA;
  FDR desc1145(.Q(post_norm_mul_output[21:21]),.D(s_output_o_0[21:21]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1146(.I0(s_frac_rnd[21:21]),.I1(s_frac_rnd[22:22]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[21:21]));
defparam desc1146.INIT=32'h0CCC0AAA;
  FDR desc1147(.Q(post_norm_mul_output[11:11]),.D(s_output_o_0[11:11]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1148(.I0(s_frac_rnd[11:11]),.I1(s_frac_rnd[12:12]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[11:11]));
defparam desc1148.INIT=32'h0CCC0AAA;
  FDR desc1149(.Q(post_norm_mul_output[6:6]),.D(s_output_o_0[6:6]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1150(.I0(s_frac_rnd[6:6]),.I1(s_frac_rnd[7:7]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[6:6]));
defparam desc1150.INIT=32'h0CCC0AAA;
  FDR desc1151(.Q(post_norm_mul_output[18:18]),.D(s_output_o_0[18:18]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1152(.I0(s_frac_rnd[18:18]),.I1(s_frac_rnd[19:19]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[18:18]));
defparam desc1152.INIT=32'h0CCC0AAA;
  FDR desc1153(.Q(post_norm_mul_output[9:9]),.D(s_output_o_0[9:9]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1154(.I0(s_frac_rnd[9:9]),.I1(s_frac_rnd[10:10]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[9:9]));
defparam desc1154.INIT=32'h0CCC0AAA;
  FDR desc1155(.Q(post_norm_mul_output[16:16]),.D(s_output_o_0[16:16]),.C(clk_i),.R(s_output_o_sm0));
  LUT5 desc1156(.I0(s_frac_rnd[16:16]),.I1(s_frac_rnd[17:17]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.O(s_output_o_0[16:16]));
defparam desc1156.INIT=32'h0CCC0AAA;
  LUT6 desc1157(.I0(N_247),.I1(N_1247),.I2(N_1249),.I3(N_1261),.I4(N_1277),.I5(N_1372),.O(s_zeros_2_0[3:3]));
defparam desc1157.INIT=64'h0003000200030000;
  LUT6 desc1158(.I0(N_315),.I1(N_1251),.I2(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I3(N_1277),.I4(N_1372),.I5(s_fract_48_i[15:15]),.O(N_414_i_0));
defparam desc1158.INIT=64'h0055005500540055;
  LUT6 desc1159(.I0(s_fract_48_i[38:38]),.I1(v_count_0_sqmuxa_47_0),.I2(v_count_0_sqmuxa_47_1_0),.I3(v_count_0_sqmuxa_47_3_3),.I4(v_count_0_sqmuxa_47_3_4),.I5(v_count_0_sqmuxa_47_4_4),.O(v_count_0_sqmuxa_47_1));
defparam desc1159.INIT=64'h4000000000000000;
  LUT6 desc1160(.I0(N_23_0_3),.I1(N_23_0_4),.I2(N_23_4),.I3(N_1247),.I4(s_fract_48_i[40:40]),.I5(s_fract_48_i[43:43]),.O(N_23_i_0));
defparam desc1160.INIT=64'h0101010101000101;
  LUT6 desc1161(.I0(N_62_1),.I1(N_425),.I2(N_1254),.I3(s_fract_48_i[43:43]),.I4(s_fract_48_i[44:44]),.I5(s_fract_48_i[45:45]),.O(N_62_i_0));
defparam desc1161.INIT=64'h0000000005050501;
  LUT2 s_expo2b_axb_1_cZ(.I0(s_expo1[1:1]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_1));
defparam s_expo2b_axb_1_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_2_cZ(.I0(s_expo1[2:2]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_2));
defparam s_expo2b_axb_2_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_3_cZ(.I0(s_expo1[3:3]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_3));
defparam s_expo2b_axb_3_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_4_cZ(.I0(s_expo1[4:4]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_4));
defparam s_expo2b_axb_4_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_5_cZ(.I0(s_expo1[5:5]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_5));
defparam s_expo2b_axb_5_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_6_cZ(.I0(s_expo1[6:6]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_6));
defparam s_expo2b_axb_6_cZ.INIT=4'h9;
  LUT4 desc1162(.I0(s_exp_10_i[0:0]),.I1(s_exp_10_i[1:1]),.I2(s_fract_48_i[47:47]),.I3(s_zeros[1:1]),.O(s_exp_10b_axb_1));
defparam desc1162.INIT=16'h6C93;
  LUT1 s_frac_rnd_3_0_axb_1_cZ(.I0(s_frac2a[24:24]),.O(s_frac_rnd_3_0_axb_1));
defparam s_frac_rnd_3_0_axb_1_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_2_cZ(.I0(s_frac2a[25:25]),.O(s_frac_rnd_3_0_axb_2));
defparam s_frac_rnd_3_0_axb_2_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_3_cZ(.I0(s_frac2a[26:26]),.O(s_frac_rnd_3_0_axb_3));
defparam s_frac_rnd_3_0_axb_3_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_4_cZ(.I0(s_frac2a[27:27]),.O(s_frac_rnd_3_0_axb_4));
defparam s_frac_rnd_3_0_axb_4_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_5_cZ(.I0(s_frac2a[28:28]),.O(s_frac_rnd_3_0_axb_5));
defparam s_frac_rnd_3_0_axb_5_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_6_cZ(.I0(s_frac2a[29:29]),.O(s_frac_rnd_3_0_axb_6));
defparam s_frac_rnd_3_0_axb_6_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_7_cZ(.I0(s_frac2a[30:30]),.O(s_frac_rnd_3_0_axb_7));
defparam s_frac_rnd_3_0_axb_7_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_8_cZ(.I0(s_frac2a[31:31]),.O(s_frac_rnd_3_0_axb_8));
defparam s_frac_rnd_3_0_axb_8_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_9_cZ(.I0(s_frac2a[32:32]),.O(s_frac_rnd_3_0_axb_9));
defparam s_frac_rnd_3_0_axb_9_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_10_cZ(.I0(s_frac2a[33:33]),.O(s_frac_rnd_3_0_axb_10));
defparam s_frac_rnd_3_0_axb_10_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_11_cZ(.I0(s_frac2a[34:34]),.O(s_frac_rnd_3_0_axb_11));
defparam s_frac_rnd_3_0_axb_11_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_12_cZ(.I0(s_frac2a[35:35]),.O(s_frac_rnd_3_0_axb_12));
defparam s_frac_rnd_3_0_axb_12_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_13_cZ(.I0(s_frac2a[36:36]),.O(s_frac_rnd_3_0_axb_13));
defparam s_frac_rnd_3_0_axb_13_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_14_cZ(.I0(s_frac2a[37:37]),.O(s_frac_rnd_3_0_axb_14));
defparam s_frac_rnd_3_0_axb_14_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_15_cZ(.I0(s_frac2a[38:38]),.O(s_frac_rnd_3_0_axb_15));
defparam s_frac_rnd_3_0_axb_15_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_16_cZ(.I0(s_frac2a[39:39]),.O(s_frac_rnd_3_0_axb_16));
defparam s_frac_rnd_3_0_axb_16_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_17_cZ(.I0(s_frac2a[40:40]),.O(s_frac_rnd_3_0_axb_17));
defparam s_frac_rnd_3_0_axb_17_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_18_cZ(.I0(s_frac2a[41:41]),.O(s_frac_rnd_3_0_axb_18));
defparam s_frac_rnd_3_0_axb_18_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_19_cZ(.I0(s_frac2a[42:42]),.O(s_frac_rnd_3_0_axb_19));
defparam s_frac_rnd_3_0_axb_19_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_20_cZ(.I0(s_frac2a[43:43]),.O(s_frac_rnd_3_0_axb_20));
defparam s_frac_rnd_3_0_axb_20_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_21_cZ(.I0(s_frac2a[44:44]),.O(s_frac_rnd_3_0_axb_21));
defparam s_frac_rnd_3_0_axb_21_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_22_cZ(.I0(s_frac2a[45:45]),.O(s_frac_rnd_3_0_axb_22));
defparam s_frac_rnd_3_0_axb_22_cZ.INIT=2'h2;
  LUT1 s_frac_rnd_3_0_axb_23_cZ(.I0(s_frac2a[46:46]),.O(s_frac_rnd_3_0_axb_23));
defparam s_frac_rnd_3_0_axb_23_cZ.INIT=2'h2;
  p_O_FD desc1163(.Q(s_exp_10_i[1:1]),.D(pre_norm_mul_exp_10[1:1]),.C(clk_i),.E(p_desc1163_p_O_FD));
  p_O_FD desc1164(.Q(s_exp_10_i[2:2]),.D(pre_norm_mul_exp_10[2:2]),.C(clk_i),.E(p_desc1164_p_O_FD));
  p_O_FD desc1165(.Q(s_exp_10_i[3:3]),.D(pre_norm_mul_exp_10[3:3]),.C(clk_i),.E(p_desc1165_p_O_FD));
  p_O_FD desc1166(.Q(s_exp_10_i[4:4]),.D(pre_norm_mul_exp_10[4:4]),.C(clk_i),.E(p_desc1166_p_O_FD));
  p_O_FD desc1167(.Q(s_exp_10_i[5:5]),.D(pre_norm_mul_exp_10[5:5]),.C(clk_i),.E(p_desc1167_p_O_FD));
  p_O_FD desc1168(.Q(s_exp_10_i[6:6]),.D(pre_norm_mul_exp_10[6:6]),.C(clk_i),.E(p_desc1168_p_O_FD));
  p_O_FD desc1169(.Q(s_exp_10_i[7:7]),.D(pre_norm_mul_exp_10[7:7]),.C(clk_i),.E(p_desc1169_p_O_FD));
  p_O_FD desc1170(.Q(s_exp_10_i[8:8]),.D(pre_norm_mul_exp_10[8:8]),.C(clk_i),.E(p_desc1170_p_O_FD));
  p_O_FD desc1171(.Q(s_exp_10_i[9:9]),.D(pre_norm_mul_exp_10[9:9]),.C(clk_i),.E(p_desc1171_p_O_FD));
  p_O_FD desc1172(.Q(s_exp_10_i[0:0]),.D(pre_norm_mul_exp_10[0:0]),.C(clk_i),.E(p_desc1172_p_O_FD));
  p_O_FD desc1173(.Q(s_frac2a[6:6]),.D(s_frac2a_3[6:6]),.C(clk_i),.E(p_desc1173_p_O_FD));
  p_O_FD desc1174(.Q(s_frac2a[7:7]),.D(s_frac2a_3[7:7]),.C(clk_i),.E(p_desc1174_p_O_FD));
  p_O_FD desc1175(.Q(s_frac2a[8:8]),.D(s_frac2a_3[8:8]),.C(clk_i),.E(p_desc1175_p_O_FD));
  p_O_FD desc1176(.Q(s_frac2a[9:9]),.D(s_frac2a_3[9:9]),.C(clk_i),.E(p_desc1176_p_O_FD));
  p_O_FD desc1177(.Q(s_frac2a[10:10]),.D(s_frac2a_3[10:10]),.C(clk_i),.E(p_desc1177_p_O_FD));
  p_O_FD desc1178(.Q(s_frac2a[11:11]),.D(s_frac2a_3[11:11]),.C(clk_i),.E(p_desc1178_p_O_FD));
  p_O_FD desc1179(.Q(s_frac2a[12:12]),.D(s_frac2a_3[12:12]),.C(clk_i),.E(p_desc1179_p_O_FD));
  p_O_FD desc1180(.Q(s_frac2a[13:13]),.D(s_frac2a_3[13:13]),.C(clk_i),.E(p_desc1180_p_O_FD));
  p_O_FD desc1181(.Q(s_frac2a[14:14]),.D(s_frac2a_3[14:14]),.C(clk_i),.E(p_desc1181_p_O_FD));
  p_O_FD desc1182(.Q(s_frac2a[15:15]),.D(s_frac2a_3[15:15]),.C(clk_i),.E(p_desc1182_p_O_FD));
  p_O_FD desc1183(.Q(post_norm_mul_output[31:31]),.D(s_sign_i),.C(clk_i),.E(p_desc1183_p_O_FD));
  p_O_FD desc1184(.Q(s_frac2a[0:0]),.D(s_frac2a_3[0:0]),.C(clk_i),.E(p_desc1184_p_O_FD));
  p_O_FD desc1185(.Q(s_frac2a[1:1]),.D(s_frac2a_3[1:1]),.C(clk_i),.E(p_desc1185_p_O_FD));
  p_O_FD desc1186(.Q(s_frac2a[2:2]),.D(s_frac2a_3[2:2]),.C(clk_i),.E(p_desc1186_p_O_FD));
  p_O_FD desc1187(.Q(s_frac2a[3:3]),.D(s_frac2a_3[3:3]),.C(clk_i),.E(p_desc1187_p_O_FD));
  p_O_FD desc1188(.Q(s_frac2a[4:4]),.D(s_frac2a_3[4:4]),.C(clk_i),.E(p_desc1188_p_O_FD));
  p_O_FD desc1189(.Q(s_frac2a[5:5]),.D(s_frac2a_3[5:5]),.C(clk_i),.E(p_desc1189_p_O_FD));
  p_O_FD desc1190(.Q(post_norm_mul_output[22:22]),.D(s_output_o[22:22]),.C(clk_i),.E(p_desc1190_p_O_FD));
  p_O_FD desc1191(.Q(s_frac_rnd[18:18]),.D(s_frac_rnd_3[18:18]),.C(clk_i),.E(p_desc1191_p_O_FD));
  p_O_FD desc1192(.Q(s_frac_rnd[19:19]),.D(s_frac_rnd_3[19:19]),.C(clk_i),.E(p_desc1192_p_O_FD));
  p_O_FD desc1193(.Q(s_frac_rnd[20:20]),.D(s_frac_rnd_3[20:20]),.C(clk_i),.E(p_desc1193_p_O_FD));
  p_O_FD desc1194(.Q(s_frac_rnd[21:21]),.D(s_frac_rnd_3[21:21]),.C(clk_i),.E(p_desc1194_p_O_FD));
  p_O_FD desc1195(.Q(s_frac_rnd[22:22]),.D(s_frac_rnd_3[22:22]),.C(clk_i),.E(p_desc1195_p_O_FD));
  p_O_FD desc1196(.Q(s_frac_rnd[23:23]),.D(s_frac_rnd_3[23:23]),.C(clk_i),.E(p_desc1196_p_O_FD));
  p_O_FD desc1197(.Q(s_frac_rnd[24:24]),.D(s_frac_rnd_3[24:24]),.C(clk_i),.E(p_desc1197_p_O_FD));
  p_O_FD desc1198(.Q(s_frac_rnd[3:3]),.D(s_frac_rnd_3[3:3]),.C(clk_i),.E(p_desc1198_p_O_FD));
  p_O_FD desc1199(.Q(s_frac_rnd[4:4]),.D(s_frac_rnd_3[4:4]),.C(clk_i),.E(p_desc1199_p_O_FD));
  p_O_FD desc1200(.Q(s_frac_rnd[5:5]),.D(s_frac_rnd_3[5:5]),.C(clk_i),.E(p_desc1200_p_O_FD));
  p_O_FD desc1201(.Q(s_frac_rnd[6:6]),.D(s_frac_rnd_3[6:6]),.C(clk_i),.E(p_desc1201_p_O_FD));
  p_O_FD desc1202(.Q(s_frac_rnd[7:7]),.D(s_frac_rnd_3[7:7]),.C(clk_i),.E(p_desc1202_p_O_FD));
  p_O_FD desc1203(.Q(s_frac_rnd[8:8]),.D(s_frac_rnd_3[8:8]),.C(clk_i),.E(p_desc1203_p_O_FD));
  p_O_FD desc1204(.Q(s_frac_rnd[9:9]),.D(s_frac_rnd_3[9:9]),.C(clk_i),.E(p_desc1204_p_O_FD));
  p_O_FD desc1205(.Q(s_frac_rnd[10:10]),.D(s_frac_rnd_3[10:10]),.C(clk_i),.E(p_desc1205_p_O_FD));
  p_O_FD desc1206(.Q(s_frac_rnd[11:11]),.D(s_frac_rnd_3[11:11]),.C(clk_i),.E(p_desc1206_p_O_FD));
  p_O_FD desc1207(.Q(s_frac_rnd[12:12]),.D(s_frac_rnd_3[12:12]),.C(clk_i),.E(p_desc1207_p_O_FD));
  p_O_FD desc1208(.Q(s_frac_rnd[13:13]),.D(s_frac_rnd_3[13:13]),.C(clk_i),.E(p_desc1208_p_O_FD));
  p_O_FD desc1209(.Q(s_frac_rnd[14:14]),.D(s_frac_rnd_3[14:14]),.C(clk_i),.E(p_desc1209_p_O_FD));
  p_O_FD desc1210(.Q(s_frac_rnd[15:15]),.D(s_frac_rnd_3[15:15]),.C(clk_i),.E(p_desc1210_p_O_FD));
  p_O_FD desc1211(.Q(s_frac_rnd[16:16]),.D(s_frac_rnd_3[16:16]),.C(clk_i),.E(p_desc1211_p_O_FD));
  p_O_FD desc1212(.Q(s_frac_rnd[17:17]),.D(s_frac_rnd_3[17:17]),.C(clk_i),.E(p_desc1212_p_O_FD));
  p_O_FD desc1213(.Q(s_frac_rnd[0:0]),.D(s_frac_rnd_3[0:0]),.C(clk_i),.E(p_desc1213_p_O_FD));
  p_O_FD desc1214(.Q(s_frac_rnd[1:1]),.D(s_frac_rnd_3[1:1]),.C(clk_i),.E(p_desc1214_p_O_FD));
  p_O_FD desc1215(.Q(s_frac_rnd[2:2]),.D(s_frac_rnd_3[2:2]),.C(clk_i),.E(p_desc1215_p_O_FD));
  p_O_FD desc1216(.Q(s_zeros[0:0]),.D(N_23_i_0),.C(clk_i),.E(p_desc1216_p_O_FD));
  p_O_FD desc1217(.Q(s_zeros[1:1]),.D(N_62_i_0),.C(clk_i),.E(p_desc1217_p_O_FD));
  p_O_FD desc1218(.Q(s_zeros[2:2]),.D(s_zeros_2_0[2:2]),.C(clk_i),.E(p_desc1218_p_O_FD));
  p_O_FD desc1219(.Q(s_zeros[3:3]),.D(s_zeros_2_0[3:3]),.C(clk_i),.E(p_desc1219_p_O_FD));
  p_O_FD desc1220(.Q(s_zeros[4:4]),.D(N_414_i_0),.C(clk_i),.E(p_desc1220_p_O_FD));
  p_O_FD desc1221(.Q(s_zeros[5:5]),.D(v_count_0_sqmuxa_47_1),.C(clk_i),.E(p_desc1221_p_O_FD));
  p_O_FD s_sign_i_Z(.Q(s_sign_i),.D(N_6_i),.C(clk_i),.E(p_s_sign_i_Z_p_O_FD));
  p_O_FD ine_o_Z(.Q(post_norm_mul_ine),.D(un1_s_ine_o),.C(clk_i),.E(p_ine_o_Z_p_O_FD));
  FDR desc1222(.Q(s_shl2[1:1]),.D(N_715),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  FDR desc1223(.Q(s_shl2[2:2]),.D(N_716),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  FDR desc1224(.Q(s_shl2[3:3]),.D(N_717),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  FDR desc1225(.Q(s_shl2[4:4]),.D(N_718),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  FDR desc1226(.Q(s_shl2[5:5]),.D(N_719),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  FDR desc1227(.Q(s_frac2a[36:36]),.D(N_406),.C(clk_i),.R(N_459_i));
  FDR desc1228(.Q(s_frac2a[37:37]),.D(N_411),.C(clk_i),.R(N_459_i));
  FDR desc1229(.Q(s_frac2a[38:38]),.D(N_1117),.C(clk_i),.R(N_459_i));
  FDR desc1230(.Q(s_frac2a[39:39]),.D(N_1148),.C(clk_i),.R(N_459_i));
  FDR desc1231(.Q(s_frac2a[40:40]),.D(N_441),.C(clk_i),.R(N_459_i));
  FDR desc1232(.Q(s_frac2a[41:41]),.D(N_1160),.C(clk_i),.R(N_459_i));
  FDR desc1233(.Q(s_frac2a[42:42]),.D(N_245),.C(clk_i),.R(N_459_i));
  FDR desc1234(.Q(s_frac2a[43:43]),.D(N_308),.C(clk_i),.R(N_459_i));
  FDR desc1235(.Q(s_frac2a[44:44]),.D(N_256),.C(clk_i),.R(N_459_i));
  FDR desc1236(.Q(s_frac2a[45:45]),.D(N_184),.C(clk_i),.R(N_459_i));
  FDR desc1237(.Q(s_frac2a[46:46]),.D(N_1123),.C(clk_i),.R(N_459_i));
  FDR desc1238(.Q(s_frac2a[47:47]),.D(N_1131),.C(clk_i),.R(N_459_i));
  FDR desc1239(.Q(s_frac2a[32:32]),.D(N_389),.C(clk_i),.R(N_459_i));
  FDR desc1240(.Q(s_frac2a[33:33]),.D(N_396),.C(clk_i),.R(N_459_i));
  FDR desc1241(.Q(s_frac2a[34:34]),.D(N_401),.C(clk_i),.R(N_459_i));
  FDR desc1242(.Q(s_frac2a[35:35]),.D(N_300),.C(clk_i),.R(N_459_i));
  FDR desc1243(.Q(s_shl2[0:0]),.D(N_714),.C(clk_i),.R(s_exp_10b_s_1_RNI0PGD1_O6));
  p_O_FD desc1244(.Q(s_fract_48_i[47:47]),.D(mul_24_fract_48[47:47]),.C(clk_i),.E(p_desc1244_p_O_FD));
  p_O_FD desc1245(.Q(s_fract_48_i[46:46]),.D(mul_24_fract_48[46:46]),.C(clk_i),.E(p_desc1245_p_O_FD));
  p_O_FD desc1246(.Q(s_fract_48_i[45:45]),.D(mul_24_fract_48[45:45]),.C(clk_i),.E(p_desc1246_p_O_FD));
  p_O_FD desc1247(.Q(s_fract_48_i[44:44]),.D(mul_24_fract_48[44:44]),.C(clk_i),.E(p_desc1247_p_O_FD));
  p_O_FD desc1248(.Q(s_fract_48_i[43:43]),.D(mul_24_fract_48[43:43]),.C(clk_i),.E(p_desc1248_p_O_FD));
  p_O_FD desc1249(.Q(s_fract_48_i[42:42]),.D(mul_24_fract_48[42:42]),.C(clk_i),.E(p_desc1249_p_O_FD));
  p_O_FD desc1250(.Q(s_fract_48_i[41:41]),.D(mul_24_fract_48[41:41]),.C(clk_i),.E(p_desc1250_p_O_FD));
  p_O_FD desc1251(.Q(s_fract_48_i[40:40]),.D(mul_24_fract_48[40:40]),.C(clk_i),.E(p_desc1251_p_O_FD));
  p_O_FD desc1252(.Q(s_fract_48_i[39:39]),.D(mul_24_fract_48[39:39]),.C(clk_i),.E(p_desc1252_p_O_FD));
  p_O_FD desc1253(.Q(s_fract_48_i[38:38]),.D(mul_24_fract_48[38:38]),.C(clk_i),.E(p_desc1253_p_O_FD));
  p_O_FD desc1254(.Q(s_fract_48_i[37:37]),.D(mul_24_fract_48[37:37]),.C(clk_i),.E(p_desc1254_p_O_FD));
  p_O_FD desc1255(.Q(s_fract_48_i[36:36]),.D(mul_24_fract_48[36:36]),.C(clk_i),.E(p_desc1255_p_O_FD));
  p_O_FD desc1256(.Q(s_fract_48_i[35:35]),.D(mul_24_fract_48[35:35]),.C(clk_i),.E(p_desc1256_p_O_FD));
  p_O_FD desc1257(.Q(s_fract_48_i[34:34]),.D(mul_24_fract_48[34:34]),.C(clk_i),.E(p_desc1257_p_O_FD));
  p_O_FD desc1258(.Q(s_fract_48_i[33:33]),.D(mul_24_fract_48[33:33]),.C(clk_i),.E(p_desc1258_p_O_FD));
  p_O_FD desc1259(.Q(s_fract_48_i[32:32]),.D(mul_24_fract_48[32:32]),.C(clk_i),.E(p_desc1259_p_O_FD));
  p_O_FD desc1260(.Q(s_fract_48_i[31:31]),.D(mul_24_fract_48[31:31]),.C(clk_i),.E(p_desc1260_p_O_FD));
  p_O_FD desc1261(.Q(s_fract_48_i[30:30]),.D(mul_24_fract_48[30:30]),.C(clk_i),.E(p_desc1261_p_O_FD));
  p_O_FD desc1262(.Q(s_fract_48_i[29:29]),.D(mul_24_fract_48[29:29]),.C(clk_i),.E(p_desc1262_p_O_FD));
  p_O_FD desc1263(.Q(s_fract_48_i[28:28]),.D(mul_24_fract_48[28:28]),.C(clk_i),.E(p_desc1263_p_O_FD));
  p_O_FD desc1264(.Q(s_fract_48_i[27:27]),.D(mul_24_fract_48[27:27]),.C(clk_i),.E(p_desc1264_p_O_FD));
  p_O_FD desc1265(.Q(s_fract_48_i[26:26]),.D(mul_24_fract_48[26:26]),.C(clk_i),.E(p_desc1265_p_O_FD));
  p_O_FD desc1266(.Q(s_fract_48_i[25:25]),.D(mul_24_fract_48[25:25]),.C(clk_i),.E(p_desc1266_p_O_FD));
  p_O_FD desc1267(.Q(s_fract_48_i[24:24]),.D(mul_24_fract_48[24:24]),.C(clk_i),.E(p_desc1267_p_O_FD));
  p_O_FD desc1268(.Q(s_fract_48_i[23:23]),.D(mul_24_fract_48[23:23]),.C(clk_i),.E(p_desc1268_p_O_FD));
  p_O_FD desc1269(.Q(s_fract_48_i[22:22]),.D(mul_24_fract_48[22:22]),.C(clk_i),.E(p_desc1269_p_O_FD));
  p_O_FD desc1270(.Q(s_fract_48_i[21:21]),.D(mul_24_fract_48[21:21]),.C(clk_i),.E(p_desc1270_p_O_FD));
  p_O_FD desc1271(.Q(s_fract_48_i[20:20]),.D(mul_24_fract_48[20:20]),.C(clk_i),.E(p_desc1271_p_O_FD));
  p_O_FD desc1272(.Q(s_fract_48_i[19:19]),.D(mul_24_fract_48[19:19]),.C(clk_i),.E(p_desc1272_p_O_FD));
  p_O_FD desc1273(.Q(s_fract_48_i[18:18]),.D(mul_24_fract_48[18:18]),.C(clk_i),.E(p_desc1273_p_O_FD));
  p_O_FD desc1274(.Q(s_fract_48_i[17:17]),.D(mul_24_fract_48[17:17]),.C(clk_i),.E(p_desc1274_p_O_FD));
  p_O_FD desc1275(.Q(s_fract_48_i[16:16]),.D(mul_24_fract_48[16:16]),.C(clk_i),.E(p_desc1275_p_O_FD));
  p_O_FD desc1276(.Q(s_fract_48_i[15:15]),.D(mul_24_fract_48[15:15]),.C(clk_i),.E(p_desc1276_p_O_FD));
  p_O_FD desc1277(.Q(s_fract_48_i[14:14]),.D(mul_24_fract_48[14:14]),.C(clk_i),.E(p_desc1277_p_O_FD));
  p_O_FD desc1278(.Q(s_fract_48_i[13:13]),.D(mul_24_fract_48[13:13]),.C(clk_i),.E(p_desc1278_p_O_FD));
  p_O_FD desc1279(.Q(s_fract_48_i[12:12]),.D(mul_24_fract_48[12:12]),.C(clk_i),.E(p_desc1279_p_O_FD));
  p_O_FD desc1280(.Q(s_fract_48_i[11:11]),.D(mul_24_fract_48[11:11]),.C(clk_i),.E(p_desc1280_p_O_FD));
  p_O_FD desc1281(.Q(s_fract_48_i[10:10]),.D(mul_24_fract_48[10:10]),.C(clk_i),.E(p_desc1281_p_O_FD));
  p_O_FD desc1282(.Q(s_fract_48_i[9:9]),.D(mul_24_fract_48[9:9]),.C(clk_i),.E(p_desc1282_p_O_FD));
  p_O_FD desc1283(.Q(s_fract_48_i[8:8]),.D(mul_24_fract_48[8:8]),.C(clk_i),.E(p_desc1283_p_O_FD));
  p_O_FD desc1284(.Q(s_fract_48_i[7:7]),.D(mul_24_fract_48[7:7]),.C(clk_i),.E(p_desc1284_p_O_FD));
  p_O_FD desc1285(.Q(s_fract_48_i[6:6]),.D(mul_24_fract_48[6:6]),.C(clk_i),.E(p_desc1285_p_O_FD));
  p_O_FD desc1286(.Q(s_fract_48_i[5:5]),.D(mul_24_fract_48[5:5]),.C(clk_i),.E(p_desc1286_p_O_FD));
  p_O_FD desc1287(.Q(s_fract_48_i[4:4]),.D(mul_24_fract_48[4:4]),.C(clk_i),.E(p_desc1287_p_O_FD));
  p_O_FD desc1288(.Q(s_fract_48_i[3:3]),.D(mul_24_fract_48[3:3]),.C(clk_i),.E(p_desc1288_p_O_FD));
  p_O_FD desc1289(.Q(s_fract_48_i[2:2]),.D(mul_24_fract_48[2:2]),.C(clk_i),.E(p_desc1289_p_O_FD));
  p_O_FD desc1290(.Q(s_fract_48_i[1:1]),.D(mul_24_fract_48[1:1]),.C(clk_i),.E(p_desc1290_p_O_FD));
  p_O_FD desc1291(.Q(s_fract_48_i[0:0]),.D(mul_24_fract_48[0:0]),.C(clk_i),.E(p_desc1291_p_O_FD));
  LUT6 desc1292(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[41:41]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[42:42]),.I4(s_fract_48_i[47:47]),.I5(N_1249),.O(N_315));
defparam desc1292.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc1293(.I0(s_zeros[1:1]),.I1(s_zeros[0:0]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_fract_48_i[47:47]),.I5(un1_s_exp_10a_3_1),.LO(N_715));
defparam desc1293.INIT=64'hA569695AAAAAAAAA;
  LUT4_L desc1294(.I0(s_zeros[0:0]),.I1(s_exp_10_i[0:0]),.I2(s_fract_48_i[47:47]),.I3(un1_s_exp_10a_3_1),.LO(N_714));
defparam desc1294.INIT=16'h96AA;
  LUT6_L desc1295(.I0(s_fract_48_i[7:7]),.I1(s_fract_48_i[38:38]),.I2(s_fract_48_i[39:39]),.I3(s_fract_48_i[32:32]),.I4(s_fract_48_i[33:33]),.I5(N_709),.LO(N_331_0_4));
defparam desc1295.INIT=64'h0000000000000001;
  LUT6 desc1296(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[38:38]),.I2(s_fract_48_i[45:45]),.I3(N_1317),.I4(N_1254),.I5(N_1353),.O(N_23_4));
defparam desc1296.INIT=64'hFFFFFFCEFFFFFF0A;
  LUT6_L desc1297(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[39:39]),.I2(N_464_1),.I3(N_301),.I4(N_1328),.I5(N_535),.LO(N_503_1));
defparam desc1297.INIT=64'hEEEEEEFFE0E0E0F0;
  LUT6_L desc1298(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[35:35]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(N_37),.I5(N_693),.LO(N_700_1));
defparam desc1298.INIT=64'hFFFF0000FFFE0000;
  LUT6 desc1299(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[15:15]),.I4(s_fract_48_i[25:25]),.I5(N_320_0_3),.O(N_320_0));
defparam desc1299.INIT=64'h0000000100000000;
  LUT5_L desc1300(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(un1_s_expo3),.LO(s_output_o_m0[23:23]));
defparam desc1300.INIT=32'h06660999;
  LUT6_L desc1301(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.I2(s_r_zeros[4:4]),.I3(s_r_zeros[5:5]),.I4(s_expo2b[1:1]),.I5(un1_s_expo3),.LO(s_output_o_m0[24:24]));
defparam desc1301.INIT=64'h066609990FFF0000;
  LUT5_L desc1302(.I0(s_r_zeros[4:4]),.I1(s_r_zeros[5:5]),.I2(s_expo2b[4:4]),.I3(un7_s_expo3_c4),.I4(un1_s_expo3),.LO(s_output_o_m0[27:27]));
defparam desc1302.INIT=32'h07707070;
  LUT6_L desc1303(.I0(s_r_zeros[4:4]),.I1(s_r_zeros[5:5]),.I2(s_expo2b[4:4]),.I3(s_expo2b[5:5]),.I4(un7_s_expo3_c4),.I5(un1_s_expo3),.LO(s_output_o_m0[28:28]));
defparam desc1303.INIT=64'h0770770077007700;
  LUT3_L desc1304(.I0(s_r_zeros[4:4]),.I1(s_r_zeros[5:5]),.I2(s_expo3[7:7]),.LO(s_output_o_m0[30:30]));
defparam desc1304.INIT=8'h70;
  LUT6_L desc1305(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.I4(N_286),.I5(N_307),.LO(N_308));
defparam desc1305.INIT=64'hFFFF0001FFFE0000;
  LUT6_L desc1306(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.I4(N_275),.I5(N_299),.LO(N_300));
defparam desc1306.INIT=64'h0001FFFF0000FFFE;
  LUT6_L desc1307(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.I4(N_71_0_0),.I5(N_1147),.LO(N_1148));
defparam desc1307.INIT=64'hFFFF0001FFFE0000;
  LUT6_L desc1308(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.I4(N_64_0),.I5(N_410),.LO(N_411));
defparam desc1308.INIT=64'h0001FFFF0000FFFE;
  LUT5 desc1309(.I0(s_fract_48_i[12:12]),.I1(s_fract_48_i[8:8]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[2:2]),.I4(N_673),.O(N_679));
defparam desc1309.INIT=32'h00010000;
  LUT6 desc1310(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[26:26]),.I2(s_fract_48_i[24:24]),.I3(s_fract_48_i[29:29]),.I4(s_fract_48_i[25:25]),.I5(N_1364),.O(N_1372));
defparam desc1310.INIT=64'h0000000100000000;
  LUT6 desc1311(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[26:26]),.I2(s_fract_48_i[24:24]),.I3(s_fract_48_i[27:27]),.I4(s_fract_48_i[31:31]),.I5(s_fract_48_i[25:25]),.O(N_611));
defparam desc1311.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc1312(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[2:2]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[29:29]),.I4(N_597),.I5(N_700_1),.LO(N_637));
defparam desc1312.INIT=64'hFFFFEEEFFFFF0000;
  LUT6_L desc1313(.I0(s_fract_48_i[23:23]),.I1(s_fract_48_i[28:28]),.I2(s_fract_48_i[29:29]),.I3(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I4(N_1251),.I5(N_611),.LO(N_624));
defparam desc1313.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc1314(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[41:41]),.I2(s_fract_48_i[42:42]),.I3(s_fract_48_i[43:43]),.I4(N_592),.I5(N_1254),.O(N_709));
defparam desc1314.INIT=64'h0000000000000001;
  LUT6 un1_s_overflow_2_cZ(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.I2(s_expo2b[3:3]),.I3(s_expo2b[1:1]),.I4(s_expo2b[6:6]),.I5(un1_s_expo3),.O(un1_s_overflow_2));
defparam un1_s_overflow_2_cZ.INIT=64'h60900000F0000000;
  LUT6_L desc1315(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.I2(s_output_o25_sn),.I3(s_expo2b[1:1]),.I4(s_expo2b[2:2]),.I5(un1_s_expo3),.LO(s_output_o_m0[25:25]));
defparam desc1315.INIT=64'h060F09000F0F0000;
  LUT6 desc1316(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(N_1246),.I5(N_582),.O(N_1328));
defparam desc1316.INIT=64'h00000000000F000E;
  LUT5_L desc1317(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[24:24]),.I3(N_1364),.I4(N_1358),.LO(N_1365));
defparam desc1317.INIT=32'h0F000E00;
  LUT6 desc1318(.I0(s_fract_48_i[47:47]),.I1(s_shr2[2:2]),.I2(s_shr2[3:3]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.I5(N_92),.O(N_286));
defparam desc1318.INIT=64'h0303030B00000008;
  LUT6 desc1319(.I0(s_fract_48_i[47:47]),.I1(s_shr2[2:2]),.I2(s_shr2[3:3]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.I5(s_fract_48_i_RNI21942_O6[46:46]),.O(N_1137));
defparam desc1319.INIT=64'h0003020300000200;
  LUT6 desc1320(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[4:4]),.I3(s_fract_48_i[5:5]),.I4(s_fract_48_i[6:6]),.I5(s_fract_48_i[2:2]),.O(N_1370));
defparam desc1320.INIT=64'h0000000000000001;
  LUT6_L desc1321(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[2:2]),.I2(N_1255),.I3(N_447),.I4(N_530_1),.I5(N_426),.LO(N_1267));
defparam desc1321.INIT=64'hFF00FF00FFFEFFF0;
  LUT6_L desc1322(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[25:25]),.I4(v_count_49_0_o2[4:4]),.I5(N_689),.LO(N_626));
defparam desc1322.INIT=64'hFFCDFFCDFFCDFFCC;
  LUT6_L desc1323(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_73),.I4(N_77),.I5(N_253),.LO(N_404));
defparam desc1323.INIT=64'h0A0208005F575D55;
  LUT6 desc1324(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_73),.I4(N_77),.I5(N_218),.O(N_234));
defparam desc1324.INIT=64'hAFABAEAA05010400;
  LUT6 desc1325(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[5:5]),.I3(s_fract_48_i[6:6]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_260));
defparam desc1325.INIT=64'h00FF33330F0F5555;
  LUT6 desc1326(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[38:38]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_84));
defparam desc1326.INIT=64'hFF00AAAACCCCF0F0;
  LUT6 desc1327(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[18:18]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_66_0));
defparam desc1327.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc1328(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_74),.I4(N_70),.I5(N_360),.O(N_371));
defparam desc1328.INIT=64'hAFAEABAA05040100;
  LUT5 desc1329(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[3:3]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_fract_48_i[47:47]),.O(s_exp_10_i_RNIE6AQ1[2:2]));
defparam desc1329.INIT=32'h6CCCCCCC;
  LUT6 desc1330(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[25:25]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_74_0));
defparam desc1330.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1331(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_72_0));
defparam desc1331.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1332(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_66),.I4(N_70),.I5(N_1140),.O(N_1141));
defparam desc1332.INIT=64'h5F575D550A020800;
  LUT6 desc1333(.I0(s_fract_48_i[0:0]),.I1(s_fract_48_i[1:1]),.I2(s_fract_48_i[2:2]),.I3(s_shl2[1:1]),.I4(s_shl2[0:0]),.I5(s_shl2[2:2]),.O(N_1078));
defparam desc1333.INIT=64'h0000000000CCAAF0;
  LUT6 desc1334(.I0(s_zeros[3:3]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[3:3]),.I3(s_exp_10_i[1:1]),.I4(s_exp_10_i[0:0]),.I5(s_fract_48_i[47:47]),.O(s_exp_10b_axb_3));
defparam desc1334.INIT=64'h69A5A5A5A5A5A5A5;
  LUT6 desc1335(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_80_1));
defparam desc1335.INIT=64'hAAAAF0F0FF00CCCC;
  LUT6 desc1336(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[29:29]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_76_0));
defparam desc1336.INIT=64'hAAAAF0F0FF00CCCC;
  LUT6 desc1337(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[24:24]),.I3(s_fract_48_i[23:23]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_70_0));
defparam desc1337.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6 desc1338(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[16:16]),.I2(s_fract_48_i[15:15]),.I3(s_fract_48_i[18:18]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_64_1));
defparam desc1338.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1339(.I0(s_exp_10_i[4:4]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[3:3]),.I3(s_exp_10_i[1:1]),.I4(s_exp_10_i[0:0]),.I5(s_fract_48_i[47:47]),.O(s_exp_10_i_RNI5I152[2:2]));
defparam desc1339.INIT=64'h6AAAAAAAAAAAAAAA;
  LUT6 desc1340(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[21:21]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_68_0));
defparam desc1340.INIT=64'hAAAACCCCFF00F0F0;
  LUT5 desc1341(.I0(s_fract_48_i[47:47]),.I1(s_shr2[2:2]),.I2(s_shr2[3:3]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.O(N_1090));
defparam desc1341.INIT=32'h00000002;
  LUT6 desc1342(.I0(s_fract_48_i[5:5]),.I1(s_fract_48_i[6:6]),.I2(s_fract_48_i[8:8]),.I3(s_fract_48_i[7:7]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(m40));
defparam desc1342.INIT=64'h0F0F333300FF5555;
  LUT6 desc1343(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_47),.I3(N_1124),.I4(N_56),.I5(N_60),.O(N_304));
defparam desc1343.INIT=64'h2031A8B96475ECFD;
  LUT6 desc1344(.I0(s_fract_48_i[0:0]),.I1(s_fract_48_i[1:1]),.I2(s_shl2[1:1]),.I3(s_shl2[0:0]),.I4(s_shl2[2:2]),.I5(s_shl2[5:5]),.O(N_327));
defparam desc1344.INIT=64'h0000000000000A0C;
  LUT5 desc1345(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_55_0),.I3(N_31_0),.I4(N_87),.O(N_56_0));
defparam desc1345.INIT=32'hD1F3C0E2;
  LUT6 desc1346(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_31_0),.I3(N_83),.I4(N_87),.I5(N_79),.O(N_80_0));
defparam desc1346.INIT=64'h80A2C4E691B3D5F7;
  LUT6_L desc1347(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_63),.I4(N_59),.I5(N_103),.LO(N_77_0));
defparam desc1347.INIT=64'h0F0E0B0A05040100;
  LUT6 desc1348(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_131),.I3(N_1077),.I4(N_63),.I5(N_59),.O(N_1120));
defparam desc1348.INIT=64'h0123456789ABCDEF;
  LUT6 desc1349(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[34:34]),.I3(s_fract_48_i[35:35]),.I4(s_fract_48_i[28:28]),.I5(s_fract_48_i[29:29]),.O(N_1337));
defparam desc1349.INIT=64'h000000000000FFFE;
  LUT6 desc1350(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.I3(s_fract_48_i[11:11]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_60_1));
defparam desc1350.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6 desc1351(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[43:43]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_131));
defparam desc1351.INIT=64'hFF00F0F0AAAACCCC;
  LUT6 desc1352(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[15:15]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_62_0));
defparam desc1352.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc1353(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[4:4]),.I3(s_fract_48_i[2:2]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_322));
defparam desc1353.INIT=64'h0F0F00FF33335555;
  LUT6 desc1354(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[21:21]),.I4(s_fract_48_i[16:16]),.I5(s_fract_48_i[18:18]),.O(v_count_49_i_o3_1[1:1]));
defparam desc1354.INIT=64'hFFFFCCCCFFFFCFCE;
  LUT6_L desc1355(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_61),.I4(N_57),.I5(N_101),.LO(N_206));
defparam desc1355.INIT=64'h0F0E0B0A05040100;
  LUT3 desc1356(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.O(N_1273));
defparam desc1356.INIT=8'hFE;
  LUT5 un7_s_expo3_ac0_5(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.I2(s_expo2b[3:3]),.I3(s_expo2b[1:1]),.I4(s_expo2b[2:2]),.O(un7_s_expo3_c4));
defparam un7_s_expo3_ac0_5.INIT=32'h90000000;
  LUT6_L desc1357(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(s_shr2[3:3]),.I3(N_139),.I4(N_194),.I5(N_192),.LO(s_frac2a_3[10:10]));
defparam desc1357.INIT=64'h1311575502004644;
  LUT6 desc1358(.I0(s_infb),.I1(un1_s_infa),.I2(result_5),.I3(un1_s_nan_b),.I4(result_4),.I5(un1_s_nan_a),.O(s_output_o_sn_N_5_mux));
defparam desc1358.INIT=64'h0000000000F10011;
  LUT6 un1_s_overflow_0_cZ(.I0(s_expo2b[0:0]),.I1(s_infb),.I2(un1_s_infa),.I3(s_expo2b[2:2]),.I4(s_expo3[7:7]),.I5(un1_s_expo3),.O(un1_s_overflow_0));
defparam un1_s_overflow_0_cZ.INIT=64'h0100000002000000;
  LUT6_L desc1359(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_25_0),.I4(N_1084),.I5(N_1129),.LO(N_1131));
defparam desc1359.INIT=64'hA0802000F0D07050;
  LUT6_L desc1360(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(s_shr2[3:3]),.I3(N_138),.I4(N_354),.I5(N_355),.LO(s_frac2a_3[9:9]));
defparam desc1360.INIT=64'h5755464413110200;
  LUT6 desc1361(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_36),.I3(N_12_0),.I4(N_16_0),.I5(N_20_0),.O(s_frac2a_1_134));
defparam desc1361.INIT=64'h1054327698DCBAFE;
  LUT6 desc1362(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[34:34]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[32:32]),.I4(N_1259),.I5(N_1252),.O(N_1277));
defparam desc1362.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L un1_s_ine_o_cZ(.I0(s_expo2b[4:4]),.I1(s_expo2b[5:5]),.I2(un3_s_ine_o),.I3(un3_s_op_0),.I4(un1_s_overflow_0),.I5(un1_s_overflow_2),.LO(un1_s_ine_o));
defparam un1_s_ine_o_cZ.INIT=64'hF800F000F000F000;
  LUT6 s_output_os2_1(.I0(s_infb),.I1(un1_s_infa),.I2(s_expo2b[4:4]),.I3(s_expo2b[5:5]),.I4(un1_s_overflow_0),.I5(un1_s_overflow_2),.O(s_output_o_sm0));
defparam s_output_os2_1.INIT=64'hFEEEEEEEEEEEEEEE;
  LUT6_L desc1363(.I0(s_fract_48_i[5:5]),.I1(s_fract_48_i[6:6]),.I2(N_1253),.I3(N_434_i_0),.I4(N_530_1),.I5(N_449),.LO(N_535));
defparam desc1363.INIT=64'h0F000F0001000000;
  LUT5 desc1364(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[16:16]),.I4(s_fract_48_i[18:18]),.O(N_443));
defparam desc1364.INIT=32'h50505455;
  LUT1 s_frac_rnd_3_0_axb_24_cZ(.I0(s_frac2a[47:47]),.O(s_frac_rnd_3_0_axb_24));
defparam s_frac_rnd_3_0_axb_24_cZ.INIT=2'h2;
  LUT2 s_expo2b_axb_7_cZ(.I0(s_expo1[7:7]),.I1(s_frac2a[46:46]),.O(s_expo2b_axb_7));
defparam s_expo2b_axb_7_cZ.INIT=4'h9;
  LUT2 s_expo2b_axb_0(.I0(s_expo1[0:0]),.I1(s_frac2a[46:46]),.O(s_expo2b[0:0]));
defparam s_expo2b_axb_0.INIT=4'h9;
  LUT2 desc1365(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[41:41]),.O(v_count_49_0_o2_9[4:4]));
defparam desc1365.INIT=4'hE;
  LUT2 desc1366(.I0(s_fract_48_i[28:28]),.I1(s_fract_48_i[29:29]),.O(v_count_49_0_o2[4:4]));
defparam desc1366.INIT=4'hE;
  LUT2 desc1367(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.O(v_count_49_0_o2_6[4:4]));
defparam desc1367.INIT=4'hE;
  LUT2 desc1368(.I0(s_fracta_i_20),.I1(s_fracta_i_21),.O(result_11));
defparam desc1368.INIT=4'hE;
  LUT3 desc1369(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[29:29]),.I2(s_shr2[0:0]),.O(N_30));
defparam desc1369.INIT=8'hAC;
  LUT3 desc1370(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[33:33]),.I2(s_shr2[0:0]),.O(N_273));
defparam desc1370.INIT=8'hAC;
  LUT3 desc1371(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[43:43]),.I2(s_shl2[0:0]),.O(N_279));
defparam desc1371.INIT=8'hCA;
  LUT3 desc1372(.I0(s_fract_48_i[37:37]),.I1(s_fract_48_i[38:38]),.I2(s_shr2[0:0]),.O(N_12_0));
defparam desc1372.INIT=8'h35;
  LUT3 desc1373(.I0(s_fract_48_i[23:23]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.O(N_1364));
defparam desc1373.INIT=8'h01;
  LUT4 desc1374(.I0(s_fract_48_i[0:0]),.I1(s_fract_48_i[1:1]),.I2(s_shl2[1:1]),.I3(s_shl2[0:0]),.O(N_50));
defparam desc1374.INIT=16'h0A0C;
  LUT5 un4_s_exp_10b_0_2_cZ(.I0(s_exp_10b_i),.I1(s_exp_10b[1:1]),.I2(s_exp_10b[2:2]),.I3(s_exp_10b[3:3]),.I4(s_exp_10b[4:4]),.O(un4_s_exp_10b_0_2));
defparam un4_s_exp_10b_0_2_cZ.INIT=32'h00000002;
  LUT6 un3_s_ine_o_0_0_cZ(.I0(s_frac2a[0:0]),.I1(s_frac2a[1:1]),.I2(s_frac2a[16:16]),.I3(s_frac2a[17:17]),.I4(s_frac2a[18:18]),.I5(s_frac2a[19:19]),.O(un3_s_ine_o_0_0));
defparam un3_s_ine_o_0_0_cZ.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 un3_s_ine_o_0_1_cZ(.I0(s_frac2a[2:2]),.I1(s_frac2a[3:3]),.I2(s_frac2a[4:4]),.I3(s_frac2a[5:5]),.I4(s_frac2a[6:6]),.I5(s_frac2a[7:7]),.O(un3_s_ine_o_0_1));
defparam un3_s_ine_o_0_1_cZ.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 un3_s_ine_o_0_2_cZ(.I0(s_frac2a[8:8]),.I1(s_frac2a[9:9]),.I2(s_frac2a[10:10]),.I3(s_frac2a[11:11]),.I4(s_frac2a[12:12]),.I5(s_frac2a[13:13]),.O(un3_s_ine_o_0_2));
defparam un3_s_ine_o_0_2_cZ.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc1375(.I0(s_fracta_i_0),.I1(s_fracta_i_1),.I2(s_fracta_i_2),.I3(s_fracta_i_3),.I4(s_fracta_i_4),.I5(s_fracta_i_5),.O(result_3_21_1));
defparam desc1375.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc1376(.I0(s_fracta_i_6),.I1(s_fracta_i_7),.I2(s_fracta_i_8),.I3(s_fracta_i_9),.I4(s_fracta_i_10),.I5(s_fracta_i_11),.LO(result_3_21_0));
defparam desc1376.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc1377(.I0(s_fract_48_i[0:0]),.I1(s_fract_48_i[1:1]),.I2(s_fract_48_i[3:3]),.I3(s_fract_48_i[2:2]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_49_0));
defparam desc1377.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc1378(.I0(s_fract_48_i[0:0]),.I1(s_fract_48_i[1:1]),.I2(s_fract_48_i[3:3]),.I3(s_fract_48_i[2:2]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_52));
defparam desc1378.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1379(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[4:4]),.I3(s_fract_48_i[2:2]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_53));
defparam desc1379.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1380(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[5:5]),.I3(s_fract_48_i[2:2]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_51));
defparam desc1380.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1381(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[5:5]),.I3(s_fract_48_i[2:2]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_54));
defparam desc1381.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1382(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[5:5]),.I3(s_fract_48_i[6:6]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_55_1));
defparam desc1382.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1383(.I0(s_fract_48_i[4:4]),.I1(s_fract_48_i[5:5]),.I2(s_fract_48_i[6:6]),.I3(s_fract_48_i[7:7]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_53_0));
defparam desc1383.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc1384(.I0(s_fract_48_i[4:4]),.I1(s_fract_48_i[5:5]),.I2(s_fract_48_i[6:6]),.I3(s_fract_48_i[7:7]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_56));
defparam desc1384.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1385(.I0(s_fract_48_i[5:5]),.I1(s_fract_48_i[6:6]),.I2(s_fract_48_i[8:8]),.I3(s_fract_48_i[7:7]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_57));
defparam desc1385.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1386(.I0(s_fract_48_i[6:6]),.I1(s_fract_48_i[8:8]),.I2(s_fract_48_i[9:9]),.I3(s_fract_48_i[7:7]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_55));
defparam desc1386.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc1387(.I0(s_fract_48_i[6:6]),.I1(s_fract_48_i[8:8]),.I2(s_fract_48_i[9:9]),.I3(s_fract_48_i[7:7]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_58));
defparam desc1387.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1388(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[7:7]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_59));
defparam desc1388.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1389(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(s_frac2a_1_58));
defparam desc1389.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc1390(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_60));
defparam desc1390.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1391(.I0(s_fract_48_i[12:12]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_58_0));
defparam desc1391.INIT=64'hAAAAF0F0FF00CCCC;
  LUT6 desc1392(.I0(s_fract_48_i[12:12]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_61));
defparam desc1392.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1393(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[12:12]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_59_0));
defparam desc1393.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1394(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[12:12]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_62));
defparam desc1394.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc1395(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.I3(s_fract_48_i[11:11]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_63));
defparam desc1395.INIT=64'hFF00AAAAF0F0CCCC;
  LUT6 desc1396(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.I3(s_fract_48_i[15:15]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(s_frac2a_1_62));
defparam desc1396.INIT=64'hFF00AAAACCCCF0F0;
  LUT6 desc1397(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.I3(s_fract_48_i[15:15]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_64));
defparam desc1397.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc1398(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[15:15]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_65));
defparam desc1398.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1399(.I0(s_fract_48_i[14:14]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[15:15]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_66));
defparam desc1399.INIT=64'hAAAAF0F0FF00CCCC;
  LUT6 desc1400(.I0(s_fract_48_i[14:14]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[15:15]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_63_0));
defparam desc1400.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1401(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[16:16]),.I2(s_fract_48_i[15:15]),.I3(s_fract_48_i[18:18]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_67));
defparam desc1401.INIT=64'hF0F0AAAACCCCFF00;
  LUT6 desc1402(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_68));
defparam desc1402.INIT=64'hF0F0FF00AAAACCCC;
  LUT6 desc1403(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_65_0));
defparam desc1403.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc1404(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[18:18]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_69));
defparam desc1404.INIT=64'hCCCCF0F0FF00AAAA;
  LUT6 desc1405(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[18:18]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_70));
defparam desc1405.INIT=64'hFF00AAAACCCCF0F0;
  LUT6 desc1406(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[18:18]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_67_0));
defparam desc1406.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc1407(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[19:19]),.I3(s_fract_48_i[21:21]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_71));
defparam desc1407.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc1408(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[23:23]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_72));
defparam desc1408.INIT=64'hCCCCAAAAF0F0FF00;
  LUT6 desc1409(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[23:23]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_69_1));
defparam desc1409.INIT=64'hFF00F0F0AAAACCCC;
  LUT6 desc1410(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[24:24]),.I3(s_fract_48_i[23:23]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_73));
defparam desc1410.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6 desc1411(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_74));
defparam desc1411.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc1412(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_71_0));
defparam desc1412.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc1413(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_75_0));
defparam desc1413.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc1414(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[25:25]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_76));
defparam desc1414.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc1415(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[34:34]),.I3(s_fract_48_i[35:35]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_86));
defparam desc1415.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6 desc1416(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[35:35]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_84_0));
defparam desc1416.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6 desc1417(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[38:38]),.I2(s_fract_48_i[39:39]),.I3(s_fract_48_i[41:41]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_49));
defparam desc1417.INIT=64'h333355550F0F00FF;
  LUT6 desc1418(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[39:39]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_47));
defparam desc1418.INIT=64'h55550F0F333300FF;
  LUT6 desc1419(.I0(s_fract_48_i[37:37]),.I1(s_fract_48_i[40:40]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[39:39]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(s_frac2a_2_91));
defparam desc1419.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc1420(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[7:7]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_60_0_0));
defparam desc1420.INIT=64'h0F0F5555333300FF;
  LUT6 desc1421(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[35:35]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_81_0));
defparam desc1421.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6 desc1422(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_82));
defparam desc1422.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1423(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[28:28]),.I2(s_fract_48_i[29:29]),.I3(s_fract_48_i[31:31]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_80));
defparam desc1423.INIT=64'hCCCCAAAAF0F0FF00;
  LUT6 desc1424(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[29:29]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_79_1));
defparam desc1424.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1425(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[29:29]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_78));
defparam desc1425.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1426(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[25:25]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_77));
defparam desc1426.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1427(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[47:47]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_905));
defparam desc1427.INIT=64'h00FF0F0F33335555;
  LUT6 desc1428(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[45:45]),.I2(s_fract_48_i[42:42]),.I3(s_fract_48_i[43:43]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_31_0));
defparam desc1428.INIT=64'h333300FF55550F0F;
  LUT6 desc1429(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[41:41]),.I2(s_fract_48_i[42:42]),.I3(s_fract_48_i[43:43]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_904));
defparam desc1429.INIT=64'h00FF33330F0F5555;
  LUT6 desc1430(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[38:38]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_87_0));
defparam desc1430.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc1431(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[34:34]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[33:33]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_85_0));
defparam desc1431.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc1432(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_83_0));
defparam desc1432.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1433(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[29:29]),.I2(s_fract_48_i[31:31]),.I3(s_fract_48_i[32:32]),.I4(s_shl2[1:1]),.I5(s_shl2[0:0]),.O(N_81));
defparam desc1433.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6 desc1434(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_79));
defparam desc1434.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc1435(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[28:28]),.I2(s_fract_48_i[29:29]),.I3(s_fract_48_i[31:31]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_77_1));
defparam desc1435.INIT=64'hFF00F0F0AAAACCCC;
  LUT6 desc1436(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[28:28]),.I3(s_fract_48_i[29:29]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_75));
defparam desc1436.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc1437(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[25:25]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_73_0));
defparam desc1437.INIT=64'hF0F0FF00AAAACCCC;
  LUT6 desc1438(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[38:38]),.I2(s_fract_48_i[39:39]),.I3(s_fract_48_i[41:41]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_87));
defparam desc1438.INIT=64'hFF00F0F0AAAACCCC;
  LUT6 desc1439(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[39:39]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_85));
defparam desc1439.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6 desc1440(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[34:34]),.I3(s_fract_48_i[35:35]),.I4(s_shr2[1:1]),.I5(s_shr2[0:0]),.O(N_83));
defparam desc1440.INIT=64'hCCCCFF00AAAAF0F0;
  LUT6_L un5_s_exp_10a_1_cZ(.I0(s_zeros_RNI0TNS_O5),.I1(un5_v_shr1_axb1),.I2(s_exp_10_i_RNIORIF1[2:2]),.I3(s_exp_10_i_RNIE6AQ1[2:2]),.I4(s_exp_10_i_RNI5I152[2:2]),.I5(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91),.LO(un5_s_exp_10a_1));
defparam un5_s_exp_10a_1_cZ.INIT=64'h0000000000000001;
  LUT6 desc1441(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[40:40]),.I2(s_fract_48_i[46:46]),.I3(s_fract_48_i[45:45]),.I4(s_fract_48_i[42:42]),.I5(v_count_49_0_o2_6[4:4]),.O(v_count_0_sqmuxa_47_0));
defparam desc1441.INIT=64'h0000000000000001;
  LUT5 desc1442(.I0(s_fracta_i_12),.I1(s_fracta_i_13),.I2(s_fracta_i_14),.I3(s_fracta_i_15),.I4(result_3_21_0),.O(result_3_21_3));
defparam desc1442.INIT=32'hFFFFFFFE;
  LUT5_L un2_s_lost_axbxc3_cZ(.I0(s_frac_rnd[24:24]),.I1(s_shr2[2:2]),.I2(s_shr2[3:3]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.LO(un2_s_lost_axbxc3));
defparam un2_s_lost_axbxc3_cZ.INIT=32'h78F0F0F0;
  LUT5 un2_s_exp_10a_ac0_5(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[3:3]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_fract_48_i[47:47]),.O(un2_s_exp_10a_c4));
defparam un2_s_exp_10a_ac0_5.INIT=32'h80000000;
  LUT5 desc1443(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[28:28]),.I4(s_fract_48_i[25:25]),.O(N_1305));
defparam desc1443.INIT=32'hFF0AFF0E;
  LUT5 desc1444(.I0(s_fract_48_i[0:0]),.I1(s_shl2[1:1]),.I2(s_shl2[0:0]),.I3(s_shl2[3:3]),.I4(s_shl2[2:2]),.O(N_318));
defparam desc1444.INIT=32'h00000002;
  LUT6 desc1445(.I0(s_fract_48_i[0:0]),.I1(s_shl2[1:1]),.I2(s_shl2[0:0]),.I3(s_shl2[2:2]),.I4(N_3),.I5(N_55_1),.O(N_103));
defparam desc1445.INIT=64'h3BFF08FF3B000800;
  LUT5 desc1446(.I0(s_fract_48_i[0:0]),.I1(s_shl2[1:1]),.I2(s_shl2[0:0]),.I3(s_shl2[2:2]),.I4(N_53),.O(N_101));
defparam desc1446.INIT=32'h02FF0200;
  LUT6 desc1447(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_903),.I3(N_35_0),.I4(s_fract_48_i_RNI21942_O6[46:46]),.I5(N_20_0),.O(N_138));
defparam desc1447.INIT=64'hAE268C04BF379D15;
  LUT6 desc1448(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[47:47]),.I2(s_shr2[2:2]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.I5(N_31_0),.O(N_139));
defparam desc1448.INIT=64'h00C000A00FCF0FAF;
  LUT5 desc1449(.I0(s_shl2[1:1]),.I1(s_shl2[2:2]),.I2(N_279),.I3(N_1288),.I4(s_frac2a_2_91),.O(N_250));
defparam desc1449.INIT=32'h0123CDEF;
  LUT5 desc1450(.I0(s_shl2[1:1]),.I1(s_shl2[2:2]),.I2(N_1289),.I3(N_1076),.I4(N_49),.O(N_1150));
defparam desc1450.INIT=32'hCEDF0213;
  LUT5 desc1451(.I0(s_shl2[1:1]),.I1(s_shl2[2:2]),.I2(N_269),.I3(N_1076),.I4(N_1124),.O(N_1125));
defparam desc1451.INIT=32'hFEDC3210;
  LUT3 desc1452(.I0(s_shl2[2:2]),.I1(N_56),.I2(N_60),.O(s_frac2a_2_111));
defparam desc1452.INIT=8'hD8;
  LUT3_L desc1453(.I0(s_shl2[2:2]),.I1(N_53),.I2(N_57),.LO(N_105));
defparam desc1453.INIT=8'hD8;
  LUT6 desc1454(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_903),.I3(N_12_0),.I4(N_16_0),.I5(N_20_0),.O(N_134));
defparam desc1454.INIT=64'h08194C5D2A3B6E7F;
  LUT6 desc1455(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_273),.I3(N_36),.I4(N_12_0),.I5(N_16_0),.O(s_frac2a_1_132));
defparam desc1455.INIT=64'h54107632DC98FEBA;
  LUT6 desc1456(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_30),.I3(N_273),.I4(N_40),.I5(N_36),.O(N_126));
defparam desc1456.INIT=64'hBA98FEDC32107654;
  LUT5 desc1457(.I0(s_shr2[2:2]),.I1(s_shr2[1:1]),.I2(N_30),.I3(N_40),.I4(N_74_0),.O(s_frac2a_1_124));
defparam desc1457.INIT=32'h75FD20A8;
  LUT3 desc1458(.I0(s_shr2[2:2]),.I1(N_59_0),.I2(N_63_0),.O(s_frac2a_1_109));
defparam desc1458.INIT=8'hE4;
  LUT6 desc1459(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[34:34]),.I2(N_1367),.I3(N_1252),.I4(N_1260),.I5(N_1353),.O(N_23_0_2));
defparam desc1459.INIT=64'h00FCAAFE00000000;
  LUT6_L desc1460(.I0(s_fract_48_i[35:35]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[47:47]),.I3(N_320_2),.I4(v_count_0_sqmuxa_47_1_4),.I5(v_count_0_sqmuxa_47_2_4),.LO(v_count_0_sqmuxa_47_1_0));
defparam desc1460.INIT=64'h0100000000000000;
  LUT6_L desc1461(.I0(N_592),.I1(v_count_49_0_o2_9[4:4]),.I2(N_591),.I3(s_zeros_2_0_i_a2_3_lut6_2_O5),.I4(v_count_49_0_o2_6[4:4]),.I5(N_1254),.LO(N_693));
defparam desc1461.INIT=64'h00000F0C00000F0D;
  LUT5 un4_s_lost_c2_cZ(.I0(s_r_zeros[0:0]),.I1(s_r_zeros[1:1]),.I2(s_frac_rnd[24:24]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.O(un4_s_lost_c2));
defparam un4_s_lost_c2_cZ.INIT=32'h07317310;
  LUT6 desc1462(.I0(s_fract_48_i[11:11]),.I1(s_fract_48_i[15:15]),.I2(N_1273),.I3(N_449),.I4(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I5(N_1251),.O(N_247));
defparam desc1462.INIT=64'hFFFFFFFFFFFFCCCD;
  LUT6_L desc1463(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[4:4]),.I3(s_fract_48_i[5:5]),.I4(s_fract_48_i[6:6]),.I5(s_fract_48_i[2:2]),.LO(N_1264));
defparam desc1463.INIT=64'hFFFF00F3FFFF00F1;
  LUT6_L desc1464(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[42:42]),.I4(s_fract_48_i[43:43]),.I5(s_fract_48_i[47:47]),.LO(N_686));
defparam desc1464.INIT=64'h00FF005100FF0050;
  LUT4 desc1465(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_66),.I3(N_70),.O(N_1093));
defparam desc1465.INIT=16'h3120;
  LUT6 desc1466(.I0(s_fract_48_i[9:9]),.I1(s_fract_48_i[31:31]),.I2(N_663_3),.I3(N_426),.I4(N_1273),.I5(N_1370),.O(v_count_0_sqmuxa_46_0));
defparam desc1466.INIT=64'h0000001000000000;
  LUT6_L desc1467(.I0(s_fract_48_i[23:23]),.I1(N_614),.I2(v_count_49_0_o2_6[4:4]),.I3(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I4(N_1251),.I5(N_331_0_4),.LO(N_331_0));
defparam desc1467.INIT=64'h0000000100000000;
  LUT6 desc1468(.I0(N_588),.I1(N_331_1),.I2(N_239),.I3(N_1308),.I4(N_1337),.I5(v_count_49_i_o3_i_a2_lut6_2_O5[3:3]),.O(N_669_0));
defparam desc1468.INIT=64'h0000000400000000;
  LUT6 desc1469(.I0(s_fract_48_i[6:6]),.I1(s_fract_48_i[8:8]),.I2(s_fract_48_i[9:9]),.I3(s_fract_48_i[7:7]),.I4(N_704),.I5(N_1308),.O(N_662));
defparam desc1469.INIT=64'h0000000000550054;
  LUT6 desc1470(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[7:7]),.I3(s_fract_48_i[2:2]),.I4(v_count_49_i_o3_i_a2_lut6_2_O6[3:3]),.I5(N_708),.O(N_650));
defparam desc1470.INIT=64'h00FF000000F40000;
  LUT5 un3_s_ine_o_0_3(.I0(s_frac2a[14:14]),.I1(s_frac2a[15:15]),.I2(un3_s_ine_o_0_0),.I3(un3_s_ine_o_0_1),.I4(un3_s_ine_o_0_2),.O(un3_s_ine_o_0));
defparam un3_s_ine_o_0_3.INIT=32'hFFFFFFFE;
  LUT6 desc1471(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_260),.I3(N_60_0_0),.I4(N_60_1),.I5(N_64_1),.O(N_263));
defparam desc1471.INIT=64'h32107654BA98FEDC;
  LUT6 desc1472(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(N_53),.I3(N_65),.I4(N_61),.I5(N_57),.O(N_161_0));
defparam desc1472.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc1473(.I0(s_fract_48_i[0:0]),.I1(s_shl2[1:1]),.I2(s_shl2[0:0]),.I3(s_shl2[3:3]),.I4(s_shl2[2:2]),.I5(N_105),.O(N_153));
defparam desc1473.INIT=64'h00FF02FF00000200;
  LUT6 desc1474(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_85),.I3(N_77_1),.I4(N_81_0),.I5(N_73_0),.O(N_169));
defparam desc1474.INIT=64'hF7D5B391E6C4A280;
  LUT6 desc1475(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_frac2a_1_58),.I3(s_frac2a_1_62),.I4(N_69_1),.I5(N_65_0),.O(N_423));
defparam desc1475.INIT=64'h012389AB4567CDEF;
  LUT5 desc1476(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_50),.I3(N_82),.I4(N_78),.O(N_1154));
defparam desc1476.INIT=32'h8C9DAEBF;
  LUT6 desc1477(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_905),.I3(N_85),.I4(N_904),.I5(N_81_0),.O(N_382));
defparam desc1477.INIT=64'hC4E680A2D5F791B3;
  LUT6 desc1478(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_58_0),.I3(N_62_0),.I4(N_70_0),.I5(N_66_0),.O(N_349));
defparam desc1478.INIT=64'hFEDC7654BA983210;
  LUT6 desc1479(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_53_0),.I3(s_frac2a_1_58),.I4(s_frac2a_1_62),.I5(N_65_0),.O(N_342));
defparam desc1479.INIT=64'h0123456789ABCDEF;
  LUT5 desc1480(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_70_0),.I3(N_66_0),.I4(s_frac2a_1_124),.O(N_333));
defparam desc1480.INIT=32'hFDEC3120;
  LUT6_L desc1481(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_322),.I3(m40),.I4(N_58_0),.I5(N_62_0),.LO(N_325));
defparam desc1481.INIT=64'hCDEF89AB45670123;
  LUT5 desc1482(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_80),.I3(N_84_0),.I4(N_52),.O(N_296));
defparam desc1482.INIT=32'h8A9BCEDF;
  LUT5 desc1483(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_76_0),.I3(N_80_1),.I4(s_frac2a_1_134),.O(N_284));
defparam desc1483.INIT=32'h0123CDEF;
  LUT6 desc1484(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_60_1),.I3(N_68_0),.I4(N_64_1),.I5(N_72_0),.O(N_278));
defparam desc1484.INIT=64'h0145236789CDABEF;
  LUT6 desc1485(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(N_35_0),.I4(N_92),.I5(s_frac2a_1_134),.O(N_275));
defparam desc1485.INIT=64'h8088C4CCB3BBF7FF;
  LUT6 desc1486(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_68_0),.I3(N_76_0),.I4(N_80_1),.I5(N_72_0),.O(N_271));
defparam desc1486.INIT=64'h014589CD2367ABEF;
  LUT5 desc1487(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_85_0),.I3(N_81),.I4(N_101),.O(N_253));
defparam desc1487.INIT=32'h0123CDEF;
  LUT5 desc1488(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_83_0),.I3(N_79_1),.I4(N_1078),.O(N_242));
defparam desc1488.INIT=32'hFEDC3210;
  LUT6 desc1489(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_87_0),.I3(N_1077),.I4(N_55_1),.I5(N_59),.O(N_240));
defparam desc1489.INIT=64'h02138A9B4657CEDF;
  LUT6 desc1490(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_69_1),.I3(N_77_1),.I4(N_81_0),.I5(N_73_0),.O(N_217));
defparam desc1490.INIT=64'h014589CD2367ABEF;
  LUT6 desc1491(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_85),.I3(N_904),.I4(N_77_1),.I5(N_81_0),.O(N_211));
defparam desc1491.INIT=64'h8C049D15AE26BF37;
  LUT6 desc1492(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_frac2a_1_62),.I3(N_69_1),.I4(N_65_0),.I5(N_73_0),.O(N_201));
defparam desc1492.INIT=64'h0145236789CDABEF;
  LUT6 desc1493(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_83),.I3(N_87),.I4(N_79),.I5(N_75),.O(N_194));
defparam desc1493.INIT=64'h048C26AE159D37BF;
  LUT6 desc1494(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_50),.I3(N_86),.I4(N_82),.I5(N_54),.O(N_1152));
defparam desc1494.INIT=64'h08192A3B4C5D6E7F;
  LUT6 desc1495(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_47),.I3(N_84_0),.I4(N_52),.I5(N_56),.O(N_1128));
defparam desc1495.INIT=64'h103298BA5476DCFE;
  LUT5 desc1496(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_87_0),.I3(N_83_0),.I4(N_103),.O(N_1114));
defparam desc1496.INIT=32'h0123CDEF;
  LUT6 desc1497(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_68_0),.I3(N_76_0),.I4(N_64_1),.I5(N_72_0),.O(N_85_0_0));
defparam desc1497.INIT=64'h028A139B46CE57DF;
  LUT6 desc1498(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_63_0),.I3(N_71_0),.I4(N_67_0),.I5(N_75),.O(N_74_0_0));
defparam desc1498.INIT=64'h0145236789CDABEF;
  LUT6 desc1499(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(N_35_0),.I4(N_88),.I5(N_92),.O(N_71_0_0));
defparam desc1499.INIT=64'h3733262215110400;
  LUT6 desc1500(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_84),.I3(N_76_0),.I4(N_80_1),.I5(N_72_0),.O(N_69_0));
defparam desc1500.INIT=64'h082A4C6E193B5D7F;
  LUT6 desc1501(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_60_0_0),.I3(N_60_1),.I4(N_68_0),.I5(N_64_1),.O(N_64_0_0));
defparam desc1501.INIT=64'h103298BA5476DCFE;
  LUT6 desc1502(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_83),.I3(N_71_0),.I4(N_79),.I5(N_75),.O(N_52_0));
defparam desc1502.INIT=64'h08194C5D2A3B6E7F;
  LUT6 desc1503(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_59_0),.I3(N_55),.I4(N_63_0),.I5(N_67_0),.O(N_44_1));
defparam desc1503.INIT=64'h021346578A9BCEDF;
  LUT6 desc1504(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_84),.I3(N_88),.I4(N_92),.I5(N_80_1),.O(N_1083));
defparam desc1504.INIT=64'h02468ACE13579BDF;
  LUT5 desc1505(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_83),.I3(N_87),.I4(N_139),.O(s_frac2a_1_141_RNIA10R));
defparam desc1505.INIT=32'h0123CDEF;
  LUT6 desc1506(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_69_1),.I3(N_77_1),.I4(N_65_0),.I5(N_73_0),.O(N_161));
defparam desc1506.INIT=64'hFD75EC64B931A820;
  LUT6 desc1507(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(N_35_0),.I4(s_fract_48_i_RNI21942_O6[46:46]),.I5(N_134),.O(N_64_0));
defparam desc1507.INIT=64'h88C88CCCBBFBBFFF;
  LUT5 desc1508(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_74_0),.I3(N_70_0),.I4(N_126),.O(N_60_0));
defparam desc1508.INIT=32'h0213CEDF;
  LUT6 desc1509(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(m40),.I3(N_58_0),.I4(N_62_0),.I5(N_66_0),.O(N_938));
defparam desc1509.INIT=64'h1032547698BADCFE;
  LUT6_L desc1510(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_49_0),.I3(N_53_0),.I4(s_frac2a_1_58),.I5(s_frac2a_1_62),.LO(N_7_0));
defparam desc1510.INIT=64'h0123456789ABCDEF;
  LUT6 desc1511(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_74_0),.I3(N_62_0),.I4(N_70_0),.I5(N_66_0),.O(N_158));
defparam desc1511.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc1512(.I0(N_505_1_2),.I1(N_446),.I2(N_1371),.I3(N_173),.I4(N_301),.I5(N_543),.O(s_zeros_2_2[2:2]));
defparam desc1512.INIT=64'h0000CECC00000000;
  LUT5_L desc1513(.I0(s_fract_48_i[15:15]),.I1(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I2(N_1251),.I3(v_count_0_sqmuxa_46_0),.I4(N_1372),.LO(v_count_0_sqmuxa_46));
defparam desc1513.INIT=32'h01000000;
  LUT6 desc1514(.I0(s_fract_48_i[23:23]),.I1(v_count_49_0_o2[4:4]),.I2(N_610),.I3(s_zeros_2_0_i_a2_1_2_lut6_2_O5),.I4(N_1251),.I5(N_611),.O(N_1281_2));
defparam desc1514.INIT=64'hF0F0F0F5F0F0F0F4;
  LUT6_L desc1515(.I0(v_count_49_0_o2_9[4:4]),.I1(N_614),.I2(N_591),.I3(s_zeros_2_0_i_a2_3_lut6_2_O5),.I4(N_599),.I5(v_count_49_0_o2_6[4:4]),.LO(N_687));
defparam desc1515.INIT=64'h3333333302030202;
  LUT6 un1_s_exp_10a_3_1_cZ(.I0(s_exp_10b[5:5]),.I1(s_exp_10b[6:6]),.I2(un4_s_exp_10b_0_2),.I3(s_exp_10b[7:7]),.I4(s_exp_10b[9:9]),.I5(s_exp_10b[8:8]),.O(un1_s_exp_10a_3_1));
defparam un1_s_exp_10a_3_1_cZ.INIT=64'hFFFF0000FFFF0010;
  LUT6 desc1516(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_65),.I4(N_61),.I5(N_121),.O(N_1167));
defparam desc1516.INIT=64'h0F0D07050A080200;
  LUT6 desc1517(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_55_1),.I4(N_59),.I5(N_115),.O(N_368));
defparam desc1517.INIT=64'h0F070D050A020800;
  LUT6 desc1518(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_71),.I4(N_75_0),.I5(N_115),.O(N_228));
defparam desc1518.INIT=64'h0F0B0E0A05010400;
  LUT6 desc1519(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_1078),.I4(N_55_1),.I5(N_59),.O(N_190));
defparam desc1519.INIT=64'h0F050B010E040A00;
  LUT6 desc1520(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_79_1),.I4(N_75_0),.I5(N_1102),.O(N_116));
defparam desc1520.INIT=64'hAFAEABAA05040100;
  LUT5_L desc1521(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_318),.I3(N_129),.I4(N_121),.LO(i40_mux));
defparam desc1521.INIT=32'hF3E2D1C0;
  LUT5_L desc1522(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_1157),.I3(N_1154),.I4(N_106),.LO(N_1158));
defparam desc1522.INIT=32'hBA10FE54;
  LUT6 desc1523(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_71),.I4(N_75_0),.I5(N_242),.O(N_399));
defparam desc1523.INIT=64'h5F575D550A020800;
  LUT5_L desc1524(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_250),.I3(N_109),.I4(N_253),.LO(N_254));
defparam desc1524.INIT=32'hBAFE1054;
  LUT5_L desc1525(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_1150),.I3(N_110),.I4(N_1152),.LO(N_1153));
defparam desc1525.INIT=32'hBAFE1054;
  LUT5_L desc1526(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_1125),.I3(s_frac2a_2_115_lut6_2_O6),.I4(N_1128),.LO(N_1129));
defparam desc1526.INIT=32'hABEF0145;
  LUT6_L desc1527(.I0(s_shl2[3:3]),.I1(s_shl2[2:2]),.I2(s_shl2[5:5]),.I3(N_79_1),.I4(N_75_0),.I5(N_1114),.LO(N_1115));
defparam desc1527.INIT=64'h0A0802005F5D5755;
  LUT5_L desc1528(.I0(s_shl2[4:4]),.I1(s_shl2[5:5]),.I2(N_318),.I3(un1_s_shr2_1_4),.I4(N_7_0),.LO(N_921));
defparam desc1528.INIT=32'h100010FF;
  LUT5_L desc1529(.I0(s_shr2[4:4]),.I1(s_shr2[3:3]),.I2(N_99),.I3(s_frac2a_1_109),.I4(N_977),.LO(N_195));
defparam desc1529.INIT=32'h5410FEBA;
  LUT5 desc1530(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[19:19]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.I4(N_679),.O(v_count_49_1_3));
defparam desc1530.INIT=32'h0A0E0000;
  LUT6_L desc1531(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[23:23]),.I3(N_239),.I4(N_443),.I5(N_1261),.LO(N_1340));
defparam desc1531.INIT=64'h0000000000F500F4;
  LUT5 un2_s_exp_10a_ac0_1_lut6_2_RNI37EH3(.I0(s_zeros[3:3]),.I1(s_zeros[2:2]),.I2(s_exp_10_i_RNIORIF1[2:2]),.I3(v_shl1_5_0_0_c2),.I4(s_exp_10_i_RNIE6AQ1[2:2]),.O(v_shl1_5_0_0_c4));
defparam un2_s_exp_10a_ac0_1_lut6_2_RNI37EH3.INIT=32'h8A08EFAE;
  LUT6 un2_s_exp_10a_ac0_13(.I0(s_exp_10_i[7:7]),.I1(s_exp_10_i[6:6]),.I2(s_exp_10_i[5:5]),.I3(s_exp_10_i[4:4]),.I4(s_exp_10_i[3:3]),.I5(un2_s_exp_10a_c3),.O(un2_s_exp_10a_c8));
defparam un2_s_exp_10a_ac0_13.INIT=64'h8000000000000000;
  LUT5 desc1532(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.I4(N_679),.O(N_688));
defparam desc1532.INIT=32'h00010000;
  LUT5 desc1533(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.I4(N_679),.O(N_658));
defparam desc1533.INIT=32'h00040000;
  LUT5 desc1534(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_327),.I3(un1_s_shr2_1_4),.I4(N_325),.O(N_330));
defparam desc1534.INIT=32'h10FF1000;
  LUT6_L desc1535(.I0(s_zeros[3:3]),.I1(s_zeros[2:2]),.I2(s_exp_10_i_RNIORIF1[2:2]),.I3(v_shl1_5_0_0_c2),.I4(s_exp_10_i_RNIE6AQ1[2:2]),.I5(un1_s_exp_10a_3_1),.LO(N_717));
defparam desc1535.INIT=64'h65A69A59AAAAAAAA;
  LUT4_L desc1536(.I0(s_zeros[2:2]),.I1(s_exp_10_i_RNIORIF1[2:2]),.I2(v_shl1_5_0_0_c2),.I3(un1_s_exp_10a_3_1),.LO(N_716));
defparam desc1536.INIT=16'h69AA;
  LUT5_L desc1537(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_263),.I4(N_265),.LO(N_268));
defparam desc1537.INIT=32'h101F000F;
  LUT5_L desc1538(.I0(s_shl2[3:3]),.I1(s_shl2[5:5]),.I2(N_137),.I3(N_129),.I4(N_153),.LO(i104_mux));
defparam desc1538.INIT=32'h0123CDEF;
  LUT4_L desc1539(.I0(s_shl2[4:4]),.I1(s_shl2[5:5]),.I2(N_153),.I3(N_1167),.LO(N_1168));
defparam desc1539.INIT=16'h7520;
  LUT6_L desc1540(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_297),.I3(N_265),.I4(N_289),.I5(N_280),.LO(N_376));
defparam desc1540.INIT=64'hFE76BA32DC549810;
  LUT6_L desc1541(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_327),.I3(N_370),.I4(N_360),.I5(N_361),.LO(N_372));
defparam desc1541.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc1542(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_327),.I4(N_106),.I5(N_360),.O(N_363));
defparam desc1542.INIT=64'h3715331126042200;
  LUT6_L desc1543(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(s_frac2a_2_111),.I4(N_265),.I5(N_289),.LO(N_291));
defparam desc1543.INIT=64'h3733151126220400;
  LUT6_L desc1544(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_101),.I4(N_109),.I5(N_234),.LO(N_235));
defparam desc1544.INIT=64'h5F575D550A020800;
  LUT3_L desc1545(.I0(s_shl2[4:4]),.I1(N_190),.I2(N_228),.LO(N_229));
defparam desc1545.INIT=8'hD8;
  LUT6_L desc1546(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_101),.I4(N_218),.I5(N_109),.LO(N_221));
defparam desc1546.INIT=64'h1715060413110200;
  LUT6_L desc1547(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_1140),.I3(N_1096),.I4(N_1093),.I5(N_1094),.LO(N_1142));
defparam desc1547.INIT=64'hFE76BA32DC549810;
  LUT6_L desc1548(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_103),.I4(N_111),.I5(N_116),.LO(N_1112));
defparam desc1548.INIT=64'h5F575D550A020800;
  LUT5_L desc1549(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_1084),.I3(N_1085),.I4(N_1086),.LO(N_1109));
defparam desc1549.INIT=32'h76325410;
  LUT6_L desc1550(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_1102),.I4(N_103),.I5(N_111),.LO(N_1104));
defparam desc1550.INIT=64'h1706150413021100;
  LUT5_L desc1551(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_1096),.I3(N_1093),.I4(N_1094),.LO(N_1098));
defparam desc1551.INIT=32'h75643120;
  LUT6_L desc1552(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_25_0),.I3(N_1084),.I4(N_1085),.I5(N_1086),.LO(N_1087));
defparam desc1552.INIT=64'hFEBADC9876325410;
  LUT4_L desc1553(.I0(s_shl2[4:4]),.I1(s_shl2[5:5]),.I2(N_318),.I3(N_161_0),.LO(N_78_0));
defparam desc1553.INIT=16'h3120;
  LUT5_L un4_s_lost_c4_cZ(.I0(s_r_zeros[2:2]),.I1(s_r_zeros[3:3]),.I2(un4_s_lost_c2),.I3(un2_s_lost_ac0_5_lut6_2_O5),.I4(un2_s_lost_axbxc3),.LO(un4_s_lost_c4));
defparam un4_s_lost_c4_cZ.INIT=32'hF7733110;
  LUT6 un1_s_expo3_cZ(.I0(s_frac_rnd[24:24]),.I1(s_expo2b[7:7]),.I2(s_expo2b[6:6]),.I3(s_expo2b[4:4]),.I4(s_expo2b[5:5]),.I5(un7_s_expo3_c4),.O(un1_s_expo3));
defparam un1_s_expo3_cZ.INIT=64'h2AAAAAAAAAAAAAAA;
  LUT6_L desc1554(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_1140),.I3(N_1093),.I4(N_1094),.I5(N_1152),.LO(N_410));
defparam desc1554.INIT=64'hEAC86240FBD97351;
  LUT6_L desc1555(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_1154),.I3(N_370),.I4(N_360),.I5(N_361),.LO(N_1156));
defparam desc1555.INIT=64'hEFABCD8967234501;
  LUT6_L desc1556(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(un1_s_shr2_1_4),.I4(N_342),.I5(N_101),.LO(N_344));
defparam desc1556.INIT=64'h010001FF000000FF;
  LUT6_L desc1557(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_297),.I3(N_304),.I4(N_289),.I5(N_296),.LO(N_307));
defparam desc1557.INIT=64'hA8B92031ECFD6475;
  LUT6_L desc1558(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_297),.I3(N_289),.I4(N_280),.I5(N_296),.LO(N_299));
defparam desc1558.INIT=64'hEAC86240FBD97351;
  LUT6_L desc1559(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_25_0),.I3(N_1084),.I4(N_1085),.I5(N_1128),.LO(N_1147));
defparam desc1559.INIT=64'hEAC86240FBD97351;
  LUT5_L desc1560(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_64_0_0),.I4(N_1086),.LO(N_67_0_0));
defparam desc1560.INIT=32'h101F000F;
  LUT6_L desc1561(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(un1_s_shr2_1_4),.I4(N_44_1),.I5(N_103),.LO(N_49_0_0));
defparam desc1561.INIT=64'h010001FF000000FF;
  LUT5_L desc1562(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_938),.I4(N_1096),.LO(N_57_0));
defparam desc1562.INIT=32'h101F000F;
  LUT5_L desc1563(.I0(s_shl2[4:4]),.I1(s_shl2[5:5]),.I2(un1_s_shr2_1_4),.I3(N_423),.I4(N_153),.LO(N_1163));
defparam desc1563.INIT=32'h101F000F;
  LUT6 desc1564(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(N_327),.I3(un1_s_shr2_1_4),.I4(N_349),.I5(N_361),.O(N_354));
defparam desc1564.INIT=64'h51FF510040FF4000;
  LUT6_L desc1565(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_278),.I4(N_265),.I5(N_280),.LO(N_283));
defparam desc1565.INIT=64'h505F101F404F000F;
  LUT4_L desc1566(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_201),.I3(N_206),.LO(N_208));
defparam desc1566.INIT=16'h4703;
  LUT6_L desc1567(.I0(s_shl2[4:4]),.I1(s_shr2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_115_i),.I4(s_frac2a_1_109),.I5(N_190),.LO(N_192));
defparam desc1567.INIT=64'h535F505C030F000C;
  LUT6_L desc1568(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_158),.I4(N_1096),.I5(N_1094),.LO(N_1134));
defparam desc1568.INIT=64'h5F501F104F400F00;
  LUT6_L desc1569(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(un1_s_shr2_1_4),.I3(N_85_0_0),.I4(N_1085),.I5(N_1086),.LO(N_87_0_0));
defparam desc1569.INIT=64'h505F404F101F000F;
  LUT4_L desc1570(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_74_0_0),.I3(N_77_0),.LO(N_79_0));
defparam desc1570.INIT=16'h4703;
  LUT6 un2_s_exp_10a_ac0_5_RNISRBP1(.I0(s_exp_10_i[8:8]),.I1(s_exp_10_i[7:7]),.I2(s_exp_10_i[6:6]),.I3(s_exp_10_i[5:5]),.I4(s_exp_10_i[4:4]),.I5(un2_s_exp_10a_c4),.O(N_6484_i));
defparam un2_s_exp_10a_ac0_5_RNISRBP1.INIT=64'h9555555555555555;
  LUT6_L desc1571(.I0(N_1245),.I1(m107_i_a2_7_0),.I2(N_1253),.I3(N_434_i_0),.I4(N_1246),.I5(N_1267),.LO(N_1358));
defparam desc1571.INIT=64'h0000EEEA0000EAEA;
  LUT6_L desc1572(.I0(s_fract_48_i[37:37]),.I1(s_fract_48_i[40:40]),.I2(s_fract_48_i[38:38]),.I3(s_fract_48_i[39:39]),.I4(s_fract_48_i[41:41]),.I5(N_686),.LO(N_622));
defparam desc1572.INIT=64'hAFABAFABAFABAFAA;
  LUT5_L desc1573(.I0(s_fract_48_i[1:1]),.I1(N_677),.I2(N_709),.I3(N_669_0),.I4(N_668_3),.LO(v_count_49[4:4]));
defparam desc1573.INIT=32'hCCCC4000;
  LUT4_L desc1574(.I0(s_zeros[4:4]),.I1(s_exp_10_i_RNI5I152[2:2]),.I2(v_shl1_5_0_0_c4),.I3(un1_s_exp_10a_3_1),.LO(N_718));
defparam desc1574.INIT=16'h69AA;
  LUT6 desc1575(.I0(s_frac_rnd[24:24]),.I1(s_expo2b[7:7]),.I2(s_expo2b[6:6]),.I3(s_expo2b[4:4]),.I4(s_expo2b[5:5]),.I5(un7_s_expo3_c4),.O(s_expo3[7:7]));
defparam desc1575.INIT=64'hECCCCCCCCCCCCCCC;
  LUT5_L desc1576(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_223),.I3(N_219),.I4(N_404),.LO(N_406));
defparam desc1576.INIT=32'hFC74B830;
  LUT5_L desc1577(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_399),.I3(N_368),.I4(s_frac2a_1_141_RNIA10R),.LO(N_401));
defparam desc1577.INIT=32'hC840FB73;
  LUT6_L desc1578(.I0(s_shl2[4:4]),.I1(s_shl2[5:5]),.I2(un1_s_shr2_1_4),.I3(N_161_0),.I4(N_382),.I5(i40_mux),.LO(N_389));
defparam desc1578.INIT=64'h70507F5F20002F0F;
  LUT5_L desc1579(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_214),.I3(N_234),.I4(N_254),.LO(N_256));
defparam desc1579.INIT=32'hB830FC74;
  LUT5_L desc1580(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_1137),.I3(N_1141),.I4(N_1153),.LO(N_184));
defparam desc1580.INIT=32'hB830FC74;
  LUT5_L desc1581(.I0(s_shl2[4:4]),.I1(N_82_0),.I2(un1_s_shr2_1_4),.I3(N_116),.I4(N_1121),.LO(N_1123));
defparam desc1581.INIT=32'hAC0CFC5C;
  LUT5_L desc1582(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_56_0),.I3(N_1103),.I4(N_1115),.LO(N_1117));
defparam desc1582.INIT=32'hFC74B830;
  LUT6_L desc1583(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(un1_s_shr2_1_4),.I3(N_1081),.I4(s_frac2a_1_141_RNIA10R),.I5(N_195),.LO(s_frac2a_3[2:2]));
defparam desc1583.INIT=64'h5545776710003222;
  LUT5_L desc1584(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_161),.I3(N_382),.I4(N_921),.LO(s_frac2a_3[0:0]));
defparam desc1584.INIT=32'h51734062;
  LUT3 s_exp_10b_s_9_RNO(.I0(s_exp_10_i[9:9]),.I1(s_exp_10_i[8:8]),.I2(un2_s_exp_10a_c8),.O(N_6485_i));
defparam s_exp_10b_s_9_RNO.INIT=8'h95;
  LUT6_L desc1585(.I0(s_fract_48_i[7:7]),.I1(s_fract_48_i[15:15]),.I2(N_1273),.I3(N_1370),.I4(N_1281_2),.I5(N_331_0),.LO(v_count_49_i_i[3:3]));
defparam desc1585.INIT=64'hFF00FF0055005400;
  LUT5_L desc1586(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_330),.I3(N_333),.I4(N_337),.LO(s_frac2a_3[1:1]));
defparam desc1586.INIT=32'h76325410;
  LUT6 un6_s_exp_10a_cZ(.I0(s_exp_10_i[9:9]),.I1(s_exp_10_i[8:8]),.I2(un2_s_exp_10a_c8),.I3(N_6482_i),.I4(N_6483_i),.I5(un5_s_exp_10a_1),.O(un6_s_exp_10a));
defparam un6_s_exp_10a_cZ.INIT=64'hEB6A6A6A6A6A6A6A;
  LUT6_L desc1587(.I0(s_expo2b[0:0]),.I1(s_output_o25_sn),.I2(s_expo2b[3:3]),.I3(s_expo2b[1:1]),.I4(s_expo2b[2:2]),.I5(un1_s_expo3),.LO(s_output_o_m0[26:26]));
defparam desc1587.INIT=64'h1230303030303030;
  LUT6_L desc1588(.I0(s_output_o25_sn),.I1(s_expo2b[6:6]),.I2(s_expo2b[4:4]),.I3(s_expo2b[5:5]),.I4(un7_s_expo3_c4),.I5(un1_s_expo3),.LO(s_output_o_m0[29:29]));
defparam desc1588.INIT=64'h1444444444444444;
  LUT5_L desc1589(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_271),.I3(N_275),.I4(N_268),.LO(s_frac2a_3[3:3]));
defparam desc1589.INIT=32'h15370426;
  LUT5_L desc1590(.I0(s_shl2[4:4]),.I1(un1_s_shr2_1_4),.I2(N_1165),.I3(N_1167),.I4(i104_mux),.LO(N_441));
defparam desc1590.INIT=32'hB830FC74;
  LUT6_L desc1591(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.I4(N_658),.I5(N_688),.LO(v_count_49_0_4));
defparam desc1591.INIT=64'hFFFFFBFAFFFFAAAA;
  LUT6_L desc1592(.I0(s_fract_48_i[27:27]),.I1(s_fract_48_i[25:25]),.I2(N_326_2),.I3(N_1252),.I4(N_326_0_3),.I5(N_1340),.LO(N_326_2_0));
defparam desc1592.INIT=64'h0000000000100000;
  LUT6 un2_s_exp_10a_ac0_3_lut6_2_RNIQPBD7(.I0(un5_v_shr1_c3),.I1(s_exp_10_i_RNIE6AQ1[2:2]),.I2(s_exp_10_i_RNI5I152[2:2]),.I3(N_6482_i),.I4(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91),.I5(un6_s_exp_10a),.O(v_shr1_4[6:6]));
defparam un2_s_exp_10a_ac0_3_lut6_2_RNIQPBD7.INIT=64'hFF00FD0200000000;
  LUT5_L desc1593(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_223),.I3(N_217),.I4(N_344),.LO(s_frac2a_3[4:4]));
defparam desc1593.INIT=32'h31752064;
  LUT5_L desc1594(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_71_0_0),.I3(N_69_0),.I4(N_67_0_0),.LO(s_frac2a_3[7:7]));
defparam desc1594.INIT=32'h31752064;
  LUT5_L desc1595(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_56_0),.I3(N_52_0),.I4(N_49_0_0),.LO(s_frac2a_3[6:6]));
defparam desc1595.INIT=32'h31752064;
  LUT5_L desc1596(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_60_0),.I3(N_64_0),.I4(N_57_0),.LO(s_frac2a_3[5:5]));
defparam desc1596.INIT=32'h15370426;
  LUT6_L desc1597(.I0(s_zeros[5:5]),.I1(s_zeros[4:4]),.I2(s_exp_10_i_RNI5I152[2:2]),.I3(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91),.I4(v_shl1_5_0_0_c4),.I5(un1_s_exp_10a_3_1),.LO(N_719));
defparam desc1597.INIT=64'h659AA659AAAAAAAA;
  LUT5_L desc1598(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_1165),.I3(N_169),.I4(N_1163),.LO(s_frac2a_3[8:8]));
defparam desc1598.INIT=32'h75316420;
  LUT5_L desc1599(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_286),.I3(N_284),.I4(N_283),.LO(s_frac2a_3[11:11]));
defparam desc1599.INIT=32'h31752064;
  LUT5_L desc1600(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_214),.I3(N_211),.I4(N_208),.LO(s_frac2a_3[12:12]));
defparam desc1600.INIT=32'h31752064;
  LUT5_L desc1601(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_1137),.I3(s_frac2a_1_124_RNIEJB51_O6),.I4(N_1134),.LO(s_frac2a_3[13:13]));
defparam desc1601.INIT=32'h31752064;
  LUT5_L desc1602(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_1090),.I3(N_1083),.I4(N_87_0_0),.LO(s_frac2a_3[15:15]));
defparam desc1602.INIT=32'h31752064;
  LUT6_L desc1603(.I0(s_fract_48_i[27:27]),.I1(N_707),.I2(N_582),.I3(N_650),.I4(N_688),.I5(v_count_49_0_4),.LO(v_count_49_0));
defparam desc1603.INIT=64'hFFFFFFFFFF0EFF00;
  LUT6_L desc1604(.I0(v_count_49_i_o2_1_i_a2_lut6_2_O6[2:2]),.I1(v_count_49_i_o2_0_i_a2_lut6_2_O6[2:2]),.I2(N_638),.I3(N_673),.I4(N_677),.I5(N_637),.LO(s_r_zeros_RNO_0[2:2]));
defparam desc1604.INIT=64'hF8000000F0000000;
  LUT6 un4_s_lost_c6_cZ(.I0(s_r_zeros[4:4]),.I1(s_r_zeros[5:5]),.I2(s_shr2[5:5]),.I3(s_shr2[4:4]),.I4(un2_s_lost_c4),.I5(un4_s_lost_c4),.O(un4_s_lost_c6));
defparam un4_s_lost_c6_cZ.INIT=64'h17F3F37103717130;
  LUT6_L desc1605(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.I2(s_fract_48_i[12:12]),.I3(s_fract_48_i[10:10]),.I4(s_fract_48_i[11:11]),.I5(N_1350),.LO(N_1271));
defparam desc1605.INIT=64'hDCDCDDDDDCDCDDDC;
  LUT5 un16_s_roundup_cZ(.I0(s_frac2a[20:20]),.I1(s_frac2a[21:21]),.I2(s_frac2a[23:23]),.I3(un3_s_ine_o_0),.I4(un4_s_lost_c6),.O(un16_s_roundup));
defparam un16_s_roundup_cZ.INIT=32'hFFFFFFFE;
  LUT5 un3_s_ine_o_cZ(.I0(s_frac2a[20:20]),.I1(s_frac2a[21:21]),.I2(s_frac2a[22:22]),.I3(un3_s_ine_o_0),.I4(un4_s_lost_c6),.O(un3_s_ine_o));
defparam un3_s_ine_o_cZ.INIT=32'hFFFFFFFE;
  LUT6_L desc1606(.I0(s_fract_48_i[19:19]),.I1(s_fract_48_i[18:18]),.I2(N_663_3),.I3(v_count_49_i_o2_0_i_a2_lut6_2_O6[2:2]),.I4(v_count_49_i_o3_1[1:1]),.I5(N_626),.LO(N_663_2));
defparam desc1606.INIT=64'hF0F01000F0F00000;
  LUT6_L desc1607(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(N_1353),.I3(N_326_1),.I4(N_23_0_2),.I5(N_326_2_0),.LO(N_23_0_4));
defparam desc1607.INIT=64'hFFFFFF20FFFF2020;
  LUT6_L desc1608(.I0(s_fract_48_i[31:31]),.I1(s_fract_48_i[32:32]),.I2(N_314_1),.I3(N_1361),.I4(N_173),.I5(N_1365),.LO(N_314));
defparam desc1608.INIT=64'hF1F1F1F1F1F0F1F1;
  LUT6 desc1609(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[34:34]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[32:32]),.I4(N_641_1),.I5(N_622),.O(N_641));
defparam desc1609.INIT=64'hFFFF0031FFFF0030;
  LUT6 desc1610(.I0(s_fract_48_i[29:29]),.I1(N_1260),.I2(N_1305),.I3(N_1353),.I4(N_320_0),.I5(N_1271),.O(N_23_0_3));
defparam desc1610.INIT=64'h3300100010001000;
  LUT6_L desc1611(.I0(s_fract_48_i[5:5]),.I1(s_fract_48_i[7:7]),.I2(v_count_49_i_o3_i_a2_lut6_2_O6[3:3]),.I3(s_fract_48_i_RNIEUJ9_O5[3:3]),.I4(N_610),.I5(s_r_zeros_RNO_0[2:2]),.LO(N_566_i));
defparam desc1611.INIT=64'h00000000EF00FF00;
  LUT6_L desc1612(.I0(s_frac_rnd[23:23]),.I1(s_frac_rnd[22:22]),.I2(s_output_o25_sn),.I3(s_output_o_sn_N_5_mux),.I4(un1_s_expo3),.I5(s_output_o_sm0),.LO(s_output_o[22:22]));
defparam desc1612.INIT=64'h00FF00FF0A0A0C0C;
  LUT6_L desc1613(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[38:38]),.I4(N_1249),.I5(N_314),.LO(N_62_1));
defparam desc1613.INIT=64'h0000FFCD0000FFCC;
  LUT6 un16_s_roundup_RNIMA661(.I0(s_frac2a[22:22]),.I1(s_sign_i),.I2(s_rmode_i[0:0]),.I3(s_rmode_i[1:1]),.I4(un16_s_roundup),.I5(un3_s_ine_o),.O(s_roundup));
defparam un16_s_roundup_RNIMA661.INIT=64'hC30AC300000A0000;
  LUT6 desc1614(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[28:28]),.I2(N_653),.I3(N_582),.I4(N_641),.I5(N_688),.O(v_count_49_1_1));
defparam desc1614.INIT=64'hF0F1F0F0F0F0F0F0;
  LUT3_L desc1615(.I0(s_frac2a[39:39]),.I1(s_frac_rnd_3_0_s_16),.I2(s_roundup),.LO(s_frac_rnd_3[16:16]));
defparam desc1615.INIT=8'hCA;
  LUT6_L desc1616(.I0(N_672),.I1(v_count_49_i_a2_0_lut6_2_O6[1:1]),.I2(N_1308),.I3(v_count_49_i_0[1:1]),.I4(N_662),.I5(N_663_2),.LO(N_564_i));
defparam desc1616.INIT=64'h000000F7000000FF;
  LUT6_L desc1617(.I0(s_fract_48_i[15:15]),.I1(N_654),.I2(N_679),.I3(v_count_49_1_3),.I4(v_count_49_1_1),.I5(v_count_49_0),.LO(v_count_49[0:0]));
defparam desc1617.INIT=64'hFFFFFFFFFFFFFFEC;
  LUT3 desc1618(.I0(s_exp_10_i[1:1]),.I1(s_exp_10_i[0:0]),.I2(s_fract_48_i[47:47]),.O(un5_v_shr1_axb1));
defparam desc1618.INIT=8'h6A;
  LUT5 desc1619(.I0(s_zeros[2:2]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_fract_48_i[47:47]),.O(s_exp_10b_axb_2));
defparam desc1619.INIT=32'h69999999;
  LUT4 desc1620(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(s_exp_10_i[0:0]),.I3(s_fract_48_i[47:47]),.O(s_exp_10_i_RNIORIF1[2:2]));
defparam desc1620.INIT=16'h6AAA;
  LUT5 un2_s_exp_10a_ac0_1_lut6_2_RNIDG351(.I0(s_zeros[4:4]),.I1(s_exp_10_i[4:4]),.I2(s_exp_10_i[2:2]),.I3(s_exp_10_i[3:3]),.I4(un2_s_exp_10a_c2),.O(s_exp_10b_axb_4));
defparam un2_s_exp_10a_ac0_1_lut6_2_RNIDG351.INIT=32'h69999999;
  LUT5 desc1621(.I0(s_zeros[5:5]),.I1(s_exp_10_i[5:5]),.I2(s_exp_10_i[4:4]),.I3(s_exp_10_i[3:3]),.I4(un2_s_exp_10a_c3),.O(s_exp_10b_axb_5));
defparam desc1621.INIT=32'h69999999;
  LUT4 un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91_cZ(.I0(s_exp_10_i[5:5]),.I1(s_exp_10_i[4:4]),.I2(s_exp_10_i[3:3]),.I3(un2_s_exp_10a_c3),.O(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91));
defparam un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91_cZ.INIT=16'h6AAA;
  LUT5 un2_s_exp_10a_ac0_3_lut6_2_RNIMNHK1(.I0(s_exp_10_i[6:6]),.I1(s_exp_10_i[5:5]),.I2(s_exp_10_i[4:4]),.I3(s_exp_10_i[3:3]),.I4(un2_s_exp_10a_c3),.O(N_6482_i));
defparam un2_s_exp_10a_ac0_3_lut6_2_RNIMNHK1.INIT=32'h95555555;
  LUT5 s_exp_10b_cry_6_RNO_cZ(.I0(s_exp_10_i[6:6]),.I1(s_exp_10_i[5:5]),.I2(s_exp_10_i[4:4]),.I3(s_exp_10_i[3:3]),.I4(un2_s_exp_10a_c3),.O(s_exp_10b_cry_6_RNO));
defparam s_exp_10b_cry_6_RNO_cZ.INIT=32'h6AAAAAAA;
  LUT5 un2_s_exp_10a_ac0_5_RNI1CKE1(.I0(s_exp_10_i[7:7]),.I1(s_exp_10_i[6:6]),.I2(s_exp_10_i[5:5]),.I3(s_exp_10_i[4:4]),.I4(un2_s_exp_10a_c4),.O(N_6483_i));
defparam un2_s_exp_10a_ac0_5_RNI1CKE1.INIT=32'h95555555;
  LUT5 s_exp_10b_cry_7_RNO_cZ(.I0(s_exp_10_i[7:7]),.I1(s_exp_10_i[6:6]),.I2(s_exp_10_i[5:5]),.I3(s_exp_10_i[4:4]),.I4(un2_s_exp_10a_c4),.O(s_exp_10b_cry_7_RNO));
defparam s_exp_10b_cry_7_RNO_cZ.INIT=32'h6AAAAAAA;
  XORCY s_frac_rnd_3_0_s_24_cZ(.LI(s_frac_rnd_3_0_axb_24),.CI(s_frac_rnd_3_0_cry_23),.O(s_frac_rnd_3_0_s_24));
  XORCY s_frac_rnd_3_0_s_23_cZ(.LI(s_frac_rnd_3_0_axb_23),.CI(s_frac_rnd_3_0_cry_22),.O(s_frac_rnd_3_0_s_23));
  MUXCY_L s_frac_rnd_3_0_cry_23_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_22),.S(s_frac_rnd_3_0_axb_23),.LO(s_frac_rnd_3_0_cry_23));
  XORCY s_frac_rnd_3_0_s_22_cZ(.LI(s_frac_rnd_3_0_axb_22),.CI(s_frac_rnd_3_0_cry_21),.O(s_frac_rnd_3_0_s_22));
  MUXCY_L s_frac_rnd_3_0_cry_22_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_21),.S(s_frac_rnd_3_0_axb_22),.LO(s_frac_rnd_3_0_cry_22));
  XORCY s_frac_rnd_3_0_s_21_cZ(.LI(s_frac_rnd_3_0_axb_21),.CI(s_frac_rnd_3_0_cry_20),.O(s_frac_rnd_3_0_s_21));
  MUXCY_L s_frac_rnd_3_0_cry_21_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_20),.S(s_frac_rnd_3_0_axb_21),.LO(s_frac_rnd_3_0_cry_21));
  XORCY s_frac_rnd_3_0_s_20_cZ(.LI(s_frac_rnd_3_0_axb_20),.CI(s_frac_rnd_3_0_cry_19),.O(s_frac_rnd_3_0_s_20));
  MUXCY_L s_frac_rnd_3_0_cry_20_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_19),.S(s_frac_rnd_3_0_axb_20),.LO(s_frac_rnd_3_0_cry_20));
  XORCY s_frac_rnd_3_0_s_19_cZ(.LI(s_frac_rnd_3_0_axb_19),.CI(s_frac_rnd_3_0_cry_18),.O(s_frac_rnd_3_0_s_19));
  MUXCY_L s_frac_rnd_3_0_cry_19_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_18),.S(s_frac_rnd_3_0_axb_19),.LO(s_frac_rnd_3_0_cry_19));
  XORCY s_frac_rnd_3_0_s_18_cZ(.LI(s_frac_rnd_3_0_axb_18),.CI(s_frac_rnd_3_0_cry_17),.O(s_frac_rnd_3_0_s_18));
  MUXCY_L s_frac_rnd_3_0_cry_18_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_17),.S(s_frac_rnd_3_0_axb_18),.LO(s_frac_rnd_3_0_cry_18));
  XORCY s_frac_rnd_3_0_s_17_cZ(.LI(s_frac_rnd_3_0_axb_17),.CI(s_frac_rnd_3_0_cry_16),.O(s_frac_rnd_3_0_s_17));
  MUXCY_L s_frac_rnd_3_0_cry_17_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_16),.S(s_frac_rnd_3_0_axb_17),.LO(s_frac_rnd_3_0_cry_17));
  XORCY s_frac_rnd_3_0_s_16_cZ(.LI(s_frac_rnd_3_0_axb_16),.CI(s_frac_rnd_3_0_cry_15),.O(s_frac_rnd_3_0_s_16));
  MUXCY_L s_frac_rnd_3_0_cry_16_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_15),.S(s_frac_rnd_3_0_axb_16),.LO(s_frac_rnd_3_0_cry_16));
  XORCY s_frac_rnd_3_0_s_15_cZ(.LI(s_frac_rnd_3_0_axb_15),.CI(s_frac_rnd_3_0_cry_14),.O(s_frac_rnd_3_0_s_15));
  MUXCY_L s_frac_rnd_3_0_cry_15_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_14),.S(s_frac_rnd_3_0_axb_15),.LO(s_frac_rnd_3_0_cry_15));
  XORCY s_frac_rnd_3_0_s_14_cZ(.LI(s_frac_rnd_3_0_axb_14),.CI(s_frac_rnd_3_0_cry_13),.O(s_frac_rnd_3_0_s_14));
  MUXCY_L s_frac_rnd_3_0_cry_14_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_13),.S(s_frac_rnd_3_0_axb_14),.LO(s_frac_rnd_3_0_cry_14));
  XORCY s_frac_rnd_3_0_s_13_cZ(.LI(s_frac_rnd_3_0_axb_13),.CI(s_frac_rnd_3_0_cry_12),.O(s_frac_rnd_3_0_s_13));
  MUXCY_L s_frac_rnd_3_0_cry_13_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_12),.S(s_frac_rnd_3_0_axb_13),.LO(s_frac_rnd_3_0_cry_13));
  XORCY s_frac_rnd_3_0_s_12_cZ(.LI(s_frac_rnd_3_0_axb_12),.CI(s_frac_rnd_3_0_cry_11),.O(s_frac_rnd_3_0_s_12));
  MUXCY_L s_frac_rnd_3_0_cry_12_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_11),.S(s_frac_rnd_3_0_axb_12),.LO(s_frac_rnd_3_0_cry_12));
  XORCY s_frac_rnd_3_0_s_11_cZ(.LI(s_frac_rnd_3_0_axb_11),.CI(s_frac_rnd_3_0_cry_10),.O(s_frac_rnd_3_0_s_11));
  MUXCY_L s_frac_rnd_3_0_cry_11_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_10),.S(s_frac_rnd_3_0_axb_11),.LO(s_frac_rnd_3_0_cry_11));
  XORCY s_frac_rnd_3_0_s_10_cZ(.LI(s_frac_rnd_3_0_axb_10),.CI(s_frac_rnd_3_0_cry_9),.O(s_frac_rnd_3_0_s_10));
  MUXCY_L s_frac_rnd_3_0_cry_10_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_9),.S(s_frac_rnd_3_0_axb_10),.LO(s_frac_rnd_3_0_cry_10));
  XORCY s_frac_rnd_3_0_s_9_cZ(.LI(s_frac_rnd_3_0_axb_9),.CI(s_frac_rnd_3_0_cry_8),.O(s_frac_rnd_3_0_s_9));
  MUXCY_L s_frac_rnd_3_0_cry_9_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_8),.S(s_frac_rnd_3_0_axb_9),.LO(s_frac_rnd_3_0_cry_9));
  XORCY s_frac_rnd_3_0_s_8_cZ(.LI(s_frac_rnd_3_0_axb_8),.CI(s_frac_rnd_3_0_cry_7),.O(s_frac_rnd_3_0_s_8));
  MUXCY_L s_frac_rnd_3_0_cry_8_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_7),.S(s_frac_rnd_3_0_axb_8),.LO(s_frac_rnd_3_0_cry_8));
  XORCY s_frac_rnd_3_0_s_7_cZ(.LI(s_frac_rnd_3_0_axb_7),.CI(s_frac_rnd_3_0_cry_6),.O(s_frac_rnd_3_0_s_7));
  MUXCY_L s_frac_rnd_3_0_cry_7_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_6),.S(s_frac_rnd_3_0_axb_7),.LO(s_frac_rnd_3_0_cry_7));
  XORCY s_frac_rnd_3_0_s_6_cZ(.LI(s_frac_rnd_3_0_axb_6),.CI(s_frac_rnd_3_0_cry_5),.O(s_frac_rnd_3_0_s_6));
  MUXCY_L s_frac_rnd_3_0_cry_6_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_5),.S(s_frac_rnd_3_0_axb_6),.LO(s_frac_rnd_3_0_cry_6));
  XORCY s_frac_rnd_3_0_s_5_cZ(.LI(s_frac_rnd_3_0_axb_5),.CI(s_frac_rnd_3_0_cry_4),.O(s_frac_rnd_3_0_s_5));
  MUXCY_L s_frac_rnd_3_0_cry_5_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_4),.S(s_frac_rnd_3_0_axb_5),.LO(s_frac_rnd_3_0_cry_5));
  XORCY s_frac_rnd_3_0_s_4_cZ(.LI(s_frac_rnd_3_0_axb_4),.CI(s_frac_rnd_3_0_cry_3),.O(s_frac_rnd_3_0_s_4));
  MUXCY_L s_frac_rnd_3_0_cry_4_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_3),.S(s_frac_rnd_3_0_axb_4),.LO(s_frac_rnd_3_0_cry_4));
  XORCY s_frac_rnd_3_0_s_3_cZ(.LI(s_frac_rnd_3_0_axb_3),.CI(s_frac_rnd_3_0_cry_2),.O(s_frac_rnd_3_0_s_3));
  MUXCY_L s_frac_rnd_3_0_cry_3_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_2),.S(s_frac_rnd_3_0_axb_3),.LO(s_frac_rnd_3_0_cry_3));
  XORCY s_frac_rnd_3_0_s_2_cZ(.LI(s_frac_rnd_3_0_axb_2),.CI(s_frac_rnd_3_0_cry_1),.O(s_frac_rnd_3_0_s_2));
  MUXCY_L s_frac_rnd_3_0_cry_2_cZ(.DI(GND),.CI(s_frac_rnd_3_0_cry_1),.S(s_frac_rnd_3_0_axb_2),.LO(s_frac_rnd_3_0_cry_2));
  XORCY s_frac_rnd_3_0_s_1_cZ(.LI(s_frac_rnd_3_0_axb_1),.CI(s_frac2a[23:23]),.O(s_frac_rnd_3_0_s_1));
  MUXCY_L s_frac_rnd_3_0_cry_1_cZ(.DI(GND),.CI(s_frac2a[23:23]),.S(s_frac_rnd_3_0_axb_1),.LO(s_frac_rnd_3_0_cry_1));
  XORCY s_exp_10b_s_9(.LI(N_6485_i),.CI(s_exp_10b_cry_8),.O(s_exp_10b[9:9]));
  XORCY s_exp_10b_s_8(.LI(N_6484_i),.CI(s_exp_10b_cry_7),.O(s_exp_10b[8:8]));
  MUXCY_L s_exp_10b_cry_8_cZ(.DI(VCC),.CI(s_exp_10b_cry_7),.S(N_6484_i),.LO(s_exp_10b_cry_8));
  XORCY s_exp_10b_s_7(.LI(N_6483_i),.CI(s_exp_10b_cry_6),.O(s_exp_10b[7:7]));
  MUXCY_L s_exp_10b_cry_7_cZ(.DI(s_exp_10b_cry_7_RNO),.CI(s_exp_10b_cry_6),.S(N_6483_i),.LO(s_exp_10b_cry_7));
  XORCY s_exp_10b_s_6(.LI(N_6482_i),.CI(s_exp_10b_cry_5),.O(s_exp_10b[6:6]));
  MUXCY_L s_exp_10b_cry_6_cZ(.DI(s_exp_10b_cry_6_RNO),.CI(s_exp_10b_cry_5),.S(N_6482_i),.LO(s_exp_10b_cry_6));
  XORCY s_exp_10b_s_5(.LI(s_exp_10b_axb_5),.CI(s_exp_10b_cry_4),.O(s_exp_10b[5:5]));
  MUXCY_L s_exp_10b_cry_5_cZ(.DI(un2_s_exp_10a_ac0_3_lut6_2_RNIT9Q91),.CI(s_exp_10b_cry_4),.S(s_exp_10b_axb_5),.LO(s_exp_10b_cry_5));
  XORCY s_exp_10b_s_4(.LI(s_exp_10b_axb_4),.CI(s_exp_10b_cry_3),.O(s_exp_10b[4:4]));
  MUXCY_L s_exp_10b_cry_4_cZ(.DI(s_exp_10_i_RNI5I152[2:2]),.CI(s_exp_10b_cry_3),.S(s_exp_10b_axb_4),.LO(s_exp_10b_cry_4));
  XORCY s_exp_10b_s_3(.LI(s_exp_10b_axb_3),.CI(s_exp_10b_cry_2),.O(s_exp_10b[3:3]));
  MUXCY_L s_exp_10b_cry_3_cZ(.DI(s_exp_10_i_RNIE6AQ1[2:2]),.CI(s_exp_10b_cry_2),.S(s_exp_10b_axb_3),.LO(s_exp_10b_cry_3));
  XORCY s_exp_10b_s_2(.LI(s_exp_10b_axb_2),.CI(s_exp_10b_cry_1),.O(s_exp_10b[2:2]));
  MUXCY_L s_exp_10b_cry_2_cZ(.DI(s_exp_10_i_RNIORIF1[2:2]),.CI(s_exp_10b_cry_1),.S(s_exp_10b_axb_2),.LO(s_exp_10b_cry_2));
  XORCY s_exp_10b_s_1(.LI(s_exp_10b_axb_1),.CI(s_exp_10b_cry_0),.O(s_exp_10b[1:1]));
  MUXCY_L s_exp_10b_cry_1_cZ(.DI(un5_v_shr1_axb1),.CI(s_exp_10b_cry_0),.S(s_exp_10b_axb_1),.LO(s_exp_10b_cry_1));
  MUXCY_L s_exp_10b_cry_0_cZ(.DI(s_zeros_RNI0TNS_O5),.CI(VCC),.S(s_exp_10b_i),.LO(s_exp_10b_cry_0));
  XORCY s_expo2b_s_7(.LI(s_expo2b_axb_7),.CI(s_expo2b_cry_6),.O(s_expo2b[7:7]));
  XORCY s_expo2b_s_6(.LI(s_expo2b_axb_6),.CI(s_expo2b_cry_5),.O(s_expo2b[6:6]));
  MUXCY_L s_expo2b_cry_6_cZ(.DI(s_expo1[6:6]),.CI(s_expo2b_cry_5),.S(s_expo2b_axb_6),.LO(s_expo2b_cry_6));
  XORCY s_expo2b_s_5(.LI(s_expo2b_axb_5),.CI(s_expo2b_cry_4),.O(s_expo2b[5:5]));
  MUXCY_L s_expo2b_cry_5_cZ(.DI(s_expo1[5:5]),.CI(s_expo2b_cry_4),.S(s_expo2b_axb_5),.LO(s_expo2b_cry_5));
  XORCY s_expo2b_s_4(.LI(s_expo2b_axb_4),.CI(s_expo2b_cry_3),.O(s_expo2b[4:4]));
  MUXCY_L s_expo2b_cry_4_cZ(.DI(s_expo1[4:4]),.CI(s_expo2b_cry_3),.S(s_expo2b_axb_4),.LO(s_expo2b_cry_4));
  XORCY s_expo2b_s_3(.LI(s_expo2b_axb_3),.CI(s_expo2b_cry_2),.O(s_expo2b[3:3]));
  MUXCY_L s_expo2b_cry_3_cZ(.DI(s_expo1[3:3]),.CI(s_expo2b_cry_2),.S(s_expo2b_axb_3),.LO(s_expo2b_cry_3));
  XORCY s_expo2b_s_2(.LI(s_expo2b_axb_2),.CI(s_expo2b_cry_1),.O(s_expo2b[2:2]));
  MUXCY_L s_expo2b_cry_2_cZ(.DI(s_expo1[2:2]),.CI(s_expo2b_cry_1),.S(s_expo2b_axb_2),.LO(s_expo2b_cry_2));
  XORCY s_expo2b_s_1(.LI(s_expo2b_axb_1),.CI(s_expo2b_cry_0),.O(s_expo2b[1:1]));
  MUXCY_L s_expo2b_cry_1_cZ(.DI(s_expo1[1:1]),.CI(s_expo2b_cry_0),.S(s_expo2b_axb_1),.LO(s_expo2b_cry_1));
  MUXCY_L s_expo2b_cry_0_cZ(.DI(s_expo1[0:0]),.CI(GND),.S(s_expo2b[0:0]),.LO(s_expo2b_cry_0));
  FDS desc1622(.Q(post_norm_mul_output[23:23]),.D(s_output_o_m0[23:23]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1623(.Q(post_norm_mul_output[24:24]),.D(s_output_o_m0[24:24]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1624(.Q(post_norm_mul_output[25:25]),.D(s_output_o_m0[25:25]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1625(.Q(post_norm_mul_output[26:26]),.D(s_output_o_m0[26:26]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1626(.Q(post_norm_mul_output[27:27]),.D(s_output_o_m0[27:27]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1627(.Q(post_norm_mul_output[28:28]),.D(s_output_o_m0[28:28]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1628(.Q(post_norm_mul_output[29:29]),.D(s_output_o_m0[29:29]),.C(clk_i),.S(s_output_o_sm0));
  FDS desc1629(.Q(post_norm_mul_output[30:30]),.D(s_output_o_m0[30:30]),.C(clk_i),.S(s_output_o_sm0));
  FDR desc1630(.Q(s_r_zeros[5:5]),.D(v_count_0_sqmuxa_46),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1631(.Q(s_r_zeros[4:4]),.D(v_count_49[4:4]),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1632(.Q(s_r_zeros[3:3]),.D(v_count_49_i_i[3:3]),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1633(.Q(s_r_zeros[2:2]),.D(N_566_i),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1634(.Q(s_r_zeros[1:1]),.D(N_564_i),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1635(.Q(s_r_zeros[0:0]),.D(v_count_49[0:0]),.C(clk_i),.R(s_fract_48_i[0:0]));
  FDR desc1636(.Q(s_expo1[7:7]),.D(s_expo1_5[7:7]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1637(.Q(s_expo1[6:6]),.D(s_expo1_5[6:6]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1638(.Q(s_expo1[5:5]),.D(s_expo1_5[5:5]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1639(.Q(s_expo1[4:4]),.D(s_expo1_5[4:4]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1640(.Q(s_expo1[3:3]),.D(s_expo1_5[3:3]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1641(.Q(s_expo1[2:2]),.D(s_expo1_5[2:2]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  FDR desc1642(.Q(s_expo1[1:1]),.D(s_expo1_5[1:1]),.C(clk_i),.R(un1_s_exp_10a_3_lut6_2_O6));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT5 un6_s_exp_10a_RNILFHJ8_o6(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[3:3]),.I2(s_exp_10_i[1:1]),.I3(un6_s_exp_10a),.I4(v_shr1_4[6:6]),.O(v_shr1_4_e[3:3]));
defparam un6_s_exp_10a_RNILFHJ8_o6.INIT=32'hFFFF3600;
  LUT4 un6_s_exp_10a_RNILFHJ8_o5(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(un6_s_exp_10a),.I3(v_shr1_4[6:6]),.O(v_shr1_4_e[2:2]));
defparam un6_s_exp_10a_RNILFHJ8_o5.INIT=16'hFF60;
  LUT4 desc1643(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[47:47]),.O(N_599));
defparam desc1643.INIT=16'hFAFB;
  LUT5 desc1644(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[46:46]),.I2(s_fract_48_i[45:45]),.I3(s_fract_48_i[43:43]),.I4(s_fract_48_i[47:47]),.O(N_543));
defparam desc1644.INIT=32'h00000001;
  LUT3 desc1645(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[42:42]),.I2(s_fract_48_i[47:47]),.O(N_1261));
defparam desc1645.INIT=8'hFE;
  LUT5 desc1646(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[39:39]),.I2(s_fract_48_i[42:42]),.I3(s_fract_48_i[43:43]),.I4(s_fract_48_i[47:47]),.O(N_326_0_3));
defparam desc1646.INIT=32'hFFFFAAFB;
  LUT2 desc1647(.I0(s_fract_48_i[39:39]),.I1(s_fract_48_i[33:33]),.O(N_331_1));
defparam desc1647.INIT=4'h1;
  LUT4 desc1648(.I0(s_fract_48_i[40:40]),.I1(s_fract_48_i[39:39]),.I2(s_fract_48_i[41:41]),.I3(s_fract_48_i[42:42]),.O(N_481));
defparam desc1648.INIT=16'hFFFE;
  LUT2 desc1649(.I0(s_fract_48_i[27:27]),.I1(s_fract_48_i[28:28]),.O(N_505_1_2));
defparam desc1649.INIT=4'h1;
  LUT5 desc1650(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[21:21]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[28:28]),.I4(s_fract_48_i[18:18]),.O(v_count_0_sqmuxa_47_3_4));
defparam desc1650.INIT=32'h00000001;
  LUT2 desc1651(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[4:4]),.O(N_530_1));
defparam desc1651.INIT=4'h1;
  LUT3 desc1652(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[2:2]),.O(s_fract_48_i_RNIEUJ9_O5[3:3]));
defparam desc1652.INIT=8'h01;
  LUT2 desc1653(.I0(s_r_zeros[4:4]),.I1(s_r_zeros[5:5]),.O(s_output_o25_sn));
defparam desc1653.INIT=4'h8;
  LUT5 desc1654(.I0(s_frac_rnd[0:0]),.I1(s_frac_rnd[1:1]),.I2(un1_s_expo3),.I3(s_r_zeros[4:4]),.I4(s_r_zeros[5:5]),.O(s_output_o_0[0:0]));
defparam desc1654.INIT=32'h00CACACA;
  LUT2 desc1655(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[2:2]),.O(N_1308));
defparam desc1655.INIT=4'hE;
  LUT5 desc1656(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[3:3]),.I2(s_fract_48_i[4:4]),.I3(s_fract_48_i[5:5]),.I4(s_fract_48_i[2:2]),.O(v_count_49_i_0[1:1]));
defparam desc1656.INIT=32'hAAAABBBA;
  LUT2 desc1657(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[15:15]),.O(N_320_2));
defparam desc1657.INIT=4'h1;
  LUT3 desc1658(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[16:16]),.I2(s_fract_48_i[18:18]),.O(s_zeros_2_0_i_a2_1_2_lut6_2_O5));
defparam desc1658.INIT=8'hFE;
  LUT2 desc1659(.I0(s_fract_48_i[10:10]),.I1(s_fract_48_i[11:11]),.O(N_663_3));
defparam desc1659.INIT=4'h1;
  LUT5 desc1660(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[12:12]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.I4(s_fract_48_i[8:8]),.O(N_708));
defparam desc1660.INIT=32'h00000F02;
  LUT2 desc1661(.I0(s_fract_48_i[38:38]),.I1(s_fract_48_i[32:32]),.O(N_239));
defparam desc1661.INIT=4'hE;
  LUT4 desc1662(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[37:37]),.I2(s_fract_48_i[35:35]),.I3(s_fract_48_i[38:38]),.O(N_301));
defparam desc1662.INIT=16'hFFFE;
  LUT2 desc1663(.I0(s_fract_48_i[31:31]),.I1(s_fract_48_i[33:33]),.O(N_1259));
defparam desc1663.INIT=4'hE;
  LUT5 desc1664(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.I4(N_687),.O(N_689));
defparam desc1664.INIT=32'h11111110;
  LUT2 desc1665(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[14:14]),.O(N_1253));
defparam desc1665.INIT=4'hE;
  LUT4 desc1666(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[12:12]),.I2(s_fract_48_i[10:10]),.I3(s_fract_48_i[11:11]),.O(N_704));
defparam desc1666.INIT=16'h000E;
  LUT2 desc1667(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[19:19]),.O(N_1246));
defparam desc1667.INIT=4'hE;
  LUT4 desc1668(.I0(s_fract_48_i[19:19]),.I1(s_fract_48_i[17:17]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[18:18]),.O(N_638));
defparam desc1668.INIT=16'hFFFE;
  LUT2 desc1669(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[18:18]),.O(N_1245));
defparam desc1669.INIT=4'hE;
  LUT4 desc1670(.I0(s_fract_48_i[17:17]),.I1(s_fract_48_i[16:16]),.I2(s_fract_48_i[18:18]),.I3(s_fract_48_i[15:15]),.O(N_464_1));
defparam desc1670.INIT=16'hFFFE;
  LUT2 desc1671(.I0(s_fract_48_i[38:38]),.I1(s_fract_48_i[39:39]),.O(N_591));
defparam desc1671.INIT=4'hE;
  LUT4 desc1672(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[40:40]),.I2(s_fract_48_i[39:39]),.I3(s_fract_48_i[43:43]),.O(N_1249));
defparam desc1672.INIT=16'hFFFE;
  LUT2 desc1673(.I0(s_fract_48_i[32:32]),.I1(s_fract_48_i[33:33]),.O(N_1367));
defparam desc1673.INIT=4'h2;
  LUT4 desc1674(.I0(s_fract_48_i[37:37]),.I1(s_fract_48_i[35:35]),.I2(s_fract_48_i[31:31]),.I3(s_fract_48_i[33:33]),.O(N_1260));
defparam desc1674.INIT=16'hFFFE;
  LUT2 desc1675(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[23:23]),.O(v_count_49_i_o2_0_i_a2_lut6_2_O6[2:2]));
defparam desc1675.INIT=4'h1;
  LUT4 desc1676(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[23:23]),.I3(s_fract_48_i[25:25]),.O(N_1371));
defparam desc1676.INIT=16'h0001;
  LUT2 desc1677(.I0(s_fract_48_i[12:12]),.I1(s_fract_48_i[11:11]),.O(N_434_i_0));
defparam desc1677.INIT=4'h1;
  LUT4 desc1678(.I0(s_fract_48_i[11:11]),.I1(s_fract_48_i[8:8]),.I2(s_fract_48_i[9:9]),.I3(s_fract_48_i[10:10]),.O(N_610));
defparam desc1678.INIT=16'hFFFE;
  LUT2 desc1679(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[21:21]),.O(v_count_49_i_o2_1_i_a2_lut6_2_O6[2:2]));
defparam desc1679.INIT=4'h1;
  LUT4 desc1680(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[20:20]),.I2(s_fract_48_i[21:21]),.I3(s_fract_48_i[19:19]),.O(N_1251));
defparam desc1680.INIT=16'hFFFE;
  LUT2 desc1681(.I0(s_fract_48_i[4:4]),.I1(s_fract_48_i[6:6]),.O(v_count_49_i_o3_i_a2_lut6_2_O6[3:3]));
defparam desc1681.INIT=4'h1;
  LUT5 desc1682(.I0(s_fract_48_i[14:14]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[6:6]),.I3(s_fract_48_i[8:8]),.I4(s_fract_48_i[10:10]),.O(v_count_49_i_o3_i_a2_lut6_2_O5[3:3]));
defparam desc1682.INIT=32'h00000001;
  LUT2 desc1683(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[31:31]),.O(N_37));
defparam desc1683.INIT=4'h1;
  LUT4 desc1684(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[31:31]),.I2(s_fract_48_i[32:32]),.I3(s_fract_48_i[33:33]),.O(N_446));
defparam desc1684.INIT=16'hFFFE;
  LUT2 desc1685(.I0(s_fract_48_i[7:7]),.I1(s_fract_48_i[15:15]),.O(v_count_49_i_a2_0_lut6_2_O6[1:1]));
defparam desc1685.INIT=4'h1;
  LUT5 desc1686(.I0(s_fract_48_i[13:13]),.I1(s_fract_48_i[12:12]),.I2(s_fract_48_i[5:5]),.I3(s_fract_48_i[7:7]),.I4(s_fract_48_i[15:15]),.O(N_677));
defparam desc1686.INIT=32'h00000001;
  LUT2 desc1687(.I0(s_fract_48_i[14:14]),.I1(s_fract_48_i[6:6]),.O(N_672));
defparam desc1687.INIT=4'h1;
  LUT3 desc1688(.I0(s_fract_48_i[14:14]),.I1(s_fract_48_i[4:4]),.I2(s_fract_48_i[6:6]),.O(N_673));
defparam desc1688.INIT=8'h01;
  LUT2 desc1689(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.O(N_582));
defparam desc1689.INIT=4'hE;
  LUT4 desc1690(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[24:24]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[25:25]),.O(N_597));
defparam desc1690.INIT=16'hFFFE;
  LUT2 desc1691(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[7:7]),.O(N_426));
defparam desc1691.INIT=4'hE;
  LUT4 desc1692(.I0(s_fract_48_i[8:8]),.I1(s_fract_48_i[9:9]),.I2(s_fract_48_i[7:7]),.I3(N_1264),.O(N_1350));
defparam desc1692.INIT=16'h2322;
  LUT2 desc1693(.I0(s_fract_48_i[9:9]),.I1(s_fract_48_i[10:10]),.O(N_447));
defparam desc1693.INIT=4'hE;
  LUT4 desc1694(.I0(s_fract_48_i[9:9]),.I1(s_fract_48_i[10:10]),.I2(s_fract_48_i[8:8]),.I3(s_fract_48_i[7:7]),.O(N_449));
defparam desc1694.INIT=16'hFFFE;
  LUT2 desc1695(.I0(s_fract_48_i[28:28]),.I1(s_fract_48_i[29:29]),.O(N_707));
defparam desc1695.INIT=4'h4;
  LUT4 desc1696(.I0(s_fract_48_i[26:26]),.I1(s_fract_48_i[28:28]),.I2(s_fract_48_i[27:27]),.I3(s_fract_48_i[25:25]),.O(N_1361));
defparam desc1696.INIT=16'h0302;
  LUT2 desc1697(.I0(s_exp_10b[6:6]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[6:6]));
defparam desc1697.INIT=4'hE;
  LUT2 desc1698(.I0(s_exp_10b[7:7]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[7:7]));
defparam desc1698.INIT=4'hE;
  LUT2 desc1699(.I0(s_exp_10b[4:4]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[4:4]));
defparam desc1699.INIT=4'hE;
  LUT2 desc1700(.I0(s_exp_10b[5:5]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[5:5]));
defparam desc1700.INIT=4'hE;
  LUT2 desc1701(.I0(s_exp_10b[2:2]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[2:2]));
defparam desc1701.INIT=4'hE;
  LUT2 desc1702(.I0(s_exp_10b[3:3]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[3:3]));
defparam desc1702.INIT=4'hE;
  LUT2 desc1703(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[45:45]),.O(N_592));
defparam desc1703.INIT=4'hE;
  LUT4 desc1704(.I0(s_fract_48_i[45:45]),.I1(s_fract_48_i[39:39]),.I2(s_fract_48_i[41:41]),.I3(s_fract_48_i[43:43]),.O(N_1353));
defparam desc1704.INIT=16'h0001;
  LUT2 desc1705(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[35:35]),.O(N_614));
defparam desc1705.INIT=4'hE;
  LUT2 desc1706(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[32:32]),.O(v_count_0_sqmuxa_47_3_3));
defparam desc1706.INIT=4'h1;
  LUT2 desc1707(.I0(s_fract_48_i[9:9]),.I1(s_fract_48_i[11:11]),.O(N_588));
defparam desc1707.INIT=4'hE;
  LUT5 desc1708(.I0(s_fract_48_i[9:9]),.I1(s_fract_48_i[11:11]),.I2(s_fract_48_i_RNIEUJ9_O5[3:3]),.I3(v_count_49_i_o3_i_a2_lut6_2_O5[3:3]),.I4(N_624),.O(N_668_3));
defparam desc1708.INIT=32'h10000000;
  LUT2 v_count_0_sqmuxa_47_13_lut6_2_o6(.I0(s_fract_48_i[29:29]),.I1(s_fract_48_i[31:31]),.O(N_326_2));
defparam v_count_0_sqmuxa_47_13_lut6_2_o6.INIT=4'h1;
  LUT5 v_count_0_sqmuxa_47_13_lut6_2_o5(.I0(s_fract_48_i[20:20]),.I1(s_fract_48_i[29:29]),.I2(s_fract_48_i[31:31]),.I3(s_fract_48_i[25:25]),.I4(s_fract_48_i[33:33]),.O(v_count_0_sqmuxa_47_2_4));
defparam v_count_0_sqmuxa_47_13_lut6_2_o5.INIT=32'h00000001;
  LUT3 desc1709(.I0(s_fract_48_i[1:1]),.I1(s_fract_48_i[2:2]),.I2(s_shl2[0:0]),.O(N_3));
defparam desc1709.INIT=8'hAC;
  LUT2 desc1710(.I0(s_fract_48_i[3:3]),.I1(s_fract_48_i[2:2]),.O(N_653));
defparam desc1710.INIT=4'h2;
  LUT3 desc1711(.I0(s_fract_48_i[36:36]),.I1(s_fract_48_i[35:35]),.I2(s_shr2[0:0]),.O(N_36));
defparam desc1711.INIT=8'hAC;
  LUT2 desc1712(.I0(s_fract_48_i[37:37]),.I1(s_fract_48_i[35:35]),.O(N_1252));
defparam desc1712.INIT=4'hE;
  LUT3 desc1713(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[45:45]),.I2(s_shr2[0:0]),.O(s_fract_48_i_RNI21942_O6[46:46]));
defparam desc1713.INIT=8'hAC;
  LUT3 desc1714(.I0(s_fract_48_i[44:44]),.I1(s_fract_48_i[45:45]),.I2(s_shl2[0:0]),.O(N_1076));
defparam desc1714.INIT=8'hAC;
  LUT3 desc1715(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[47:47]),.I2(s_shl2[0:0]),.O(N_269));
defparam desc1715.INIT=8'hAC;
  LUT2 desc1716(.I0(s_fract_48_i[46:46]),.I1(s_fract_48_i[47:47]),.O(N_1254));
defparam desc1716.INIT=4'hE;
  LUT3 desc1717(.I0(s_fract_48_i[31:31]),.I1(s_fract_48_i[32:32]),.I2(s_shr2[0:0]),.O(N_40));
defparam desc1717.INIT=8'h35;
  LUT3 desc1718(.I0(s_fract_48_i[41:41]),.I1(s_fract_48_i[42:42]),.I2(s_shr2[0:0]),.O(N_20_0));
defparam desc1718.INIT=8'h35;
  LUT3 desc1719(.I0(s_fract_48_i[23:23]),.I1(s_fract_48_i[27:27]),.I2(s_fract_48_i[29:29]),.O(N_320_0_3));
defparam desc1719.INIT=8'h01;
  LUT2 desc1720(.I0(s_fract_48_i[30:30]),.I1(s_fract_48_i[29:29]),.O(N_173));
defparam desc1720.INIT=4'h1;
  LUT3 desc1721(.I0(s_fract_48_i[31:31]),.I1(s_fract_48_i[32:32]),.I2(s_fract_48_i[33:33]),.O(N_641_1));
defparam desc1721.INIT=8'hBA;
  LUT2 desc1722(.I0(s_fract_48_i[34:34]),.I1(s_fract_48_i[33:33]),.O(N_314_1));
defparam desc1722.INIT=4'hE;
  LUT4 desc1723(.I0(s_fract_48_i[19:19]),.I1(s_fract_48_i[39:39]),.I2(s_fract_48_i[41:41]),.I3(s_fract_48_i[43:43]),.O(v_count_0_sqmuxa_47_1_4));
defparam desc1723.INIT=16'h0001;
  LUT2 desc1724(.I0(s_fract_48_i[41:41]),.I1(s_fract_48_i[42:42]),.O(N_425));
defparam desc1724.INIT=4'hE;
  LUT4 desc1725(.I0(s_fract_48_i[22:22]),.I1(s_fract_48_i[26:26]),.I2(s_fract_48_i[16:16]),.I3(s_fract_48_i[23:23]),.O(v_count_0_sqmuxa_47_4_4));
defparam desc1725.INIT=16'h0001;
  LUT2 desc1726(.I0(s_fract_48_i[16:16]),.I1(s_fract_48_i[15:15]),.O(m107_i_a2_7_0));
defparam desc1726.INIT=4'h1;
  LUT4 un1_s_shr2_1_4_lut6_2_o6(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.O(un1_s_shr2_1_4));
defparam un1_s_shr2_1_4_lut6_2_o6.INIT=16'h0001;
  LUT2 un1_s_shr2_1_4_lut6_2_o5(.I0(s_fract_48_i[47:47]),.I1(s_shr2[0:0]),.O(N_35_0));
defparam un1_s_shr2_1_4_lut6_2_o5.INIT=4'h2;
  LUT3 desc1727(.I0(s_fract_48_i[45:45]),.I1(s_fract_48_i[42:42]),.I2(s_fract_48_i[43:43]),.O(N_1317));
defparam desc1727.INIT=8'h04;
  LUT2 desc1728(.I0(s_fract_48_i[42:42]),.I1(s_fract_48_i[43:43]),.O(s_zeros_2_0_i_a2_3_lut6_2_O5));
defparam desc1728.INIT=4'hE;
  LUT3 desc1729(.I0(s_fract_48_i[4:4]),.I1(s_fract_48_i[5:5]),.I2(s_fract_48_i[2:2]),.O(N_654));
defparam desc1729.INIT=8'h04;
  LUT2 desc1730(.I0(s_fract_48_i[5:5]),.I1(s_fract_48_i[6:6]),.O(N_1255));
defparam desc1730.INIT=4'hE;
  LUT3 un2_s_exp_10a_ac0_1_lut6_2_o6(.I0(s_exp_10_i[1:1]),.I1(s_exp_10_i[0:0]),.I2(s_fract_48_i[47:47]),.O(un2_s_exp_10a_c2));
defparam un2_s_exp_10a_ac0_1_lut6_2_o6.INIT=8'h80;
  LUT5 un2_s_exp_10a_ac0_1_lut6_2_o5(.I0(s_zeros[1:1]),.I1(s_zeros[0:0]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_fract_48_i[47:47]),.O(v_shl1_5_0_0_c2));
defparam un2_s_exp_10a_ac0_1_lut6_2_o5.INIT=32'hFA8E8EAF;
  LUT4 un2_s_exp_10a_ac0_3_lut6_2_o6(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(s_exp_10_i[0:0]),.I3(s_fract_48_i[47:47]),.O(un2_s_exp_10a_c3));
defparam un2_s_exp_10a_ac0_3_lut6_2_o6.INIT=16'h8000;
  LUT4 un2_s_exp_10a_ac0_3_lut6_2_o5(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(s_exp_10_i[0:0]),.I3(s_fract_48_i[47:47]),.O(un5_v_shr1_c3));
defparam un2_s_exp_10a_ac0_3_lut6_2_o5.INIT=16'h9111;
  LUT5 un2_s_lost_ac0_5_lut6_2_o6(.I0(s_frac_rnd[24:24]),.I1(s_shr2[2:2]),.I2(s_shr2[3:3]),.I3(s_shr2[1:1]),.I4(s_shr2[0:0]),.O(un2_s_lost_c4));
defparam un2_s_lost_ac0_5_lut6_2_o6.INIT=32'h80000000;
  LUT4 un2_s_lost_ac0_5_lut6_2_o5(.I0(s_frac_rnd[24:24]),.I1(s_shr2[2:2]),.I2(s_shr2[1:1]),.I3(s_shr2[0:0]),.O(un2_s_lost_ac0_5_lut6_2_O5));
defparam un2_s_lost_ac0_5_lut6_2_o5.INIT=16'h6CCC;
  LUT3 desc1731(.I0(s_shl2[2:2]),.I1(N_85_0),.I2(s_frac2a_2_91),.O(N_137));
defparam desc1731.INIT=8'hD8;
  LUT3 desc1732(.I0(s_shl2[2:2]),.I1(N_86),.I2(N_49),.O(N_1157));
defparam desc1732.INIT=8'h72;
  LUT3 desc1733(.I0(s_shl2[2:2]),.I1(N_61),.I2(N_57),.O(N_109));
defparam desc1733.INIT=8'hE4;
  LUT3 desc1734(.I0(s_shl2[2:2]),.I1(N_67),.I2(N_63),.O(N_115));
defparam desc1734.INIT=8'hE4;
  LUT3 desc1735(.I0(s_shl2[2:2]),.I1(N_64),.I2(N_60),.O(s_frac2a_2_115_lut6_2_O6));
defparam desc1735.INIT=8'hE4;
  LUT3 desc1736(.I0(s_shl2[2:2]),.I1(N_63),.I2(N_59),.O(N_111));
defparam desc1736.INIT=8'hE4;
  LUT3 desc1737(.I0(s_shl2[2:2]),.I1(N_62),.I2(N_58),.O(N_110));
defparam desc1737.INIT=8'hE4;
  LUT3 desc1738(.I0(s_shl2[2:2]),.I1(N_81),.I2(N_77),.O(N_129));
defparam desc1738.INIT=8'hE4;
  LUT3 desc1739(.I0(s_shl2[2:2]),.I1(N_54),.I2(N_58),.O(N_106));
defparam desc1739.INIT=8'hD8;
  LUT3 desc1740(.I0(s_shl2[2:2]),.I1(N_73),.I2(N_69),.O(N_121));
defparam desc1740.INIT=8'hE4;
  LUT3 desc1741(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_905),.O(N_214));
defparam desc1741.INIT=8'h01;
  LUT3 desc1742(.I0(s_shr2[2:2]),.I1(N_51),.I2(N_55),.O(N_99));
defparam desc1742.INIT=8'hE4;
  LUT4 desc1743(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_78),.I3(N_74),.O(N_1140));
defparam desc1743.INIT=16'h3210;
  LUT4 desc1744(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_74),.I3(N_70),.O(N_370));
defparam desc1744.INIT=16'h3210;
  LUT4 desc1745(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_50),.I3(N_54),.O(N_1096));
defparam desc1745.INIT=16'h3120;
  LUT4 desc1746(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_54),.I3(N_58),.O(N_361));
defparam desc1746.INIT=16'h3120;
  LUT4 desc1747(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_62),.I3(N_58),.O(N_1094));
defparam desc1747.INIT=16'h3210;
  LUT4 desc1748(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_62),.I3(N_66),.O(N_360));
defparam desc1748.INIT=16'h3120;
  LUT4 desc1749(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_52),.I3(N_56),.O(N_1086));
defparam desc1749.INIT=16'h3120;
  LUT4 desc1750(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_56),.I3(N_60),.O(N_280));
defparam desc1750.INIT=16'h3120;
  LUT4 desc1751(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_64),.I3(N_60),.O(N_1085));
defparam desc1751.INIT=16'h3210;
  LUT4 desc1752(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_68),.I3(N_64),.O(N_289));
defparam desc1752.INIT=16'h3210;
  LUT4 desc1753(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_72),.I3(N_68),.O(N_1084));
defparam desc1753.INIT=16'h3210;
  LUT3 desc1754(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_52),.O(N_265));
defparam desc1754.INIT=8'h10;
  LUT4 desc1755(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_80),.I3(N_76),.O(N_25_0));
defparam desc1755.INIT=16'h3210;
  LUT4 desc1756(.I0(s_shl2[2:2]),.I1(s_shl2[5:5]),.I2(N_72),.I3(N_76),.O(N_297));
defparam desc1756.INIT=16'h3120;
  LUT3 desc1757(.I0(s_shr2[3:3]),.I1(s_frac2a_1_132),.I2(N_138),.O(N_337));
defparam desc1757.INIT=8'hE4;
  LUT5 desc1758(.I0(s_shr2[3:3]),.I1(un1_s_shr2_1_4),.I2(s_frac2a_1_132),.I3(N_138),.I4(N_1156),.O(N_396));
defparam desc1758.INIT=32'hFEDC3210;
  LUT5 desc1759(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_85),.I3(N_905),.I4(N_904),.O(N_223));
defparam desc1759.INIT=32'h10543276;
  LUT4 desc1760(.I0(s_shr2[2:2]),.I1(s_shr2[3:3]),.I2(N_905),.I3(N_904),.O(N_1165));
defparam desc1760.INIT=16'h0213;
  LUT3 desc1761(.I0(s_shr2[3:3]),.I1(N_126),.I2(N_134),.O(s_frac2a_1_124_RNIEJB51_O6));
defparam desc1761.INIT=8'h1B;
  LUT3 desc1762(.I0(s_shr2[3:3]),.I1(s_frac2a_1_132),.I2(s_frac2a_1_124),.O(N_355));
defparam desc1762.INIT=8'hD8;
  LUT3 desc1763(.I0(s_shl2[3:3]),.I1(N_1120),.I2(N_1114),.O(N_1121));
defparam desc1763.INIT=8'hE4;
  LUT3 desc1764(.I0(s_shl2[3:3]),.I1(N_240),.I2(N_242),.O(N_243));
defparam desc1764.INIT=8'hB1;
  LUT5 desc1765(.I0(N_368),.I1(s_shl2[4:4]),.I2(s_shl2[3:3]),.I3(s_shl2[5:5]),.I4(N_1078),.O(m368_lut6_2_O6));
defparam desc1765.INIT=32'h222E2222;
  LUT4 desc1766(.I0(s_shl2[4:4]),.I1(s_shl2[3:3]),.I2(s_shl2[5:5]),.I3(N_1078),.O(N_1081));
defparam desc1766.INIT=16'h0100;
  LUT3 s_exp_10b_s_1_RNI0PGD1_o6(.I0(s_exp_10b[9:9]),.I1(un6_s_exp_10a),.I2(s_exp_10b[8:8]),.O(s_exp_10b_s_1_RNI0PGD1_O6));
defparam s_exp_10b_s_1_RNI0PGD1_o6.INIT=8'hDC;
  LUT2 s_exp_10b_s_1_RNI0PGD1_o5(.I0(s_exp_10b[1:1]),.I1(s_exp_10b[8:8]),.O(s_expo1_5[1:1]));
defparam s_exp_10b_s_1_RNI0PGD1_o5.INIT=4'hE;
  LUT2 un1_s_exp_10a_3_lut6_2_o6(.I0(un6_s_exp_10a),.I1(un1_s_exp_10a_3_1),.O(un1_s_exp_10a_3_lut6_2_O6));
defparam un1_s_exp_10a_3_lut6_2_o6.INIT=4'hE;
  LUT3 un1_s_exp_10a_3_lut6_2_o5(.I0(s_exp_10_i[1:1]),.I1(un6_s_exp_10a),.I2(v_shr1_4[6:6]),.O(v_shr1_4_e[1:1]));
defparam un1_s_exp_10a_3_lut6_2_o5.INIT=8'hF8;
  LUT2 desc1767(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.O(N_459_i));
defparam desc1767.INIT=4'hE;
  LUT5 desc1768(.I0(s_shr2[5:5]),.I1(s_shr2[4:4]),.I2(N_82_0),.I3(N_80_0),.I4(N_79_0),.O(s_frac2a_3[14:14]));
defparam desc1768.INIT=32'h31752064;
  LUT3 desc1769(.I0(s_frac2a[46:46]),.I1(s_frac_rnd_3_0_s_23),.I2(s_roundup),.O(s_frac_rnd_3[23:23]));
defparam desc1769.INIT=8'hCA;
  LUT3 desc1770(.I0(s_frac2a[47:47]),.I1(s_frac_rnd_3_0_s_24),.I2(s_roundup),.O(s_frac_rnd_3[24:24]));
defparam desc1770.INIT=8'hCA;
  LUT3 desc1771(.I0(s_frac2a[44:44]),.I1(s_frac_rnd_3_0_s_21),.I2(s_roundup),.O(s_frac_rnd_3[21:21]));
defparam desc1771.INIT=8'hCA;
  LUT3 desc1772(.I0(s_frac2a[45:45]),.I1(s_frac_rnd_3_0_s_22),.I2(s_roundup),.O(s_frac_rnd_3[22:22]));
defparam desc1772.INIT=8'hCA;
  LUT3 desc1773(.I0(s_frac2a[42:42]),.I1(s_frac_rnd_3_0_s_19),.I2(s_roundup),.O(s_frac_rnd_3[19:19]));
defparam desc1773.INIT=8'hCA;
  LUT3 desc1774(.I0(s_frac2a[43:43]),.I1(s_frac_rnd_3_0_s_20),.I2(s_roundup),.O(s_frac_rnd_3[20:20]));
defparam desc1774.INIT=8'hCA;
  LUT3 desc1775(.I0(s_frac2a[40:40]),.I1(s_frac_rnd_3_0_s_17),.I2(s_roundup),.O(s_frac_rnd_3[17:17]));
defparam desc1775.INIT=8'hCA;
  LUT3 desc1776(.I0(s_frac2a[41:41]),.I1(s_frac_rnd_3_0_s_18),.I2(s_roundup),.O(s_frac_rnd_3[18:18]));
defparam desc1776.INIT=8'hCA;
  LUT3 desc1777(.I0(s_frac2a[37:37]),.I1(s_frac_rnd_3_0_s_14),.I2(s_roundup),.O(s_frac_rnd_3[14:14]));
defparam desc1777.INIT=8'hCA;
  LUT3 desc1778(.I0(s_frac2a[38:38]),.I1(s_frac_rnd_3_0_s_15),.I2(s_roundup),.O(s_frac_rnd_3[15:15]));
defparam desc1778.INIT=8'hCA;
  LUT3 desc1779(.I0(s_frac2a[35:35]),.I1(s_frac_rnd_3_0_s_12),.I2(s_roundup),.O(s_frac_rnd_3[12:12]));
defparam desc1779.INIT=8'hCA;
  LUT3 desc1780(.I0(s_frac2a[36:36]),.I1(s_frac_rnd_3_0_s_13),.I2(s_roundup),.O(s_frac_rnd_3[13:13]));
defparam desc1780.INIT=8'hCA;
  LUT3 desc1781(.I0(s_frac2a[33:33]),.I1(s_frac_rnd_3_0_s_10),.I2(s_roundup),.O(s_frac_rnd_3[10:10]));
defparam desc1781.INIT=8'hCA;
  LUT3 desc1782(.I0(s_frac2a[34:34]),.I1(s_frac_rnd_3_0_s_11),.I2(s_roundup),.O(s_frac_rnd_3[11:11]));
defparam desc1782.INIT=8'hCA;
  LUT3 desc1783(.I0(s_frac2a[31:31]),.I1(s_frac_rnd_3_0_s_8),.I2(s_roundup),.O(s_frac_rnd_3[8:8]));
defparam desc1783.INIT=8'hCA;
  LUT3 desc1784(.I0(s_frac2a[32:32]),.I1(s_frac_rnd_3_0_s_9),.I2(s_roundup),.O(s_frac_rnd_3[9:9]));
defparam desc1784.INIT=8'hCA;
  LUT3 desc1785(.I0(s_frac2a[29:29]),.I1(s_frac_rnd_3_0_s_6),.I2(s_roundup),.O(s_frac_rnd_3[6:6]));
defparam desc1785.INIT=8'hCA;
  LUT3 desc1786(.I0(s_frac2a[30:30]),.I1(s_frac_rnd_3_0_s_7),.I2(s_roundup),.O(s_frac_rnd_3[7:7]));
defparam desc1786.INIT=8'hCA;
  LUT3 desc1787(.I0(s_frac2a[27:27]),.I1(s_frac_rnd_3_0_s_4),.I2(s_roundup),.O(s_frac_rnd_3[4:4]));
defparam desc1787.INIT=8'hCA;
  LUT3 desc1788(.I0(s_frac2a[28:28]),.I1(s_frac_rnd_3_0_s_5),.I2(s_roundup),.O(s_frac_rnd_3[5:5]));
defparam desc1788.INIT=8'hCA;
  LUT3 desc1789(.I0(s_frac2a[25:25]),.I1(s_frac_rnd_3_0_s_2),.I2(s_roundup),.O(s_frac_rnd_3[2:2]));
defparam desc1789.INIT=8'hCA;
  LUT3 desc1790(.I0(s_frac2a[26:26]),.I1(s_frac_rnd_3_0_s_3),.I2(s_roundup),.O(s_frac_rnd_3[3:3]));
defparam desc1790.INIT=8'hCA;
  LUT3 desc1791(.I0(s_frac2a[24:24]),.I1(s_frac_rnd_3_0_s_1),.I2(s_roundup),.O(s_frac_rnd_3[1:1]));
defparam desc1791.INIT=8'hCA;
  LUT2 desc1792(.I0(s_frac2a[23:23]),.I1(s_roundup),.O(s_frac_rnd_3[0:0]));
defparam desc1792.INIT=4'h6;
  LUT3 desc1793(.I0(s_zeros[0:0]),.I1(s_exp_10_i[0:0]),.I2(s_fract_48_i[47:47]),.O(s_exp_10b_i));
defparam desc1793.INIT=8'h69;
  LUT2 desc1794(.I0(s_exp_10_i[0:0]),.I1(s_fract_48_i[47:47]),.O(s_zeros_RNI0TNS_O5));
defparam desc1794.INIT=4'h6;
endmodule
module pre_norm_div_inj (v_count_3,v_count_2,v_count_1_0_0_a2_0,v_count_2_0,s_exp_10_o_0,s_exp_10_o,pre_norm_div_dvsor_0,v_count_1_0_1,v_count_1_0_2,v_count_0_4,v_count_0_1,v_count_0_0,v_count_i,s_opb_i,s_opb_i_0_0,s_opb_i_0_3,s_opb_i_0_4,s_opb_i_0_2,s_opb_i_0_5,s_opa_i_0,s_opa_i,v_count_1_0_a2_7_i_0,pre_norm_div_dvsor,pre_norm_div_dvdnd_0,pre_norm_div_dvdnd_11,un11_s_exp_10_o_0,N_1083,N_143_mux,N_48_0,N_59,N_54,N_1630,N_55,N_63,N_1278_i,s_dvdnd_50_o_105_0_e,N_987,s_expa_lt_expb,N_2240,N_1232_i,un2_s_snan_o_22,N_1174,result_i_o3_lut6_2_O6,result_3_0_0_i,N_1055,N_1077,N_399,un4_s_infa_1,N_1140,N_1051,N_2220,N_1170,un4_s_expb_in_2_i_o2_2,un4_s_expb_in_2_i_o2_2_lut6_2_O5,N_1041,result_2_16,s_dvdnd_50_o_104_0_e,un4_s_expb_in_2_i_0_e,clk_i,s_dvdnd_50_o_103_0_e,s_dvdnd_50_o_102_0_e,s_dvdnd_50_o_106_0_e,s_dvdnd_50_o_108_0_e,N_1236,N_2103,s_dvdnd_50_o_107_0_e,un4_s_expb_in_2_i_o2_0,un4_s_expb_in_2_i_o2_1,result_1_i_o3_0_e,N_1227,N_378_i,N_396,result_1_i_o3,N_1084_i,un11_s_exp_10_o_axb_0_i,N_1050,N_1087,un2_s_snan_o_8,result_2_10,N_1617,N_41_0,N_43_0,N_44,N_45_0,N_1628,N_1624,N_1619,N_46,N_1620,N_95_0,N_70_0,N_27_0,N_1238);
input v_count_3 ;
input v_count_2 ;
output [1:1] v_count_1_0_0_a2_0 ;
output [4:4] v_count_2_0 ;
input [1:0] s_exp_10_o_0 ;
output [1:1] s_exp_10_o ;
output [23:23] pre_norm_div_dvsor_0 ;
output v_count_1_0_1 ;
output v_count_1_0_2 ;
output v_count_0_4 ;
input v_count_0_1 ;
output v_count_0_0 ;
output v_count_i ;
input [30:0] s_opb_i ;
input s_opb_i_0_0 ;
input s_opb_i_0_3 ;
input s_opb_i_0_4 ;
input s_opb_i_0_2 ;
input s_opb_i_0_5 ;
input [30:24] s_opa_i_0 ;
input [30:0] s_opa_i ;
input v_count_1_0_a2_7_i_0 ;
output [22:7] pre_norm_div_dvsor ;
output pre_norm_div_dvdnd_0 ;
output pre_norm_div_dvdnd_11 ;
output [9:1] un11_s_exp_10_o_0 ;
output N_1083 ;
input N_143_mux ;
input N_48_0 ;
output N_59 ;
output N_54 ;
output N_1630 ;
output N_55 ;
output N_63 ;
output N_1278_i ;
output s_dvdnd_50_o_105_0_e ;
input N_987 ;
input s_expa_lt_expb ;
input N_2240 ;
output N_1232_i ;
output un2_s_snan_o_22 ;
input N_1174 ;
output result_i_o3_lut6_2_O6 ;
output result_3_0_0_i ;
output N_1055 ;
output N_1077 ;
output N_399 ;
output un4_s_infa_1 ;
output N_1140 ;
input N_1051 ;
output N_2220 ;
output N_1170 ;
output un4_s_expb_in_2_i_o2_2 ;
output un4_s_expb_in_2_i_o2_2_lut6_2_O5 ;
output N_1041 ;
output result_2_16 ;
output s_dvdnd_50_o_104_0_e ;
input un4_s_expb_in_2_i_0_e ;
input clk_i ;
output s_dvdnd_50_o_103_0_e ;
output s_dvdnd_50_o_102_0_e ;
output s_dvdnd_50_o_106_0_e ;
output s_dvdnd_50_o_108_0_e ;
input N_1236 ;
output N_2103 ;
output s_dvdnd_50_o_107_0_e ;
input un4_s_expb_in_2_i_o2_0 ;
output un4_s_expb_in_2_i_o2_1 ;
output result_1_i_o3_0_e ;
output N_1227 ;
input N_378_i ;
output N_396 ;
output result_1_i_o3 ;
output N_1084_i ;
output un11_s_exp_10_o_axb_0_i ;
input N_1050 ;
input N_1087 ;
input un2_s_snan_o_8 ;
input result_2_10 ;
output N_1617 ;
output N_41_0 ;
output N_43_0 ;
output N_44 ;
output N_45_0 ;
output N_1628 ;
output N_1624 ;
output N_1619 ;
output N_46 ;
output N_1620 ;
output N_95_0 ;
input N_70_0 ;
input N_27_0 ;
input N_1238 ;
wire v_count_3 ;
wire v_count_2 ;
wire v_count_0_4 ;
wire v_count_0_1 ;
wire v_count_0_0 ;
wire s_opb_i_0_0 ;
wire s_opb_i_0_3 ;
wire s_opb_i_0_4 ;
wire s_opb_i_0_2 ;
wire s_opb_i_0_5 ;
wire pre_norm_div_dvdnd_0 ;
wire pre_norm_div_dvdnd_11 ;
wire N_1083 ;
wire N_143_mux ;
wire N_48_0 ;
wire N_59 ;
wire N_54 ;
wire N_1630 ;
wire N_55 ;
wire N_63 ;
wire N_1278_i ;
wire s_dvdnd_50_o_105_0_e ;
wire N_987 ;
wire s_expa_lt_expb ;
wire N_2240 ;
wire N_1232_i ;
wire un2_s_snan_o_22 ;
wire N_1174 ;
wire result_i_o3_lut6_2_O6 ;
wire result_3_0_0_i ;
wire N_1055 ;
wire N_1077 ;
wire N_399 ;
wire un4_s_infa_1 ;
wire N_1140 ;
wire N_1051 ;
wire N_2220 ;
wire N_1170 ;
wire un4_s_expb_in_2_i_o2_2 ;
wire un4_s_expb_in_2_i_o2_2_lut6_2_O5 ;
wire N_1041 ;
wire result_2_16 ;
wire s_dvdnd_50_o_104_0_e ;
wire un4_s_expb_in_2_i_0_e ;
wire clk_i ;
wire s_dvdnd_50_o_103_0_e ;
wire s_dvdnd_50_o_102_0_e ;
wire s_dvdnd_50_o_106_0_e ;
wire s_dvdnd_50_o_108_0_e ;
wire N_1236 ;
wire N_2103 ;
wire s_dvdnd_50_o_107_0_e ;
wire un4_s_expb_in_2_i_o2_0 ;
wire un4_s_expb_in_2_i_o2_1 ;
wire result_1_i_o3_0_e ;
wire N_1227 ;
wire N_378_i ;
wire N_396 ;
wire result_1_i_o3 ;
wire N_1084_i ;
wire un11_s_exp_10_o_axb_0_i ;
wire N_1050 ;
wire N_1087 ;
wire un2_s_snan_o_8 ;
wire result_2_10 ;
wire N_1617 ;
wire N_41_0 ;
wire N_43_0 ;
wire N_44 ;
wire N_45_0 ;
wire N_1628 ;
wire N_1624 ;
wire N_1619 ;
wire N_46 ;
wire N_1620 ;
wire N_95_0 ;
wire N_70_0 ;
wire N_27_0 ;
wire N_1238 ;
wire [9:0] un11_s_exp_10_o_5 ;
wire [4:0] v_count ;
wire [3:2] v_count_0 ;
wire v_count_1_0_a2_0 ;
wire s_expb_in ;
wire s_expa_in ;
wire [8:0] un11_s_exp_10_o_6 ;
wire [8:5] un11_s_exp_10_o_6_i ;
wire [8:8] un11_s_exp_10_o_6_1 ;
wire [8:8] un11_s_exp_10_o_6_0 ;
wire v_count_1_0_a2_1_4 ;
wire [2:2] v_count_0_0_a5_0_1_1 ;
wire GND ;
wire un11_s_exp_10_o_5_s_9_true ;
wire VCC ;
wire un11_s_exp_10_o_axb_0 ;
wire N_1622 ;
wire N_1626 ;
wire N_64 ;
wire N_62 ;
wire N_56 ;
wire N_112 ;
wire N_101 ;
wire N_76 ;
wire N_1049 ;
wire N_1219 ;
wire N_340 ;
wire N_432 ;
wire N_240_2 ;
wire N_1052 ;
wire N_304_1 ;
wire result_2_11 ;
wire N_22 ;
wire N_1216 ;
wire N_27 ;
wire N_91 ;
wire N_121 ;
wire N_25 ;
wire N_124 ;
wire un11_s_exp_10_o_6_axb_1 ;
wire un11_s_exp_10_o_6_axb_2 ;
wire un11_s_exp_10_o_6_axb_3 ;
wire un11_s_exp_10_o_6_axb_4 ;
wire un11_s_exp_10_o_6_axb_5 ;
wire un11_s_exp_10_o_6_axb_6 ;
wire un11_s_exp_10_o_6_axb_7 ;
wire un11_s_exp_10_o_5_axb_2 ;
wire un11_s_exp_10_o_5_axb_3 ;
wire un11_s_exp_10_o_5_axb_4 ;
wire un11_s_exp_10_o_5_axb_7 ;
wire N_89 ;
wire N_93 ;
wire N_95 ;
wire N_296 ;
wire N_341 ;
wire N_384 ;
wire un11_s_exp_10_o_axb_3 ;
wire un11_s_exp_10_o_axb_4 ;
wire N_104 ;
wire N_108 ;
wire N_100 ;
wire N_2194 ;
wire N_110 ;
wire N_106 ;
wire N_20 ;
wire N_18 ;
wire result_i_o2_0_0 ;
wire un11_s_exp_10_o_axb_9 ;
wire un11_s_exp_10_o_axb_8 ;
wire un11_s_exp_10_o_axb_7 ;
wire un11_s_exp_10_o_axb_6 ;
wire un11_s_exp_10_o_axb_5 ;
wire N_290 ;
wire N_1160 ;
wire N_238 ;
wire un11_s_exp_10_o_axb_2 ;
wire un11_s_exp_10_o_axb_1 ;
wire un11_s_exp_10_o_5_axb_1 ;
wire N_126 ;
wire N_128 ;
wire N_130 ;
wire N_132 ;
wire N_41 ;
wire N_43 ;
wire N_45 ;
wire N_47 ;
wire N_47_0 ;
wire N_58 ;
wire N_60 ;
wire N_66 ;
wire N_68 ;
wire N_70 ;
wire N_74 ;
wire un11_s_exp_10_o_cry_8 ;
wire un11_s_exp_10_o_cry_7 ;
wire un11_s_exp_10_o_cry_6 ;
wire un11_s_exp_10_o_cry_5 ;
wire un11_s_exp_10_o_cry_4 ;
wire un11_s_exp_10_o_cry_3 ;
wire un11_s_exp_10_o_cry_2 ;
wire un11_s_exp_10_o_cry_1 ;
wire un11_s_exp_10_o_cry_0 ;
wire un11_s_exp_10_o_5_cry_8 ;
wire un11_s_exp_10_o_5_cry_7 ;
wire un11_s_exp_10_o_5_cry_6 ;
wire un11_s_exp_10_o_5_cry_5 ;
wire un11_s_exp_10_o_5_cry_4 ;
wire un11_s_exp_10_o_5_cry_3 ;
wire un11_s_exp_10_o_5_cry_2 ;
wire un11_s_exp_10_o_5_cry_1 ;
wire un11_s_exp_10_o_5_cry_0 ;
wire un11_s_exp_10_o_6_cry_6 ;
wire un11_s_exp_10_o_6_cry_5 ;
wire un11_s_exp_10_o_6_cry_4 ;
wire un11_s_exp_10_o_6_cry_3 ;
wire un11_s_exp_10_o_6_cry_2 ;
wire un11_s_exp_10_o_6_cry_1 ;
wire un11_s_exp_10_o_6_cry_0 ;
// instances
  LUT1 un11_s_exp_10_o_5_s_9_true_cZ(.I0(GND),.O(un11_s_exp_10_o_5_s_9_true));
defparam un11_s_exp_10_o_5_s_9_true_cZ.INIT=2'h3;
  LUT6_2 desc1795(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(v_count_0[3:3]),.I3(N_112),.I4(N_101),.I5(v_count[4:4]),.O6(s_dvdnd_50_o_105_0_e),.O5(N_76));
defparam desc1795.INIT=64'h0000000005040100;
  LUT6_2 desc1796(.I0(s_opa_i[21:21]),.I1(s_opa_i[22:22]),.I2(s_opa_i[20:20]),.I3(un2_s_snan_o_22),.I4(N_1174),.I5(result_i_o3_lut6_2_O6),.O6(v_count_0_4),.O5(result_3_0_0_i));
defparam desc1796.INIT=64'h0000000000000100;
  FD desc1797(.Q(s_expb_in),.D(un4_s_expb_in_2_i_0_e),.C(clk_i));
  LUT5 desc1798(.I0(N_101),.I1(v_count[1:1]),.I2(v_count_0[2:2]),.I3(v_count_0[3:3]),.I4(v_count[4:4]),.O(s_dvdnd_50_o_103_0_e));
defparam desc1798.INIT=32'h00000002;
  LUT6 desc1799(.I0(v_count[0:0]),.I1(v_count[1:1]),.I2(v_count_0[2:2]),.I3(v_count_0[3:3]),.I4(s_opb_i[0:0]),.I5(v_count[4:4]),.O(s_dvdnd_50_o_102_0_e));
defparam desc1799.INIT=64'h0000000000010000;
  LUT5 desc1800(.I0(N_121),.I1(N_25),.I2(v_count_0[2:2]),.I3(v_count_0[3:3]),.I4(v_count[4:4]),.O(s_dvdnd_50_o_106_0_e));
defparam desc1800.INIT=32'h000000CA;
  LUT5 desc1801(.I0(N_124),.I1(N_27),.I2(v_count_0[2:2]),.I3(v_count_0[3:3]),.I4(v_count[4:4]),.O(s_dvdnd_50_o_108_0_e));
defparam desc1801.INIT=32'h000000CA;
  LUT6 desc1802(.I0(N_1236),.I1(N_2103),.I2(v_count_0_1),.I3(v_count_2),.I4(v_count_3),.I5(v_count_0_4),.O(s_dvdnd_50_o_107_0_e));
defparam desc1802.INIT=64'h0000000000000C55;
  LUT6 un4_s_expb_in_2_i_o2_1_RNI3K4D2(.I0(un4_s_expb_in_2_i_o2_0),.I1(un4_s_expb_in_2_i_o2_1),.I2(s_opb_i[24:24]),.I3(s_opb_i[27:27]),.I4(s_opb_i[28:28]),.I5(s_opb_i[23:23]),.O(result_1_i_o3_0_e));
defparam un4_s_expb_in_2_i_o2_1_RNI3K4D2.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT2 un11_s_exp_10_o_6_axb_0(.I0(s_expa_in),.I1(s_expb_in),.O(un11_s_exp_10_o_6[0:0]));
defparam un11_s_exp_10_o_6_axb_0.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_1_cZ(.I0(s_opa_i_0[24:24]),.I1(s_opb_i_0_0),.O(un11_s_exp_10_o_6_axb_1));
defparam un11_s_exp_10_o_6_axb_1_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_2_cZ(.I0(s_opa_i[25:25]),.I1(s_opb_i[25:25]),.O(un11_s_exp_10_o_6_axb_2));
defparam un11_s_exp_10_o_6_axb_2_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_3_cZ(.I0(s_opa_i_0[26:26]),.I1(s_opb_i[26:26]),.O(un11_s_exp_10_o_6_axb_3));
defparam un11_s_exp_10_o_6_axb_3_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_4_cZ(.I0(s_opa_i_0[27:27]),.I1(s_opb_i_0_3),.O(un11_s_exp_10_o_6_axb_4));
defparam un11_s_exp_10_o_6_axb_4_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_5_cZ(.I0(s_opa_i[28:28]),.I1(s_opb_i_0_4),.O(un11_s_exp_10_o_6_axb_5));
defparam un11_s_exp_10_o_6_axb_5_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_6_cZ(.I0(s_opa_i[29:29]),.I1(s_opb_i[29:29]),.O(un11_s_exp_10_o_6_axb_6));
defparam un11_s_exp_10_o_6_axb_6_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_6_axb_7_cZ(.I0(s_opa_i_0[30:30]),.I1(s_opb_i[30:30]),.O(un11_s_exp_10_o_6_axb_7));
defparam un11_s_exp_10_o_6_axb_7_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_5_axb_2_cZ(.I0(un11_s_exp_10_o_6[2:2]),.I1(v_count_2),.O(un11_s_exp_10_o_5_axb_2));
defparam un11_s_exp_10_o_5_axb_2_cZ.INIT=4'h9;
  LUT2 un11_s_exp_10_o_5_axb_3_cZ(.I0(un11_s_exp_10_o_6[3:3]),.I1(v_count_3),.O(un11_s_exp_10_o_5_axb_3));
defparam un11_s_exp_10_o_5_axb_3_cZ.INIT=4'h9;
  LUT3 un11_s_exp_10_o_5_axb_4_cZ(.I0(N_1174),.I1(N_1227),.I2(un11_s_exp_10_o_6[4:4]),.O(un11_s_exp_10_o_5_axb_4));
defparam un11_s_exp_10_o_5_axb_4_cZ.INIT=8'h4B;
  LUT1 desc1803(.I0(un11_s_exp_10_o_6[5:5]),.O(un11_s_exp_10_o_6_i[5:5]));
defparam desc1803.INIT=2'h1;
  LUT1 desc1804(.I0(un11_s_exp_10_o_6[6:6]),.O(un11_s_exp_10_o_6_i[6:6]));
defparam desc1804.INIT=2'h1;
  LUT1 un11_s_exp_10_o_5_axb_7_cZ(.I0(un11_s_exp_10_o_6[7:7]),.O(un11_s_exp_10_o_5_axb_7));
defparam un11_s_exp_10_o_5_axb_7_cZ.INIT=2'h2;
  LUT1 desc1805(.I0(un11_s_exp_10_o_6[8:8]),.O(un11_s_exp_10_o_6_i[8:8]));
defparam desc1805.INIT=2'h1;
  LUT1 un11_s_exp_10_o_6_cry_7_outextlut(.I0(GND),.O(un11_s_exp_10_o_6_1[8:8]));
defparam un11_s_exp_10_o_6_cry_7_outextlut.INIT=2'h3;
  FD desc1806(.Q(s_expa_in),.D(N_378_i),.C(clk_i));
  MUXCY un11_s_exp_10_o_6_cry_7_outext(.DI(GND),.CI(un11_s_exp_10_o_6_0[8:8]),.S(un11_s_exp_10_o_6_1[8:8]),.O(un11_s_exp_10_o_6[8:8]));
  LUT4_L desc1807(.I0(v_count_0[2:2]),.I1(v_count[4:4]),.I2(N_25),.I3(N_89),.LO(pre_norm_div_dvsor[16:16]));
defparam desc1807.INIT=16'h3340;
  LUT5_L desc1808(.I0(v_count_0[2:2]),.I1(v_count[4:4]),.I2(N_25),.I3(N_121),.I4(N_93),.LO(pre_norm_div_dvsor[20:20]));
defparam desc1808.INIT=32'h33334480;
  LUT5_L desc1809(.I0(v_count_0[2:2]),.I1(v_count[4:4]),.I2(N_124),.I3(N_27),.I4(N_95),.LO(pre_norm_div_dvsor[22:22]));
defparam desc1809.INIT=32'h33334840;
  LUT6 desc1810(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[12:12]),.I4(N_1041),.I5(N_296),.O(N_341));
defparam desc1810.INIT=64'h0303030203020302;
  LUT6 desc1811(.I0(s_expb_in),.I1(s_expa_in),.I2(N_399),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(un11_s_exp_10_o_5[0:0]));
defparam desc1811.INIT=64'h9999999999999996;
  LUT6 desc1812(.I0(s_opa_i[13:13]),.I1(s_opa_i[15:15]),.I2(s_opa_i[11:11]),.I3(s_opa_i[9:9]),.I4(N_384),.I5(N_240_2),.O(v_count_1_0_a2_1_4));
defparam desc1812.INIT=64'h0001000000000000;
  LUT6 desc1813(.I0(s_opb_i[14:14]),.I1(s_opb_i[15:15]),.I2(s_opb_i[8:8]),.I3(s_opb_i[9:9]),.I4(N_1049),.I5(N_1041),.O(N_1055));
defparam desc1813.INIT=64'h0001000000000000;
  LUT6 desc1814(.I0(s_opb_i[24:24]),.I1(s_opb_i[28:28]),.I2(s_opb_i[27:27]),.I3(s_opb_i[23:23]),.I4(un4_s_expb_in_2_i_o2_0),.I5(un4_s_expb_in_2_i_o2_1),.O(result_1_i_o3));
defparam desc1814.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 un4_s_expb_in_2_i_o2_1_RNI3K4D2_0(.I0(s_opb_i[24:24]),.I1(s_opb_i[28:28]),.I2(s_opb_i[27:27]),.I3(s_opb_i[23:23]),.I4(un4_s_expb_in_2_i_o2_0),.I5(un4_s_expb_in_2_i_o2_1),.O(N_1084_i));
defparam un4_s_expb_in_2_i_o2_1_RNI3K4D2_0.INIT=64'h0000000000000001;
  LUT6 desc1815(.I0(s_opa_i[22:22]),.I1(s_opa_i[24:24]),.I2(N_1077),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(v_count_0_0));
defparam desc1815.INIT=64'hFFFFFFFFFFFFFF02;
  LUT6 desc1816(.I0(s_opa_i[22:22]),.I1(s_opa_i[24:24]),.I2(N_1077),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(v_count_i));
defparam desc1816.INIT=64'h00000000000000FD;
  LUT6 un11_s_exp_10_o_axb_3_cZ(.I0(s_opb_i[16:16]),.I1(s_opb_i[18:18]),.I2(N_340),.I3(N_1055),.I4(v_count_2_0[4:4]),.I5(un11_s_exp_10_o_5[3:3]),.O(un11_s_exp_10_o_axb_3));
defparam un11_s_exp_10_o_axb_3_cZ.INIT=64'hEFEEFFFF10110000;
  LUT5 un11_s_exp_10_o_axb_4_cZ(.I0(s_opb_i[16:16]),.I1(s_opb_i[18:18]),.I2(N_1055),.I3(v_count_2_0[4:4]),.I4(un11_s_exp_10_o_5[4:4]),.O(un11_s_exp_10_o_axb_4));
defparam un11_s_exp_10_o_axb_4_cZ.INIT=32'hEFFF1000;
  LUT6 desc1817(.I0(s_opb_i[0:0]),.I1(s_opb_i[22:22]),.I2(s_opb_i[23:23]),.I3(N_1083),.I4(N_143_mux),.I5(v_count[1:1]),.O(N_25));
defparam desc1817.INIT=64'h000000008880AAA2;
  LUT6 desc1818(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_112));
defparam desc1818.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1819(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_104));
defparam desc1819.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1820(.I0(s_opb_i[6:6]),.I1(s_opb_i[7:7]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_108));
defparam desc1820.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1821(.I0(s_opb_i[13:13]),.I1(s_opb_i[12:12]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_100));
defparam desc1821.INIT=64'hACACACCCAAAAAACA;
  LUT6 desc1822(.I0(s_opb_i[14:14]),.I1(s_opb_i[15:15]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_2194));
defparam desc1822.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1823(.I0(s_opb_i[4:4]),.I1(s_opb_i[5:5]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_110));
defparam desc1823.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1824(.I0(s_opb_i[8:8]),.I1(s_opb_i[9:9]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_106));
defparam desc1824.INIT=64'hCACACAAACCCCCCAC;
  LUT6 desc1825(.I0(s_opb_i[1:1]),.I1(s_opb_i[0:0]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_101));
defparam desc1825.INIT=64'hACACACCCAAAAAACA;
  LUT6 desc1826(.I0(s_opb_i[19:19]),.I1(s_opb_i[18:18]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_20));
defparam desc1826.INIT=64'hACACACCCAAAAAACA;
  LUT6 desc1827(.I0(s_opb_i[17:17]),.I1(s_opb_i[16:16]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.I5(N_143_mux),.O(N_18));
defparam desc1827.INIT=64'hACACACCCAAAAAACA;
  LUT5 un4_s_expb_in_2_i_o3_RNIODKRI_0(.I0(s_opb_i[22:22]),.I1(s_opb_i[23:23]),.I2(N_1083),.I3(N_143_mux),.I4(un11_s_exp_10_o_5[0:0]),.O(un11_s_exp_10_o_axb_0_i));
defparam un4_s_expb_in_2_i_o3_RNIODKRI_0.INIT=32'h5702A8FD;
  LUT2_L desc1828(.I0(s_opa_i_0[28:28]),.I1(s_opa_i_0[25:25]),.LO(result_i_o2_0_0));
defparam desc1828.INIT=4'hE;
  LUT2 un4_s_expb_in_2_i_o2_1_c(.I0(s_opb_i_0_2),.I1(s_opb_i_0_5),.O(un4_s_expb_in_2_i_o2_1));
defparam un4_s_expb_in_2_i_o2_1_c.INIT=4'hE;
  LUT1_L un11_s_exp_10_o_axb_9_cZ(.I0(un11_s_exp_10_o_5[9:9]),.LO(un11_s_exp_10_o_axb_9));
defparam un11_s_exp_10_o_axb_9_cZ.INIT=2'h2;
  LUT1_L un11_s_exp_10_o_axb_8_cZ(.I0(un11_s_exp_10_o_5[8:8]),.LO(un11_s_exp_10_o_axb_8));
defparam un11_s_exp_10_o_axb_8_cZ.INIT=2'h2;
  LUT1_L un11_s_exp_10_o_axb_7_cZ(.I0(un11_s_exp_10_o_5[7:7]),.LO(un11_s_exp_10_o_axb_7));
defparam un11_s_exp_10_o_axb_7_cZ.INIT=2'h2;
  LUT1_L un11_s_exp_10_o_axb_6_cZ(.I0(un11_s_exp_10_o_5[6:6]),.LO(un11_s_exp_10_o_axb_6));
defparam un11_s_exp_10_o_axb_6_cZ.INIT=2'h2;
  LUT1_L un11_s_exp_10_o_axb_5_cZ(.I0(un11_s_exp_10_o_5[5:5]),.LO(un11_s_exp_10_o_axb_5));
defparam un11_s_exp_10_o_axb_5_cZ.INIT=2'h2;
  LUT3 desc1829(.I0(s_opa_i[6:6]),.I1(s_opa_i[7:7]),.I2(s_opa_i[8:8]),.O(N_384));
defparam desc1829.INIT=8'hF2;
  LUT6 desc1830(.I0(s_opa_i[30:30]),.I1(s_opa_i_0[29:29]),.I2(s_opa_i[26:26]),.I3(s_opa_i[27:27]),.I4(s_opa_i[23:23]),.I5(result_i_o2_0_0),.O(N_1077));
defparam desc1830.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc1831(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[1:1]),.I4(s_opb_i[5:5]),.I5(s_opb_i[0:0]),.LO(N_290));
defparam desc1831.INIT=64'hFFFFF1F1FFFFF1F0;
  LUT6 desc1832(.I0(s_opb_i[21:21]),.I1(s_opb_i[17:17]),.I2(s_opb_i[19:19]),.I3(s_opb_i[20:20]),.I4(s_opb_i[22:22]),.I5(N_1084_i),.O(v_count_2_0[4:4]));
defparam desc1832.INIT=64'h0000000100000000;
  LUT6_L desc1833(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[1:1]),.I3(s_opa_i[4:4]),.I4(s_opa_i[0:0]),.I5(s_opa_i[5:5]),.LO(N_1160));
defparam desc1833.INIT=64'hFFFFFFFFFF11FF10;
  LUT6 un4_s_expb_in_2_i_o3(.I0(s_opb_i_0_2),.I1(s_opb_i_0_5),.I2(s_opb_i[24:24]),.I3(s_opb_i[28:28]),.I4(s_opb_i[27:27]),.I5(un4_s_expb_in_2_i_o2_0),.O(N_1083));
defparam un4_s_expb_in_2_i_o3.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT5_L desc1834(.I0(s_opb_i[6:6]),.I1(s_opb_i[8:8]),.I2(s_opb_i[9:9]),.I3(s_opb_i[7:7]),.I4(N_290),.LO(N_296));
defparam desc1834.INIT=32'hFCFDFCFC;
  LUT5 desc1835(.I0(s_opb_i[4:4]),.I1(N_1050),.I2(N_1052),.I3(N_2220),.I4(N_1051),.O(v_count_0_0_a5_0_1_1[2:2]));
defparam desc1835.INIT=32'h0C0C4C0C;
  LUT6 desc1836(.I0(s_opa_i[16:16]),.I1(s_opa_i[14:14]),.I2(s_opa_i[15:15]),.I3(N_240_2),.I4(v_count_1_0_a2_1_4),.I5(N_432),.O(v_count_1_0_2));
defparam desc1836.INIT=64'hFFFFAE0000000000;
  LUT5 desc1837(.I0(s_opa_i[7:7]),.I1(s_opa_i[4:4]),.I2(s_opa_i[10:10]),.I3(s_opa_i[5:5]),.I4(N_1087),.O(N_238));
defparam desc1837.INIT=32'h0F0B0F0A;
  LUT6_L desc1838(.I0(s_opa_i[8:8]),.I1(s_opa_i[10:10]),.I2(s_opa_i[11:11]),.I3(s_opa_i[9:9]),.I4(un2_s_snan_o_8),.I5(N_1160),.LO(N_1216));
defparam desc1838.INIT=64'h0303030203020302;
  LUT6 desc1839(.I0(s_opa_i[18:18]),.I1(s_opa_i[19:19]),.I2(s_opa_i[21:21]),.I3(s_opa_i[20:20]),.I4(s_opa_i[24:24]),.I5(N_1077),.O(v_count_1_0_1));
defparam desc1839.INIT=64'h0000000000000F02;
  LUT6 desc1840(.I0(s_opa_i[21:21]),.I1(s_opa_i[22:22]),.I2(s_opa_i[20:20]),.I3(s_opa_i[24:24]),.I4(un2_s_snan_o_22),.I5(N_1077),.O(N_1227));
defparam desc1840.INIT=64'h0000000000010000;
  LUT6 desc1841(.I0(s_opa_i[12:12]),.I1(v_count_1_0_a2_0),.I2(v_count_1_0_a2_7_i_0),.I3(N_240_2),.I4(N_238),.I5(N_432),.O(N_396));
defparam desc1841.INIT=64'h88008C0000000000;
  LUT6 desc1842(.I0(s_opb_i[21:21]),.I1(s_opb_i[20:20]),.I2(s_opb_i[22:22]),.I3(result_2_16),.I4(v_count_0_0_a5_0_1_1[2:2]),.I5(N_1084_i),.O(v_count_0[2:2]));
defparam desc1842.INIT=64'h0101010000000000;
  LUT2_L un11_s_exp_10_o_axb_2_cZ(.I0(v_count_0[2:2]),.I1(un11_s_exp_10_o_5[2:2]),.LO(un11_s_exp_10_o_axb_2));
defparam un11_s_exp_10_o_axb_2_cZ.INIT=4'h6;
  LUT6 desc1843(.I0(s_opb_i[22:22]),.I1(result_2_11),.I2(N_304_1),.I3(result_2_10),.I4(N_341),.I5(N_1084_i),.O(v_count[1:1]));
defparam desc1843.INIT=64'h4455445400000000;
  LUT6 desc1844(.I0(s_opa_i[2:2]),.I1(s_opa_i[1:1]),.I2(N_399),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(N_1617));
defparam desc1844.INIT=64'hCCCCCCCCCCCCCCCA;
  LUT6 desc1845(.I0(s_opa_i[1:1]),.I1(s_opa_i[0:0]),.I2(N_399),.I3(v_count_1_0_1),.I4(N_396),.I5(v_count_1_0_2),.O(N_2103));
defparam desc1845.INIT=64'hCCCCCCCCCCCCCCCA;
  LUT2_L un11_s_exp_10_o_axb_1_cZ(.I0(v_count[1:1]),.I1(un11_s_exp_10_o_5[1:1]),.LO(un11_s_exp_10_o_axb_1));
defparam un11_s_exp_10_o_axb_1_cZ.INIT=4'h6;
  LUT6 un11_s_exp_10_o_5_axb_1_cZ(.I0(s_opa_i[21:21]),.I1(s_opa_i[22:22]),.I2(s_opa_i[20:20]),.I3(un11_s_exp_10_o_6[1:1]),.I4(v_count_1_0_0_a2_0[1:1]),.I5(result_i_o3_lut6_2_O6),.O(un11_s_exp_10_o_5_axb_1));
defparam un11_s_exp_10_o_5_axb_1_cZ.INIT=64'h00FF00FF33CC32CD;
  LUT6 desc1846(.I0(s_opb_i[2:2]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[1:1]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_121));
defparam desc1846.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1847(.I0(s_opb_i[6:6]),.I1(s_opb_i[3:3]),.I2(s_opb_i[4:4]),.I3(s_opb_i[5:5]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_124));
defparam desc1847.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1848(.I0(s_opb_i[6:6]),.I1(s_opb_i[8:8]),.I2(s_opb_i[5:5]),.I3(s_opb_i[7:7]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_126));
defparam desc1848.INIT=64'hF0F0FF00AAAACCCC;
  LUT6 desc1849(.I0(s_opb_i[10:10]),.I1(s_opb_i[8:8]),.I2(s_opb_i[9:9]),.I3(s_opb_i[7:7]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_128));
defparam desc1849.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc1850(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[12:12]),.I3(s_opb_i[9:9]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_130));
defparam desc1850.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1851(.I0(s_opb_i[11:11]),.I1(s_opb_i[13:13]),.I2(s_opb_i[14:14]),.I3(s_opb_i[12:12]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_132));
defparam desc1851.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1852(.I0(s_opb_i[13:13]),.I1(s_opb_i[14:14]),.I2(s_opb_i[15:15]),.I3(s_opb_i[16:16]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_41));
defparam desc1852.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1853(.I0(s_opb_i[15:15]),.I1(s_opb_i[17:17]),.I2(s_opb_i[16:16]),.I3(s_opb_i[18:18]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_43));
defparam desc1853.INIT=64'hAAAACCCCF0F0FF00;
  LUT6 desc1854(.I0(s_opb_i[17:17]),.I1(s_opb_i[19:19]),.I2(s_opb_i[20:20]),.I3(s_opb_i[18:18]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_45));
defparam desc1854.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1855(.I0(s_opb_i[21:21]),.I1(s_opb_i[19:19]),.I2(s_opb_i[20:20]),.I3(s_opb_i[22:22]),.I4(v_count[1:1]),.I5(v_count[0:0]),.O(N_47));
defparam desc1855.INIT=64'hCCCCAAAAF0F0FF00;
  LUT6 desc1856(.I0(s_opa_i[16:16]),.I1(s_opa_i[14:14]),.I2(s_opa_i[13:13]),.I3(s_opa_i[15:15]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_41_0));
defparam desc1856.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc1857(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opa_i[15:15]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_43_0));
defparam desc1857.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1858(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opa_i[19:19]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_44));
defparam desc1858.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1859(.I0(s_opa_i[17:17]),.I1(s_opa_i[18:18]),.I2(s_opa_i[19:19]),.I3(s_opa_i[20:20]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_45_0));
defparam desc1859.INIT=64'hAAAAF0F0CCCCFF00;
  LUT6 desc1860(.I0(s_opa_i[19:19]),.I1(s_opa_i[21:21]),.I2(s_opa_i[22:22]),.I3(s_opa_i[20:20]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_47_0));
defparam desc1860.INIT=64'hAAAACCCCFF00F0F0;
  LUT6 desc1861(.I0(s_opa_i[12:12]),.I1(s_opa_i[10:10]),.I2(s_opa_i[11:11]),.I3(s_opa_i[9:9]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1628));
defparam desc1861.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc1862(.I0(s_opa_i[14:14]),.I1(s_opa_i[12:12]),.I2(s_opa_i[13:13]),.I3(s_opa_i[11:11]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1630));
defparam desc1862.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc1863(.I0(s_opa_i[7:7]),.I1(s_opa_i[8:8]),.I2(s_opa_i[10:10]),.I3(s_opa_i[9:9]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1626));
defparam desc1863.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1864(.I0(s_opa_i[6:6]),.I1(s_opa_i[7:7]),.I2(s_opa_i[8:8]),.I3(s_opa_i[5:5]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1624));
defparam desc1864.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc1865(.I0(s_opa_i[6:6]),.I1(s_opa_i[3:3]),.I2(s_opa_i[4:4]),.I3(s_opa_i[5:5]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1622));
defparam desc1865.INIT=64'hCCCCFF00F0F0AAAA;
  LUT6 desc1866(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[1:1]),.I3(s_opa_i[4:4]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1619));
defparam desc1866.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc1867(.I0(s_opa_i[18:18]),.I1(s_opa_i[19:19]),.I2(s_opa_i[21:21]),.I3(s_opa_i[20:20]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_46));
defparam desc1867.INIT=64'hAAAAFF00CCCCF0F0;
  LUT6 desc1868(.I0(s_opa_i[2:2]),.I1(s_opa_i[3:3]),.I2(s_opa_i[1:1]),.I3(s_opa_i[0:0]),.I4(v_count_0_1),.I5(v_count_0_0),.O(N_1620));
defparam desc1868.INIT=64'hFF00AAAAF0F0CCCC;
  LUT5 desc1869(.I0(s_opb_i[2:2]),.I1(s_opb_i[1:1]),.I2(s_opb_i[0:0]),.I3(v_count[1:1]),.I4(v_count[0:0]),.O(N_27));
defparam desc1869.INIT=32'h00CCF0AA;
  LUT5 desc1870(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_110),.I3(N_112),.I4(N_101),.O(N_54));
defparam desc1870.INIT=32'h76325410;
  LUT6 desc1871(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_108),.I3(N_110),.I4(N_112),.I5(N_101),.O(N_56));
defparam desc1871.INIT=64'hFEBADC9876325410;
  LUT6 desc1872(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_106),.I3(N_108),.I4(N_110),.I5(N_112),.O(N_58));
defparam desc1872.INIT=64'hFEBADC9876325410;
  LUT6 desc1873(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_104),.I3(N_106),.I4(N_108),.I5(N_110),.O(N_60));
defparam desc1873.INIT=64'hFEBADC9876325410;
  LUT6 desc1874(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_100),.I3(N_104),.I4(N_106),.I5(N_108),.O(N_62));
defparam desc1874.INIT=64'hFEBADC9876325410;
  LUT6 desc1875(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_100),.I3(N_104),.I4(N_106),.I5(N_2194),.O(N_64));
defparam desc1875.INIT=64'hFBD97351EAC86240;
  LUT6 desc1876(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_18),.I3(N_100),.I4(N_104),.I5(N_2194),.O(N_66));
defparam desc1876.INIT=64'hFEDC7654BA983210;
  LUT6 desc1877(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(N_20),.I3(N_18),.I4(N_100),.I5(N_2194),.O(N_68));
defparam desc1877.INIT=64'hFEBA7632DC985410;
  LUT6 desc1878(.I0(N_22),.I1(v_count_0[2:2]),.I2(v_count[1:1]),.I3(N_20),.I4(N_18),.I5(N_2194),.O(N_70));
defparam desc1878.INIT=64'hFECEF2C23E0E3202;
  LUT6 desc1879(.I0(s_opb_i[1:1]),.I1(s_opb_i[0:0]),.I2(v_count_0[2:2]),.I3(v_count[1:1]),.I4(v_count_0[3:3]),.I5(v_count[0:0]),.O(N_74));
defparam desc1879.INIT=64'h0000000C0000000A;
  LUT6 desc1880(.I0(s_opa_i[0:0]),.I1(v_count_0_1),.I2(v_count_2),.I3(N_1617),.I4(v_count_i),.I5(N_1622),.O(N_55));
defparam desc1880.INIT=64'hBF8F3F0FB0803000;
  LUT5_L desc1881(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_25),.I3(N_126),.I4(N_121),.LO(pre_norm_div_dvsor[8:8]));
defparam desc1881.INIT=32'h73625140;
  LUT5_L desc1882(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(v_count_0[3:3]),.I3(N_101),.I4(N_58),.LO(pre_norm_div_dvsor[9:9]));
defparam desc1882.INIT=32'h1F0F1000;
  LUT6_L desc1883(.I0(v_count_0[2:2]),.I1(v_count[1:1]),.I2(v_count_0[3:3]),.I3(N_112),.I4(N_101),.I5(N_60),.LO(pre_norm_div_dvsor[11:11]));
defparam desc1883.INIT=64'h5F4F1F0F50401000;
  LUT6_L desc1884(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_41),.I3(N_130),.I4(N_126),.I5(N_121),.LO(N_89));
defparam desc1884.INIT=64'hFEDCBA9876543210;
  LUT6_L desc1885(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_43),.I3(N_132),.I4(N_128),.I5(N_124),.LO(N_91));
defparam desc1885.INIT=64'hFEDCBA9876543210;
  LUT6_L desc1886(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_45),.I3(N_41),.I4(N_130),.I5(N_126),.LO(N_93));
defparam desc1886.INIT=64'hFEDCBA9876543210;
  LUT6_L desc1887(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_47),.I3(N_43),.I4(N_132),.I5(N_128),.LO(N_95));
defparam desc1887.INIT=64'hFEDCBA9876543210;
  LUT6_L desc1888(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_25),.I3(N_130),.I4(N_126),.I5(N_121),.LO(pre_norm_div_dvsor[12:12]));
defparam desc1888.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc1889(.I0(v_count_3),.I1(v_count_2),.I2(N_47_0),.I3(N_43_0),.I4(N_1630),.I5(N_1626),.O(N_95_0));
defparam desc1889.INIT=64'hFEBADC9876325410;
  LUT5_L desc1890(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_128),.I3(N_124),.I4(N_27),.LO(pre_norm_div_dvsor[10:10]));
defparam desc1890.INIT=32'h76543210;
  LUT6_L desc1891(.I0(v_count_0[2:2]),.I1(v_count_0[3:3]),.I2(N_132),.I3(N_128),.I4(N_124),.I5(N_27),.LO(pre_norm_div_dvsor[14:14]));
defparam desc1891.INIT=64'hFEDCBA9876543210;
  LUT5_L desc1892(.I0(v_count[4:4]),.I1(v_count_0[3:3]),.I2(N_74),.I3(N_66),.I4(N_58),.LO(pre_norm_div_dvsor[17:17]));
defparam desc1892.INIT=32'hF5E4B1A0;
  LUT5_L desc1893(.I0(v_count[4:4]),.I1(v_count_0[3:3]),.I2(N_68),.I3(N_76),.I4(N_60),.LO(pre_norm_div_dvsor[19:19]));
defparam desc1893.INIT=32'hFE54BA10;
  LUT5_L desc1894(.I0(v_count[4:4]),.I1(v_count_0[3:3]),.I2(N_70),.I3(N_62),.I4(N_54),.LO(pre_norm_div_dvsor[21:21]));
defparam desc1894.INIT=32'h76325410;
  LUT5 desc1895(.I0(v_count_3),.I1(v_count_0_4),.I2(N_70_0),.I3(N_27_0),.I4(N_1238),.O(pre_norm_div_dvdnd_11));
defparam desc1895.INIT=32'h54761032;
  XORCY un11_s_exp_10_o_s_9(.LI(un11_s_exp_10_o_axb_9),.CI(un11_s_exp_10_o_cry_8),.O(un11_s_exp_10_o_0[9:9]));
  XORCY un11_s_exp_10_o_s_8(.LI(un11_s_exp_10_o_axb_8),.CI(un11_s_exp_10_o_cry_7),.O(un11_s_exp_10_o_0[8:8]));
  MUXCY_L un11_s_exp_10_o_cry_8_cZ(.DI(GND),.CI(un11_s_exp_10_o_cry_7),.S(un11_s_exp_10_o_axb_8),.LO(un11_s_exp_10_o_cry_8));
  XORCY un11_s_exp_10_o_s_7(.LI(un11_s_exp_10_o_axb_7),.CI(un11_s_exp_10_o_cry_6),.O(un11_s_exp_10_o_0[7:7]));
  MUXCY_L un11_s_exp_10_o_cry_7_cZ(.DI(GND),.CI(un11_s_exp_10_o_cry_6),.S(un11_s_exp_10_o_axb_7),.LO(un11_s_exp_10_o_cry_7));
  XORCY un11_s_exp_10_o_s_6(.LI(un11_s_exp_10_o_axb_6),.CI(un11_s_exp_10_o_cry_5),.O(un11_s_exp_10_o_0[6:6]));
  MUXCY_L un11_s_exp_10_o_cry_6_cZ(.DI(GND),.CI(un11_s_exp_10_o_cry_5),.S(un11_s_exp_10_o_axb_6),.LO(un11_s_exp_10_o_cry_6));
  XORCY un11_s_exp_10_o_s_5(.LI(un11_s_exp_10_o_axb_5),.CI(un11_s_exp_10_o_cry_4),.O(un11_s_exp_10_o_0[5:5]));
  MUXCY_L un11_s_exp_10_o_cry_5_cZ(.DI(GND),.CI(un11_s_exp_10_o_cry_4),.S(un11_s_exp_10_o_axb_5),.LO(un11_s_exp_10_o_cry_5));
  XORCY un11_s_exp_10_o_s_4(.LI(un11_s_exp_10_o_axb_4),.CI(un11_s_exp_10_o_cry_3),.O(un11_s_exp_10_o_0[4:4]));
  MUXCY_L un11_s_exp_10_o_cry_4_cZ(.DI(un11_s_exp_10_o_5[4:4]),.CI(un11_s_exp_10_o_cry_3),.S(un11_s_exp_10_o_axb_4),.LO(un11_s_exp_10_o_cry_4));
  XORCY un11_s_exp_10_o_s_3(.LI(un11_s_exp_10_o_axb_3),.CI(un11_s_exp_10_o_cry_2),.O(un11_s_exp_10_o_0[3:3]));
  MUXCY_L un11_s_exp_10_o_cry_3_cZ(.DI(un11_s_exp_10_o_5[3:3]),.CI(un11_s_exp_10_o_cry_2),.S(un11_s_exp_10_o_axb_3),.LO(un11_s_exp_10_o_cry_3));
  XORCY un11_s_exp_10_o_s_2(.LI(un11_s_exp_10_o_axb_2),.CI(un11_s_exp_10_o_cry_1),.O(un11_s_exp_10_o_0[2:2]));
  MUXCY_L un11_s_exp_10_o_cry_2_cZ(.DI(un11_s_exp_10_o_5[2:2]),.CI(un11_s_exp_10_o_cry_1),.S(un11_s_exp_10_o_axb_2),.LO(un11_s_exp_10_o_cry_2));
  XORCY un11_s_exp_10_o_s_1(.LI(un11_s_exp_10_o_axb_1),.CI(un11_s_exp_10_o_cry_0),.O(un11_s_exp_10_o_0[1:1]));
  MUXCY_L un11_s_exp_10_o_cry_1_cZ(.DI(un11_s_exp_10_o_5[1:1]),.CI(un11_s_exp_10_o_cry_0),.S(un11_s_exp_10_o_axb_1),.LO(un11_s_exp_10_o_cry_1));
  MUXCY_L un11_s_exp_10_o_cry_0_cZ(.DI(v_count[0:0]),.CI(VCC),.S(un11_s_exp_10_o_axb_0),.LO(un11_s_exp_10_o_cry_0));
  XORCY un11_s_exp_10_o_5_s_9(.LI(un11_s_exp_10_o_5_s_9_true),.CI(un11_s_exp_10_o_5_cry_8),.O(un11_s_exp_10_o_5[9:9]));
  XORCY un11_s_exp_10_o_5_s_8(.LI(un11_s_exp_10_o_6_i[8:8]),.CI(un11_s_exp_10_o_5_cry_7),.O(un11_s_exp_10_o_5[8:8]));
  MUXCY_L un11_s_exp_10_o_5_cry_8_cZ(.DI(VCC),.CI(un11_s_exp_10_o_5_cry_7),.S(un11_s_exp_10_o_6_i[8:8]),.LO(un11_s_exp_10_o_5_cry_8));
  XORCY un11_s_exp_10_o_5_s_7(.LI(un11_s_exp_10_o_5_axb_7),.CI(un11_s_exp_10_o_5_cry_6),.O(un11_s_exp_10_o_5[7:7]));
  MUXCY_L un11_s_exp_10_o_5_cry_7_cZ(.DI(GND),.CI(un11_s_exp_10_o_5_cry_6),.S(un11_s_exp_10_o_5_axb_7),.LO(un11_s_exp_10_o_5_cry_7));
  XORCY un11_s_exp_10_o_5_s_6(.LI(un11_s_exp_10_o_6_i[6:6]),.CI(un11_s_exp_10_o_5_cry_5),.O(un11_s_exp_10_o_5[6:6]));
  MUXCY_L un11_s_exp_10_o_5_cry_6_cZ(.DI(VCC),.CI(un11_s_exp_10_o_5_cry_5),.S(un11_s_exp_10_o_6_i[6:6]),.LO(un11_s_exp_10_o_5_cry_6));
  XORCY un11_s_exp_10_o_5_s_5(.LI(un11_s_exp_10_o_6_i[5:5]),.CI(un11_s_exp_10_o_5_cry_4),.O(un11_s_exp_10_o_5[5:5]));
  MUXCY_L un11_s_exp_10_o_5_cry_5_cZ(.DI(VCC),.CI(un11_s_exp_10_o_5_cry_4),.S(un11_s_exp_10_o_6_i[5:5]),.LO(un11_s_exp_10_o_5_cry_5));
  XORCY un11_s_exp_10_o_5_s_4(.LI(un11_s_exp_10_o_5_axb_4),.CI(un11_s_exp_10_o_5_cry_3),.O(un11_s_exp_10_o_5[4:4]));
  MUXCY_L un11_s_exp_10_o_5_cry_4_cZ(.DI(un11_s_exp_10_o_6[4:4]),.CI(un11_s_exp_10_o_5_cry_3),.S(un11_s_exp_10_o_5_axb_4),.LO(un11_s_exp_10_o_5_cry_4));
  XORCY un11_s_exp_10_o_5_s_3(.LI(un11_s_exp_10_o_5_axb_3),.CI(un11_s_exp_10_o_5_cry_2),.O(un11_s_exp_10_o_5[3:3]));
  MUXCY_L un11_s_exp_10_o_5_cry_3_cZ(.DI(un11_s_exp_10_o_6[3:3]),.CI(un11_s_exp_10_o_5_cry_2),.S(un11_s_exp_10_o_5_axb_3),.LO(un11_s_exp_10_o_5_cry_3));
  XORCY un11_s_exp_10_o_5_s_2(.LI(un11_s_exp_10_o_5_axb_2),.CI(un11_s_exp_10_o_5_cry_1),.O(un11_s_exp_10_o_5[2:2]));
  MUXCY_L un11_s_exp_10_o_5_cry_2_cZ(.DI(un11_s_exp_10_o_6[2:2]),.CI(un11_s_exp_10_o_5_cry_1),.S(un11_s_exp_10_o_5_axb_2),.LO(un11_s_exp_10_o_5_cry_2));
  XORCY un11_s_exp_10_o_5_s_1(.LI(un11_s_exp_10_o_5_axb_1),.CI(un11_s_exp_10_o_5_cry_0),.O(un11_s_exp_10_o_5[1:1]));
  MUXCY_L un11_s_exp_10_o_5_cry_1_cZ(.DI(un11_s_exp_10_o_6[1:1]),.CI(un11_s_exp_10_o_5_cry_0),.S(un11_s_exp_10_o_5_axb_1),.LO(un11_s_exp_10_o_5_cry_1));
  MUXCY_L un11_s_exp_10_o_5_cry_0_cZ(.DI(v_count_i),.CI(GND),.S(un11_s_exp_10_o_5[0:0]),.LO(un11_s_exp_10_o_5_cry_0));
  XORCY un11_s_exp_10_o_6_s_7(.LI(un11_s_exp_10_o_6_axb_7),.CI(un11_s_exp_10_o_6_cry_6),.O(un11_s_exp_10_o_6[7:7]));
  MUXCY un11_s_exp_10_o_6_cry_7(.DI(s_opa_i_0[30:30]),.CI(un11_s_exp_10_o_6_cry_6),.S(un11_s_exp_10_o_6_axb_7),.O(un11_s_exp_10_o_6_0[8:8]));
  XORCY un11_s_exp_10_o_6_s_6(.LI(un11_s_exp_10_o_6_axb_6),.CI(un11_s_exp_10_o_6_cry_5),.O(un11_s_exp_10_o_6[6:6]));
  MUXCY_L un11_s_exp_10_o_6_cry_6_cZ(.DI(s_opa_i[29:29]),.CI(un11_s_exp_10_o_6_cry_5),.S(un11_s_exp_10_o_6_axb_6),.LO(un11_s_exp_10_o_6_cry_6));
  XORCY un11_s_exp_10_o_6_s_5(.LI(un11_s_exp_10_o_6_axb_5),.CI(un11_s_exp_10_o_6_cry_4),.O(un11_s_exp_10_o_6[5:5]));
  MUXCY_L un11_s_exp_10_o_6_cry_5_cZ(.DI(s_opa_i[28:28]),.CI(un11_s_exp_10_o_6_cry_4),.S(un11_s_exp_10_o_6_axb_5),.LO(un11_s_exp_10_o_6_cry_5));
  XORCY un11_s_exp_10_o_6_s_4(.LI(un11_s_exp_10_o_6_axb_4),.CI(un11_s_exp_10_o_6_cry_3),.O(un11_s_exp_10_o_6[4:4]));
  MUXCY_L un11_s_exp_10_o_6_cry_4_cZ(.DI(s_opa_i_0[27:27]),.CI(un11_s_exp_10_o_6_cry_3),.S(un11_s_exp_10_o_6_axb_4),.LO(un11_s_exp_10_o_6_cry_4));
  XORCY un11_s_exp_10_o_6_s_3(.LI(un11_s_exp_10_o_6_axb_3),.CI(un11_s_exp_10_o_6_cry_2),.O(un11_s_exp_10_o_6[3:3]));
  MUXCY_L un11_s_exp_10_o_6_cry_3_cZ(.DI(s_opa_i_0[26:26]),.CI(un11_s_exp_10_o_6_cry_2),.S(un11_s_exp_10_o_6_axb_3),.LO(un11_s_exp_10_o_6_cry_3));
  XORCY un11_s_exp_10_o_6_s_2(.LI(un11_s_exp_10_o_6_axb_2),.CI(un11_s_exp_10_o_6_cry_1),.O(un11_s_exp_10_o_6[2:2]));
  MUXCY_L un11_s_exp_10_o_6_cry_2_cZ(.DI(s_opa_i[25:25]),.CI(un11_s_exp_10_o_6_cry_1),.S(un11_s_exp_10_o_6_axb_2),.LO(un11_s_exp_10_o_6_cry_2));
  XORCY un11_s_exp_10_o_6_s_1(.LI(un11_s_exp_10_o_6_axb_1),.CI(un11_s_exp_10_o_6_cry_0),.O(un11_s_exp_10_o_6[1:1]));
  MUXCY_L un11_s_exp_10_o_6_cry_1_cZ(.DI(s_opa_i_0[24:24]),.CI(un11_s_exp_10_o_6_cry_0),.S(un11_s_exp_10_o_6_axb_1),.LO(un11_s_exp_10_o_6_cry_1));
  MUXCY_L un11_s_exp_10_o_6_cry_0_cZ(.DI(s_expa_in),.CI(GND),.S(un11_s_exp_10_o_6[0:0]),.LO(un11_s_exp_10_o_6_cry_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT4 desc1896(.I0(v_count_0[2:2]),.I1(v_count[4:4]),.I2(N_27),.I3(N_91),.O(pre_norm_div_dvsor[18:18]));
defparam desc1896.INIT=16'h3340;
  LUT4 desc1897(.I0(v_count_0[3:3]),.I1(v_count_0[2:2]),.I2(v_count[4:4]),.I3(N_27),.O(s_dvdnd_50_o_104_0_e));
defparam desc1897.INIT=16'h0100;
  LUT4 desc1898(.I0(s_opb_i[16:16]),.I1(s_opb_i[18:18]),.I2(v_count_2_0[4:4]),.I3(N_56),.O(pre_norm_div_dvsor[7:7]));
defparam desc1898.INIT=16'hEF00;
  LUT5 desc1899(.I0(N_1055),.I1(s_opb_i[16:16]),.I2(s_opb_i[18:18]),.I3(v_count_2_0[4:4]),.I4(N_56),.O(pre_norm_div_dvsor_0[23:23]));
defparam desc1899.INIT=32'hFFFFFDFF;
  LUT5 desc1900(.I0(s_opa_i[14:14]),.I1(s_opa_i[13:13]),.I2(s_opa_i[12:12]),.I3(s_opa_i[15:15]),.I4(N_1216),.O(N_1219));
defparam desc1900.INIT=32'h00550054;
  LUT2 desc1901(.I0(s_opa_i[13:13]),.I1(s_opa_i[15:15]),.O(v_count_1_0_a2_0));
defparam desc1901.INIT=4'h1;
  LUT2 desc1902(.I0(s_opb_i[21:21]),.I1(s_opb_i[20:20]),.O(result_2_11));
defparam desc1902.INIT=4'hE;
  LUT5 desc1903(.I0(s_opb_i[21:21]),.I1(s_opb_i[20:20]),.I2(s_opb_i[22:22]),.I3(s_opb_i[23:23]),.I4(N_1083),.O(N_22));
defparam desc1903.INIT=32'hAAAAAACE;
  LUT2 desc1904(.I0(s_opb_i[17:17]),.I1(s_opb_i[16:16]),.O(N_304_1));
defparam desc1904.INIT=4'hE;
  LUT4 desc1905(.I0(s_opb_i[17:17]),.I1(s_opb_i[19:19]),.I2(s_opb_i[16:16]),.I3(s_opb_i[18:18]),.O(result_2_16));
defparam desc1905.INIT=16'hFFFE;
  LUT2 desc1906(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.O(N_1041));
defparam desc1906.INIT=4'h1;
  LUT4 desc1907(.I0(s_opb_i[10:10]),.I1(s_opb_i[11:11]),.I2(s_opb_i[8:8]),.I3(s_opb_i[9:9]),.O(N_1052));
defparam desc1907.INIT=16'h0001;
  LUT2 un4_s_expb_in_2_i_o2_2_lut6_2_o6(.I0(s_opb_i[28:28]),.I1(s_opb_i[27:27]),.O(un4_s_expb_in_2_i_o2_2));
defparam un4_s_expb_in_2_i_o2_2_lut6_2_o6.INIT=4'hE;
  LUT3 un4_s_expb_in_2_i_o2_2_lut6_2_o5(.I0(s_opa_i[27:27]),.I1(s_opb_i[27:27]),.I2(s_expa_lt_expb),.O(un4_s_expb_in_2_i_o2_2_lut6_2_O5));
defparam un4_s_expb_in_2_i_o2_2_lut6_2_o5.INIT=8'hAC;
  LUT2 desc1908(.I0(s_opa_i[19:19]),.I1(s_opa_i[21:21]),.O(N_240_2));
defparam desc1908.INIT=4'h1;
  LUT3 desc1909(.I0(s_opa_i[21:21]),.I1(s_opa_i[22:22]),.I2(s_opa_i[20:20]),.O(N_1170));
defparam desc1909.INIT=8'hF4;
  LUT3 desc1910(.I0(s_opb_i[6:6]),.I1(s_opb_i[5:5]),.I2(s_opb_i[7:7]),.O(N_2220));
defparam desc1910.INIT=8'h01;
  LUT5 desc1911(.I0(s_opb_i[6:6]),.I1(s_opb_i[4:4]),.I2(s_opb_i[5:5]),.I3(s_opb_i[7:7]),.I4(N_1051),.O(N_340));
defparam desc1911.INIT=32'h00010000;
  LUT2 desc1912(.I0(s_opa_i[24:24]),.I1(N_1077),.O(result_i_o3_lut6_2_O6));
defparam desc1912.INIT=4'hE;
  LUT4 desc1913(.I0(s_opa_i[24:24]),.I1(s_opb_i[23:23]),.I2(N_1077),.I3(s_expa_lt_expb),.O(N_1140));
defparam desc1913.INIT=16'h0004;
  LUT3 desc1914(.I0(s_opa_i[22:22]),.I1(s_opa_i[24:24]),.I2(N_1077),.O(N_399));
defparam desc1914.INIT=8'h02;
  LUT3 desc1915(.I0(s_opa_i[30:30]),.I1(s_opa_i[26:26]),.I2(s_opa_i[24:24]),.O(un4_s_infa_1));
defparam desc1915.INIT=8'h80;
  LUT3 desc1916(.I0(s_opa_i[17:17]),.I1(s_opa_i[24:24]),.I2(N_1077),.O(N_432));
defparam desc1916.INIT=8'h01;
  LUT4 desc1917(.I0(s_opa_i[24:24]),.I1(N_1077),.I2(s_exp_10_o_0[0:0]),.I3(s_exp_10_o_0[1:1]),.O(s_exp_10_o[1:1]));
defparam desc1917.INIT=16'hEF10;
  LUT5 desc1918(.I0(s_opb_i[16:16]),.I1(s_opb_i[18:18]),.I2(N_340),.I3(N_1055),.I4(v_count_2_0[4:4]),.O(v_count_0[3:3]));
defparam desc1918.INIT=32'h10110000;
  LUT4 desc1919(.I0(s_opb_i[16:16]),.I1(s_opb_i[18:18]),.I2(N_1055),.I3(v_count_2_0[4:4]),.O(v_count[4:4]));
defparam desc1919.INIT=16'h1000;
  LUT5 desc1920(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opa_i[19:19]),.I4(N_1219),.O(v_count_1_0_0_a2_0[1:1]));
defparam desc1920.INIT=32'h000F000E;
  LUT4 desc1921(.I0(s_opa_i[16:16]),.I1(s_opa_i[17:17]),.I2(s_opa_i[18:18]),.I3(s_opa_i[19:19]),.O(un2_s_snan_o_22));
defparam desc1921.INIT=16'h0001;
  LUT2 desc1922(.I0(s_opb_i[13:13]),.I1(s_opb_i[12:12]),.O(N_1049));
defparam desc1922.INIT=4'h1;
  LUT4 desc1923(.I0(s_opb_i[12:12]),.I1(N_987),.I2(s_expa_lt_expb),.I3(N_2240),.O(N_1232_i));
defparam desc1923.INIT=16'h3A0A;
  LUT3 desc1924(.I0(v_count_2),.I1(N_1630),.I2(N_1626),.O(N_63));
defparam desc1924.INIT=8'hE4;
  LUT5 desc1925(.I0(v_count_3),.I1(v_count_2),.I2(N_1630),.I3(N_1626),.I4(N_55),.O(N_1278_i));
defparam desc1925.INIT=32'hFEBA5410;
  LUT3 desc1926(.I0(v_count_0[3:3]),.I1(N_64),.I2(N_56),.O(pre_norm_div_dvsor[15:15]));
defparam desc1926.INIT=8'hE4;
  LUT3 desc1927(.I0(v_count_0[3:3]),.I1(N_62),.I2(N_54),.O(pre_norm_div_dvsor[13:13]));
defparam desc1927.INIT=8'hE4;
  LUT3 desc1928(.I0(v_count_2),.I1(N_1622),.I2(N_1626),.O(N_59));
defparam desc1928.INIT=8'hD8;
  LUT5 desc1929(.I0(v_count_3),.I1(v_count_2),.I2(N_48_0),.I3(N_1622),.I4(N_1626),.O(pre_norm_div_dvdnd_0));
defparam desc1929.INIT=32'hF5B1E4A0;
  LUT5 un4_s_expb_in_2_i_o3_RNIODKRI_o6(.I0(s_opb_i[22:22]),.I1(s_opb_i[23:23]),.I2(N_1083),.I3(N_143_mux),.I4(un11_s_exp_10_o_5[0:0]),.O(un11_s_exp_10_o_axb_0));
defparam un4_s_expb_in_2_i_o3_RNIODKRI_o6.INIT=32'hA8FD5702;
  LUT4 un4_s_expb_in_2_i_o3_RNIODKRI_o5(.I0(s_opb_i[22:22]),.I1(s_opb_i[23:23]),.I2(N_1083),.I3(N_143_mux),.O(v_count[0:0]));
defparam un4_s_expb_in_2_i_o3_RNIODKRI_o5.INIT=16'h5702;
endmodule
module serial_div_inj (fpu_op_i,s_state,pre_norm_div_dvdnd_0,pre_norm_div_dvdnd_8,pre_norm_div_dvdnd_9,pre_norm_div_dvdnd_10,pre_norm_div_dvdnd_11,pre_norm_div_dvdnd_12,pre_norm_div_dvdnd_13,pre_norm_div_dvdnd_14,pre_norm_div_dvdnd_0_d0,pre_norm_div_dvdnd_1,pre_norm_div_dvdnd_2,pre_norm_div_dvdnd_3,pre_norm_div_dvdnd_5,pre_norm_div_dvsor_0,pre_norm_div_dvsor_5,pre_norm_div_dvsor_6,pre_norm_div_dvsor_7,pre_norm_div_dvsor_8,pre_norm_div_dvsor_9,pre_norm_div_dvsor_10,pre_norm_div_dvsor_11,pre_norm_div_dvsor_12,pre_norm_div_dvsor_13,pre_norm_div_dvsor_14,pre_norm_div_dvsor_15,pre_norm_div_dvsor_16,pre_norm_div_dvsor_17,pre_norm_div_dvsor_0_d0,pre_norm_div_dvsor_2,pre_norm_div_dvsor_3,pre_norm_div_dvsor_4,post_norm_sqrt_output,postnorm_addsub_output_o,s_output1_6_2_i_m2,post_norm_div_output,post_norm_mul_output,serial_div_qutnt,serial_div_rmndr,N_2637_i,s_dvdnd_50_o_108_0_e,clk_i,s_dvdnd_50_o_104_0_e,s_dvdnd_50_o_106_0_e,s_dvdnd_50_o_107_0_e,s_dvdnd_50_o_108_0_e_0,s_dvdnd_50_o_106_0_e_0,m49_0_e,s_dvdnd_50_o_105_0_e,s_dvdnd_50_o_102_0_e,m46_0_e,s_dvdnd_50_o_105_0_e_0,s_dvdnd_50_o_109_0_e,s_dvdnd_50_o_102_0_e_0,s_dvdnd_50_o_103_0_e,s_start_i,div_zero_o_0_0,N_1257_i,N_1278_i,N_88,un12_s_state_0_a2_lut6_2_O5,post_norm_div_ine,post_norm_mul_ine,N_564,N_563,N_562,N_561,N_560,N_559,N_558,N_557,N_556,N_555,N_554,N_553,N_552,N_551,N_550,N_549,N_548,N_547,N_546,N_545,N_544,N_543,N_542,N_541,N_538,N_537,N_536,N_503_i,N_502_i,N_501_i,post_norm_sqrt_ine_o,postnorm_addsub_ine_o,s_ine_o_5,div_zero_o_0);
input [2:0] fpu_op_i ;
output s_state ;
input [49:49] pre_norm_div_dvdnd_0 ;
input pre_norm_div_dvdnd_8 ;
input pre_norm_div_dvdnd_9 ;
input pre_norm_div_dvdnd_10 ;
input pre_norm_div_dvdnd_11 ;
input pre_norm_div_dvdnd_12 ;
input pre_norm_div_dvdnd_13 ;
input pre_norm_div_dvdnd_14 ;
input pre_norm_div_dvdnd_0_d0 ;
input pre_norm_div_dvdnd_1 ;
input pre_norm_div_dvdnd_2 ;
input pre_norm_div_dvdnd_3 ;
input pre_norm_div_dvdnd_5 ;
input [23:23] pre_norm_div_dvsor_0 ;
input pre_norm_div_dvsor_5 ;
input pre_norm_div_dvsor_6 ;
input pre_norm_div_dvsor_7 ;
input pre_norm_div_dvsor_8 ;
input pre_norm_div_dvsor_9 ;
input pre_norm_div_dvsor_10 ;
input pre_norm_div_dvsor_11 ;
input pre_norm_div_dvsor_12 ;
input pre_norm_div_dvsor_13 ;
input pre_norm_div_dvsor_14 ;
input pre_norm_div_dvsor_15 ;
input pre_norm_div_dvsor_16 ;
input pre_norm_div_dvsor_17 ;
input pre_norm_div_dvsor_0_d0 ;
input pre_norm_div_dvsor_2 ;
input pre_norm_div_dvsor_3 ;
input pre_norm_div_dvsor_4 ;
input [31:0] post_norm_sqrt_output ;
input [31:0] postnorm_addsub_output_o ;
output [7:6] s_output1_6_2_i_m2 ;
input [31:0] post_norm_div_output ;
input [31:0] post_norm_mul_output ;
output [26:0] serial_div_qutnt ;
output [26:0] serial_div_rmndr ;
output N_2637_i ;
input s_dvdnd_50_o_108_0_e ;
input clk_i ;
input s_dvdnd_50_o_104_0_e ;
input s_dvdnd_50_o_106_0_e ;
input s_dvdnd_50_o_107_0_e ;
input s_dvdnd_50_o_108_0_e_0 ;
input s_dvdnd_50_o_106_0_e_0 ;
input m49_0_e ;
input s_dvdnd_50_o_105_0_e ;
input s_dvdnd_50_o_102_0_e ;
input m46_0_e ;
input s_dvdnd_50_o_105_0_e_0 ;
input s_dvdnd_50_o_109_0_e ;
input s_dvdnd_50_o_102_0_e_0 ;
input s_dvdnd_50_o_103_0_e ;
input s_start_i ;
output div_zero_o_0_0 ;
input N_1257_i ;
input N_1278_i ;
input N_88 ;
input un12_s_state_0_a2_lut6_2_O5 ;
input post_norm_div_ine ;
input post_norm_mul_ine ;
output N_564 ;
output N_563 ;
output N_562 ;
output N_561 ;
output N_560 ;
output N_559 ;
output N_558 ;
output N_557 ;
output N_556 ;
output N_555 ;
output N_554 ;
output N_553 ;
output N_552 ;
output N_551 ;
output N_550 ;
output N_549 ;
output N_548 ;
output N_547 ;
output N_546 ;
output N_545 ;
output N_544 ;
output N_543 ;
output N_542 ;
output N_541 ;
output N_538 ;
output N_537 ;
output N_536 ;
output N_503_i ;
output N_502_i ;
output N_501_i ;
input post_norm_sqrt_ine_o ;
input postnorm_addsub_ine_o ;
output s_ine_o_5 ;
output div_zero_o_0 ;
wire pre_norm_div_dvdnd_8 ;
wire pre_norm_div_dvdnd_9 ;
wire pre_norm_div_dvdnd_10 ;
wire pre_norm_div_dvdnd_11 ;
wire pre_norm_div_dvdnd_12 ;
wire pre_norm_div_dvdnd_13 ;
wire pre_norm_div_dvdnd_14 ;
wire pre_norm_div_dvdnd_0_d0 ;
wire pre_norm_div_dvdnd_1 ;
wire pre_norm_div_dvdnd_2 ;
wire pre_norm_div_dvdnd_3 ;
wire pre_norm_div_dvdnd_5 ;
wire pre_norm_div_dvsor_5 ;
wire pre_norm_div_dvsor_6 ;
wire pre_norm_div_dvsor_7 ;
wire pre_norm_div_dvsor_8 ;
wire pre_norm_div_dvsor_9 ;
wire pre_norm_div_dvsor_10 ;
wire pre_norm_div_dvsor_11 ;
wire pre_norm_div_dvsor_12 ;
wire pre_norm_div_dvsor_13 ;
wire pre_norm_div_dvsor_14 ;
wire pre_norm_div_dvsor_15 ;
wire pre_norm_div_dvsor_16 ;
wire pre_norm_div_dvsor_17 ;
wire pre_norm_div_dvsor_0_d0 ;
wire pre_norm_div_dvsor_2 ;
wire pre_norm_div_dvsor_3 ;
wire pre_norm_div_dvsor_4 ;
wire N_2637_i ;
wire s_dvdnd_50_o_108_0_e ;
wire clk_i ;
wire s_dvdnd_50_o_104_0_e ;
wire s_dvdnd_50_o_106_0_e ;
wire s_dvdnd_50_o_107_0_e ;
wire s_dvdnd_50_o_108_0_e_0 ;
wire s_dvdnd_50_o_106_0_e_0 ;
wire m49_0_e ;
wire s_dvdnd_50_o_105_0_e ;
wire s_dvdnd_50_o_102_0_e ;
wire m46_0_e ;
wire s_dvdnd_50_o_105_0_e_0 ;
wire s_dvdnd_50_o_109_0_e ;
wire s_dvdnd_50_o_102_0_e_0 ;
wire s_dvdnd_50_o_103_0_e ;
wire s_start_i ;
wire div_zero_o_0_0 ;
wire N_1257_i ;
wire N_1278_i ;
wire N_88 ;
wire un12_s_state_0_a2_lut6_2_O5 ;
wire post_norm_div_ine ;
wire post_norm_mul_ine ;
wire N_564 ;
wire N_563 ;
wire N_562 ;
wire N_561 ;
wire N_560 ;
wire N_559 ;
wire N_558 ;
wire N_557 ;
wire N_556 ;
wire N_555 ;
wire N_554 ;
wire N_553 ;
wire N_552 ;
wire N_551 ;
wire N_550 ;
wire N_549 ;
wire N_548 ;
wire N_547 ;
wire N_546 ;
wire N_545 ;
wire N_544 ;
wire N_543 ;
wire N_542 ;
wire N_541 ;
wire N_538 ;
wire N_537 ;
wire N_536 ;
wire N_503_i ;
wire N_502_i ;
wire N_501_i ;
wire post_norm_sqrt_ine_o ;
wire postnorm_addsub_ine_o ;
wire s_ine_o_5 ;
wire div_zero_o_0 ;
wire [23:0] s_dvsor_i ;
wire [4:0] s_count ;
wire [3:3] s_count_RNIQN9Q_O6 ;
wire [49:26] s_dvdnd_i ;
wire [25:0] un17_s_state_cry ;
wire [25:25] un17_s_state_cry_i ;
wire [26:0] s_qutnt_o ;
wire [26:1] s_dvd ;
wire [26:0] v_div_5 ;
wire [19:3] s_qutnt_o_5_iv_i_i ;
wire N_594 ;
wire N_595 ;
wire GND ;
wire VCC ;
wire un17_s_state_df1 ;
wire un17_s_state_lt1 ;
wire N_596 ;
wire N_597 ;
wire un17_s_state_df3 ;
wire un17_s_state_lt3 ;
wire N_598 ;
wire N_599 ;
wire un17_s_state_df5 ;
wire un17_s_state_lt5 ;
wire N_600 ;
wire N_601 ;
wire un17_s_state_df7 ;
wire un17_s_state_lt7 ;
wire N_602 ;
wire N_603 ;
wire un17_s_state_df9 ;
wire un17_s_state_lt9 ;
wire N_604 ;
wire N_605 ;
wire un17_s_state_df11 ;
wire un17_s_state_lt11 ;
wire N_606 ;
wire N_607 ;
wire un17_s_state_df13 ;
wire un17_s_state_lt13 ;
wire N_608 ;
wire N_609 ;
wire un17_s_state_df15 ;
wire un17_s_state_lt15 ;
wire N_610 ;
wire N_611 ;
wire un17_s_state_df17 ;
wire un17_s_state_lt17 ;
wire N_612 ;
wire N_613 ;
wire un17_s_state_df19 ;
wire un17_s_state_lt19 ;
wire N_614 ;
wire N_615 ;
wire un17_s_state_df21 ;
wire un17_s_state_lt21 ;
wire N_2620_i ;
wire N_616 ;
wire un17_s_state_df23 ;
wire un17_s_state_lt23 ;
wire N_2637_i_lut6_2_O5 ;
wire N_445 ;
wire N_453 ;
wire N_452 ;
wire N_466_i_i ;
wire m36_i_m2_lut6_2_O6 ;
wire m36_i_m2_lut6_2_O5 ;
wire m42_i_m2_lut6_2_O6 ;
wire N_497 ;
wire m45_i_m2_lut6_2_O6 ;
wire N_494 ;
wire m48_i_m2_lut6_2_O6 ;
wire N_492 ;
wire m51_i_m2_lut6_2_O6 ;
wire N_485 ;
wire m54_i_m2_lut6_2_O6 ;
wire N_484 ;
wire m57_i_m2_lut6_2_O6 ;
wire m57_i_m2_lut6_2_O5 ;
wire m69_i_m2_lut6_2_O6 ;
wire N_499 ;
wire N_481 ;
wire N_491 ;
wire N_482 ;
wire N_487 ;
wire N_483 ;
wire N_486 ;
wire N_488 ;
wire N_498 ;
wire N_489 ;
wire N_495 ;
wire N_490 ;
wire N_493 ;
wire N_496 ;
wire N_500 ;
wire N_451 ;
wire N_447 ;
wire N_448 ;
wire N_449 ;
wire N_1489_i_0 ;
wire N_1490_i ;
wire N_239_i ;
wire N_1491_i ;
wire N_237_i ;
wire m112_i_0 ;
wire m112_i_1 ;
wire m112_i_2 ;
wire m112_i_3 ;
wire m112_i_4 ;
wire v_div_5_axb_1 ;
wire v_div_5_axb_2 ;
wire v_div_5_axb_3 ;
wire v_div_5_axb_4 ;
wire v_div_5_axb_5 ;
wire v_div_5_axb_6 ;
wire v_div_5_axb_7 ;
wire v_div_5_axb_8 ;
wire v_div_5_axb_9 ;
wire v_div_5_axb_10 ;
wire v_div_5_axb_11 ;
wire v_div_5_axb_12 ;
wire v_div_5_axb_13 ;
wire v_div_5_axb_14 ;
wire v_div_5_axb_15 ;
wire v_div_5_axb_16 ;
wire v_div_5_axb_17 ;
wire v_div_5_axb_18 ;
wire v_div_5_axb_19 ;
wire v_div_5_axb_20 ;
wire v_div_5_axb_21 ;
wire v_div_5_axb_22 ;
wire v_div_5_axb_23 ;
wire N_151_i ;
wire N_2621_i ;
wire un17_s_state_df25 ;
wire v_div_5_axb_0 ;
wire N_2635_i ;
wire N_2629_i ;
wire N_2628_i ;
wire N_2634_i ;
wire N_589_i ;
wire N_2664_0_4 ;
wire N_2664_1_4 ;
wire N_2664_1_0 ;
wire v_div_5_axb_24 ;
wire v_div_5_axb_25 ;
wire v_div_5_axb_26 ;
wire N_2630_i ;
wire N_2627_i ;
wire N_2632_i ;
wire N_2664_2_4 ;
wire N_2664_3_4 ;
wire N_2664_2_0 ;
wire v_div_5_cry_0_cy ;
wire N_504 ;
wire m39_i_m2 ;
wire N_468_i ;
wire N_587_i ;
wire N_584_i ;
wire i30_mux_i ;
wire N_2633_i ;
wire N_2631_i ;
wire v_div_5_cry_0_RNO ;
wire v_div_5_cry_1_RNO ;
wire v_div_5_cry_2_RNO ;
wire v_div_5_cry_3_RNO ;
wire v_div_5_cry_4_RNO ;
wire v_div_5_cry_5_RNO ;
wire v_div_5_cry_6_RNO ;
wire v_div_5_cry_7_RNO ;
wire v_div_5_cry_8_RNO ;
wire v_div_5_cry_9_RNO ;
wire v_div_5_cry_10_RNO ;
wire v_div_5_cry_11_RNO ;
wire v_div_5_cry_12_RNO ;
wire v_div_5_cry_13_RNO ;
wire v_div_5_cry_14_RNO ;
wire v_div_5_cry_15_RNO ;
wire v_div_5_cry_16_RNO ;
wire v_div_5_cry_17_RNO ;
wire v_div_5_cry_18_RNO ;
wire v_div_5_cry_19_RNO ;
wire v_div_5_cry_20_RNO ;
wire v_div_5_cry_21_RNO ;
wire v_div_5_cry_22_RNO ;
wire v_div_5_cry_23_RNO ;
wire v_div_5_cry_25 ;
wire v_div_5_cry_24 ;
wire v_div_5_cry_23 ;
wire v_div_5_cry_22 ;
wire v_div_5_cry_21 ;
wire v_div_5_cry_20 ;
wire v_div_5_cry_19 ;
wire v_div_5_cry_18 ;
wire v_div_5_cry_17 ;
wire v_div_5_cry_16 ;
wire v_div_5_cry_15 ;
wire v_div_5_cry_14 ;
wire v_div_5_cry_13 ;
wire v_div_5_cry_12 ;
wire v_div_5_cry_11 ;
wire v_div_5_cry_10 ;
wire v_div_5_cry_9 ;
wire v_div_5_cry_8 ;
wire v_div_5_cry_7 ;
wire v_div_5_cry_6 ;
wire v_div_5_cry_5 ;
wire v_div_5_cry_4 ;
wire v_div_5_cry_3 ;
wire v_div_5_cry_2 ;
wire v_div_5_cry_1 ;
wire v_div_5_cry_0 ;
wire N_391 ;
wire N_390 ;
wire N_389 ;
wire N_388 ;
wire N_387 ;
wire N_386 ;
wire N_385 ;
wire N_384 ;
wire N_383 ;
wire N_382 ;
wire N_381 ;
wire N_380 ;
wire N_379 ;
wire N_378 ;
wire N_377 ;
wire N_376 ;
wire N_375 ;
wire N_374 ;
wire N_373 ;
wire N_372 ;
wire N_371 ;
wire N_370 ;
wire N_369 ;
wire N_368 ;
wire N_367 ;
wire N_366 ;
wire N_365 ;
wire N_364 ;
wire N_363 ;
wire N_1 ;
// instances
  FD desc1930(.Q(s_dvsor_i[6:6]),.D(s_dvdnd_50_o_108_0_e),.C(clk_i));
  FD desc1931(.Q(s_dvsor_i[2:2]),.D(s_dvdnd_50_o_104_0_e),.C(clk_i));
  FD desc1932(.Q(s_dvdnd_i[30:30]),.D(s_dvdnd_50_o_106_0_e),.C(clk_i));
  FD desc1933(.Q(s_dvdnd_i[31:31]),.D(s_dvdnd_50_o_107_0_e),.C(clk_i));
  FD desc1934(.Q(s_dvdnd_i[32:32]),.D(s_dvdnd_50_o_108_0_e_0),.C(clk_i));
  FD desc1935(.Q(s_dvsor_i[4:4]),.D(s_dvdnd_50_o_106_0_e_0),.C(clk_i));
  FD desc1936(.Q(s_dvdnd_i[28:28]),.D(m49_0_e),.C(clk_i));
  FD desc1937(.Q(s_dvdnd_i[29:29]),.D(s_dvdnd_50_o_105_0_e),.C(clk_i));
  FD desc1938(.Q(s_dvsor_i[0:0]),.D(s_dvdnd_50_o_102_0_e),.C(clk_i));
  FD desc1939(.Q(s_dvdnd_i[27:27]),.D(m46_0_e),.C(clk_i));
  FD desc1940(.Q(s_dvsor_i[3:3]),.D(s_dvdnd_50_o_105_0_e_0),.C(clk_i));
  FD desc1941(.Q(s_dvdnd_i[33:33]),.D(s_dvdnd_50_o_109_0_e),.C(clk_i));
  FD desc1942(.Q(s_dvdnd_i[26:26]),.D(s_dvdnd_50_o_102_0_e_0),.C(clk_i));
  FD desc1943(.Q(s_dvsor_i[1:1]),.D(s_dvdnd_50_o_103_0_e),.C(clk_i));
  FDRE desc1944(.Q(s_count[0:0]),.D(N_1490_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDSE desc1945(.Q(s_count[4:4]),.D(N_239_i),.C(clk_i),.S(s_start_i),.CE(s_state));
  FDSE desc1946(.Q(s_count[1:1]),.D(N_466_i_i),.C(clk_i),.S(s_start_i),.CE(s_state));
  FDRE desc1947(.Q(s_count[2:2]),.D(N_1491_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDSE desc1948(.Q(s_count[3:3]),.D(N_237_i),.C(clk_i),.S(s_start_i),.CE(s_state));
  FDS desc1949(.Q(s_state),.D(N_1489_i_0),.C(clk_i),.S(s_start_i));
  LUT6 desc1950(.I0(m112_i_0),.I1(m112_i_1),.I2(m112_i_2),.I3(m112_i_3),.I4(m112_i_4),.I5(s_dvsor_i[22:22]),.O(div_zero_o_0_0));
defparam desc1950.INIT=64'h0000000000000001;
  LUT3 desc1951(.I0(N_594),.I1(s_dvsor_i[1:1]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_1));
defparam desc1951.INIT=8'hA9;
  LUT3 desc1952(.I0(N_595),.I1(s_dvsor_i[2:2]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_2));
defparam desc1952.INIT=8'hA9;
  LUT3 desc1953(.I0(N_596),.I1(s_dvsor_i[3:3]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_3));
defparam desc1953.INIT=8'hA9;
  LUT3 desc1954(.I0(N_597),.I1(s_dvsor_i[4:4]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_4));
defparam desc1954.INIT=8'hA9;
  LUT3 desc1955(.I0(N_598),.I1(s_dvsor_i[5:5]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_5));
defparam desc1955.INIT=8'hA9;
  LUT3 desc1956(.I0(N_599),.I1(s_dvsor_i[6:6]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_6));
defparam desc1956.INIT=8'hA9;
  LUT3 desc1957(.I0(N_600),.I1(s_dvsor_i[7:7]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_7));
defparam desc1957.INIT=8'hA9;
  LUT3 desc1958(.I0(N_601),.I1(s_dvsor_i[8:8]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_8));
defparam desc1958.INIT=8'hA9;
  LUT3 desc1959(.I0(N_602),.I1(s_dvsor_i[9:9]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_9));
defparam desc1959.INIT=8'hA9;
  LUT3 desc1960(.I0(N_603),.I1(s_dvsor_i[10:10]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_10));
defparam desc1960.INIT=8'hA9;
  LUT3 desc1961(.I0(N_604),.I1(s_dvsor_i[11:11]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_11));
defparam desc1961.INIT=8'hA9;
  LUT3 desc1962(.I0(N_605),.I1(s_dvsor_i[12:12]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_12));
defparam desc1962.INIT=8'hA9;
  LUT3 desc1963(.I0(N_606),.I1(s_dvsor_i[13:13]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_13));
defparam desc1963.INIT=8'hA9;
  LUT3 desc1964(.I0(N_607),.I1(s_dvsor_i[14:14]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_14));
defparam desc1964.INIT=8'hA9;
  LUT3 desc1965(.I0(N_608),.I1(s_dvsor_i[15:15]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_15));
defparam desc1965.INIT=8'hA9;
  LUT3 desc1966(.I0(N_609),.I1(s_dvsor_i[16:16]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_16));
defparam desc1966.INIT=8'hA9;
  LUT3 desc1967(.I0(N_610),.I1(s_dvsor_i[17:17]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_17));
defparam desc1967.INIT=8'hA9;
  LUT3 desc1968(.I0(N_611),.I1(s_dvsor_i[18:18]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_18));
defparam desc1968.INIT=8'hA9;
  LUT3 desc1969(.I0(N_612),.I1(s_dvsor_i[19:19]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_19));
defparam desc1969.INIT=8'hA9;
  LUT3 desc1970(.I0(N_613),.I1(s_dvsor_i[20:20]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_20));
defparam desc1970.INIT=8'hA9;
  LUT3 desc1971(.I0(N_614),.I1(s_dvsor_i[21:21]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_21));
defparam desc1971.INIT=8'hA9;
  LUT3 desc1972(.I0(N_615),.I1(s_dvsor_i[22:22]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_22));
defparam desc1972.INIT=8'hA9;
  LUT3 desc1973(.I0(N_616),.I1(s_dvsor_i[23:23]),.I2(un17_s_state_cry[25:25]),.O(v_div_5_axb_23));
defparam desc1973.INIT=8'hA9;
  LUT1 v_div_5_cry_0_cy_RNO(.I0(un17_s_state_cry[25:25]),.O(un17_s_state_cry_i[25:25]));
defparam v_div_5_cry_0_cy_RNO.INIT=2'h1;
  LUT2 un17_s_state_df25_cZ(.I0(N_151_i),.I1(N_2621_i),.O(un17_s_state_df25));
defparam un17_s_state_df25_cZ.INIT=4'h1;
  FDR desc1974(.Q(serial_div_qutnt[0:0]),.D(s_qutnt_o[0:0]),.C(clk_i),.R(s_start_i));
  FDR desc1975(.Q(serial_div_qutnt[2:2]),.D(s_qutnt_o[2:2]),.C(clk_i),.R(s_start_i));
  FDR desc1976(.Q(serial_div_qutnt[4:4]),.D(s_qutnt_o[4:4]),.C(clk_i),.R(s_start_i));
  FDR desc1977(.Q(serial_div_qutnt[5:5]),.D(s_qutnt_o[5:5]),.C(clk_i),.R(s_start_i));
  FDR desc1978(.Q(serial_div_qutnt[16:16]),.D(s_qutnt_o[16:16]),.C(clk_i),.R(s_start_i));
  FDR desc1979(.Q(serial_div_qutnt[18:18]),.D(s_qutnt_o[18:18]),.C(clk_i),.R(s_start_i));
  FDR desc1980(.Q(serial_div_qutnt[21:21]),.D(s_qutnt_o[21:21]),.C(clk_i),.R(s_start_i));
  FDR desc1981(.Q(serial_div_qutnt[22:22]),.D(s_qutnt_o[22:22]),.C(clk_i),.R(s_start_i));
  FDR desc1982(.Q(serial_div_qutnt[23:23]),.D(s_qutnt_o[23:23]),.C(clk_i),.R(s_start_i));
  FDR desc1983(.Q(serial_div_qutnt[26:26]),.D(s_qutnt_o[26:26]),.C(clk_i),.R(s_start_i));
  FD desc1984(.Q(s_dvdnd_i[42:42]),.D(pre_norm_div_dvdnd_8),.C(clk_i));
  FD desc1985(.Q(s_dvdnd_i[43:43]),.D(pre_norm_div_dvdnd_9),.C(clk_i));
  FD desc1986(.Q(s_dvdnd_i[44:44]),.D(pre_norm_div_dvdnd_10),.C(clk_i));
  FD desc1987(.Q(s_dvdnd_i[45:45]),.D(pre_norm_div_dvdnd_11),.C(clk_i));
  FD desc1988(.Q(s_dvdnd_i[46:46]),.D(pre_norm_div_dvdnd_12),.C(clk_i));
  FD desc1989(.Q(s_dvdnd_i[47:47]),.D(pre_norm_div_dvdnd_13),.C(clk_i));
  FD desc1990(.Q(s_dvdnd_i[48:48]),.D(pre_norm_div_dvdnd_14),.C(clk_i));
  FD desc1991(.Q(s_dvdnd_i[49:49]),.D(pre_norm_div_dvdnd_0[49:49]),.C(clk_i));
  FD desc1992(.Q(s_dvdnd_i[34:34]),.D(pre_norm_div_dvdnd_0_d0),.C(clk_i));
  FD desc1993(.Q(s_dvdnd_i[35:35]),.D(pre_norm_div_dvdnd_1),.C(clk_i));
  FD desc1994(.Q(s_dvdnd_i[36:36]),.D(pre_norm_div_dvdnd_2),.C(clk_i));
  FD desc1995(.Q(s_dvdnd_i[37:37]),.D(pre_norm_div_dvdnd_3),.C(clk_i));
  FD desc1996(.Q(s_dvdnd_i[38:38]),.D(N_1257_i),.C(clk_i));
  FD desc1997(.Q(s_dvdnd_i[39:39]),.D(pre_norm_div_dvdnd_5),.C(clk_i));
  FD desc1998(.Q(s_dvdnd_i[40:40]),.D(N_1278_i),.C(clk_i));
  FD desc1999(.Q(s_dvdnd_i[41:41]),.D(N_88),.C(clk_i));
  FD desc2000(.Q(s_dvsor_i[10:10]),.D(pre_norm_div_dvsor_5),.C(clk_i));
  FD desc2001(.Q(s_dvsor_i[11:11]),.D(pre_norm_div_dvsor_6),.C(clk_i));
  FD desc2002(.Q(s_dvsor_i[12:12]),.D(pre_norm_div_dvsor_7),.C(clk_i));
  FD desc2003(.Q(s_dvsor_i[13:13]),.D(pre_norm_div_dvsor_8),.C(clk_i));
  FD desc2004(.Q(s_dvsor_i[14:14]),.D(pre_norm_div_dvsor_9),.C(clk_i));
  FD desc2005(.Q(s_dvsor_i[15:15]),.D(pre_norm_div_dvsor_10),.C(clk_i));
  FD desc2006(.Q(s_dvsor_i[16:16]),.D(pre_norm_div_dvsor_11),.C(clk_i));
  FD desc2007(.Q(s_dvsor_i[17:17]),.D(pre_norm_div_dvsor_12),.C(clk_i));
  FD desc2008(.Q(s_dvsor_i[18:18]),.D(pre_norm_div_dvsor_13),.C(clk_i));
  FD desc2009(.Q(s_dvsor_i[19:19]),.D(pre_norm_div_dvsor_14),.C(clk_i));
  FD desc2010(.Q(s_dvsor_i[20:20]),.D(pre_norm_div_dvsor_15),.C(clk_i));
  FD desc2011(.Q(s_dvsor_i[21:21]),.D(pre_norm_div_dvsor_16),.C(clk_i));
  FD desc2012(.Q(s_dvsor_i[22:22]),.D(pre_norm_div_dvsor_17),.C(clk_i));
  FD desc2013(.Q(s_dvsor_i[23:23]),.D(pre_norm_div_dvsor_0[23:23]),.C(clk_i));
  FD desc2014(.Q(s_dvsor_i[5:5]),.D(pre_norm_div_dvsor_0_d0),.C(clk_i));
  FD desc2015(.Q(s_dvsor_i[7:7]),.D(pre_norm_div_dvsor_2),.C(clk_i));
  FD desc2016(.Q(s_dvsor_i[8:8]),.D(pre_norm_div_dvsor_3),.C(clk_i));
  FD desc2017(.Q(s_dvsor_i[9:9]),.D(pre_norm_div_dvsor_4),.C(clk_i));
  FDE desc2018(.Q(s_dvd[15:15]),.D(v_div_5[14:14]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2019(.Q(s_dvd[16:16]),.D(v_div_5[15:15]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2020(.Q(s_dvd[17:17]),.D(v_div_5[16:16]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2021(.Q(s_dvd[18:18]),.D(v_div_5[17:17]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2022(.Q(s_dvd[19:19]),.D(v_div_5[18:18]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2023(.Q(s_dvd[20:20]),.D(v_div_5[19:19]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2024(.Q(s_dvd[21:21]),.D(v_div_5[20:20]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2025(.Q(s_dvd[22:22]),.D(v_div_5[21:21]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2026(.Q(s_dvd[23:23]),.D(v_div_5[22:22]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2027(.Q(s_dvd[24:24]),.D(v_div_5[23:23]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2028(.Q(s_dvd[25:25]),.D(v_div_5[24:24]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2029(.Q(s_dvd[26:26]),.D(v_div_5[25:25]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2030(.Q(s_dvd[1:1]),.D(v_div_5[0:0]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2031(.Q(s_dvd[2:2]),.D(v_div_5[1:1]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2032(.Q(s_dvd[3:3]),.D(v_div_5[2:2]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2033(.Q(s_dvd[4:4]),.D(v_div_5[3:3]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2034(.Q(s_dvd[5:5]),.D(v_div_5[4:4]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2035(.Q(s_dvd[6:6]),.D(v_div_5[5:5]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2036(.Q(s_dvd[7:7]),.D(v_div_5[6:6]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2037(.Q(s_dvd[8:8]),.D(v_div_5[7:7]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2038(.Q(s_dvd[9:9]),.D(v_div_5[8:8]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2039(.Q(s_dvd[10:10]),.D(v_div_5[9:9]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2040(.Q(s_dvd[11:11]),.D(v_div_5[10:10]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2041(.Q(s_dvd[12:12]),.D(v_div_5[11:11]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2042(.Q(s_dvd[13:13]),.D(v_div_5[12:12]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  FDE desc2043(.Q(s_dvd[14:14]),.D(v_div_5[13:13]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O5));
  MUXCY desc2044(.DI(GND),.CI(un17_s_state_cry[23:23]),.S(un17_s_state_df25),.O(un17_s_state_cry[25:25]));
  LUT6 desc2045(.I0(s_dvdnd_i[26:26]),.I1(s_dvsor_i[0:0]),.I2(s_count[3:3]),.I3(s_count[1:1]),.I4(N_445),.I5(un17_s_state_cry[25:25]),.O(v_div_5_axb_0));
defparam desc2045.INIT=64'h0000A00033339333;
  LUT6_L desc2046(.I0(serial_div_qutnt[26:26]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_state),.I4(N_445),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[26:26]));
defparam desc2046.INIT=64'hAAAA2AAAAAAAEAAA;
  LUT6_L desc2047(.I0(serial_div_qutnt[2:2]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_state),.I4(N_452),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[2:2]));
defparam desc2047.INIT=64'hAAAA8AAAAAAABAAA;
  LUT6_L desc2048(.I0(serial_div_qutnt[18:18]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_state),.I4(N_445),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[18:18]));
defparam desc2048.INIT=64'hAAAA8AAAAAAABAAA;
  LUT6_L desc2049(.I0(serial_div_qutnt[0:0]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_state),.I4(N_452),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[0:0]));
defparam desc2049.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2050(.I0(serial_div_qutnt[16:16]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_state),.I4(N_445),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[16:16]));
defparam desc2050.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2051(.I0(serial_div_qutnt[14:14]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.LO(N_2635_i));
defparam desc2051.INIT=64'hAAAAAA8AAAAAAABA;
  LUT6_L desc2052(.I0(serial_div_qutnt[15:15]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.LO(N_2629_i));
defparam desc2052.INIT=64'hAAAA8AAAAAAABAAA;
  LUT6_L desc2053(.I0(serial_div_qutnt[6:6]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_448),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o_5_iv_i_i[6:6]));
defparam desc2053.INIT=64'hAAAAAA8AAAAAAABA;
  LUT6_L desc2054(.I0(serial_div_qutnt[7:7]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_448),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o_5_iv_i_i[7:7]));
defparam desc2054.INIT=64'hAAAA8AAAAAAABAAA;
  LUT6_L desc2055(.I0(serial_div_qutnt[12:12]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_count[0:0]),.I4(N_449),.I5(un17_s_state_cry[25:25]),.LO(N_2628_i));
defparam desc2055.INIT=64'hAAAAAAA2AAAAAAAE;
  LUT6_L desc2056(.I0(serial_div_qutnt[13:13]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_count[0:0]),.I4(N_449),.I5(un17_s_state_cry[25:25]),.LO(N_2634_i));
defparam desc2056.INIT=64'hAAAAA2AAAAAAAEAA;
  LUT6_L desc2057(.I0(serial_div_qutnt[20:20]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_447),.I5(un17_s_state_cry[25:25]),.LO(N_589_i));
defparam desc2057.INIT=64'hAAAAAA2AAAAAAAEA;
  LUT6 desc2058(.I0(s_dvdnd_i[38:38]),.I1(s_dvdnd_i[39:39]),.I2(s_dvdnd_i[44:44]),.I3(s_dvdnd_i[45:45]),.I4(N_2664_0_4),.I5(N_2664_1_4),.O(N_2664_1_0));
defparam desc2058.INIT=64'h0001000000000000;
  LUT6 desc2059(.I0(s_dvd[24:24]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.O(v_div_5_axb_24));
defparam desc2059.INIT=64'hAAAAAAA25555555D;
  LUT6 desc2060(.I0(s_dvd[25:25]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.O(v_div_5_axb_25));
defparam desc2060.INIT=64'hAAAAAAA25555555D;
  LUT6_L v_div_5_axb_26_cZ(.I0(s_dvd[26:26]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.LO(v_div_5_axb_26));
defparam v_div_5_axb_26_cZ.INIT=64'hAAAAAAA25555555D;
  LUT6_L desc2061(.I0(serial_div_qutnt[24:24]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_451),.I5(un17_s_state_cry[25:25]),.LO(N_2630_i));
defparam desc2061.INIT=64'hAAAAAAA2AAAAAAAE;
  LUT6_L desc2062(.I0(serial_div_qutnt[8:8]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_451),.I5(un17_s_state_cry[25:25]),.LO(N_2627_i));
defparam desc2062.INIT=64'hAAAAAAA8AAAAAAAB;
  LUT6_L desc2063(.I0(serial_div_qutnt[10:10]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.LO(N_2632_i));
defparam desc2063.INIT=64'hAAAAAAA8AAAAAAAB;
  LUT6 desc2064(.I0(s_dvdnd_i[27:27]),.I1(s_dvdnd_i[32:32]),.I2(s_dvdnd_i[33:33]),.I3(s_dvdnd_i[26:26]),.I4(N_2664_2_4),.I5(N_2664_3_4),.O(N_2664_2_0));
defparam desc2064.INIT=64'h0001000000000000;
  LUT6 desc2065(.I0(s_dvd[25:25]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_count[4:4]),.I4(s_count[2:2]),.I5(s_count[0:0]),.O(N_2621_i));
defparam desc2065.INIT=64'hAAAAAAAAAAAA2AAA;
  LUT6 desc2066(.I0(s_dvd[24:24]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_count[4:4]),.I4(s_count[2:2]),.I5(s_count[0:0]),.O(N_2620_i));
defparam desc2066.INIT=64'hAAAAAAAAAAAA2AAA;
  MUXCY_L v_div_5_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un17_s_state_cry_i[25:25]),.LO(v_div_5_cry_0_cy));
  LUT3_L s_ine_o_5_0_i_m2(.I0(fpu_op_i[0:0]),.I1(post_norm_div_ine),.I2(post_norm_mul_ine),.LO(N_504));
defparam s_ine_o_5_0_i_m2.INIT=8'hD8;
  LUT3_L m39_i_m2_cZ(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[1:1]),.I2(postnorm_addsub_output_o[1:1]),.LO(m39_i_m2));
defparam m39_i_m2_cZ.INIT=8'h27;
  LUT4 desc2067(.I0(s_dvsor_i[18:18]),.I1(s_dvsor_i[19:19]),.I2(s_dvsor_i[20:20]),.I3(s_dvsor_i[21:21]),.O(m112_i_4));
defparam desc2067.INIT=16'hFFFE;
  LUT4 desc2068(.I0(s_dvdnd_i[34:34]),.I1(s_dvdnd_i[35:35]),.I2(s_dvdnd_i[36:36]),.I3(s_dvdnd_i[37:37]),.O(N_2664_0_4));
defparam desc2068.INIT=16'h0001;
  LUT4 desc2069(.I0(s_dvdnd_i[40:40]),.I1(s_dvdnd_i[41:41]),.I2(s_dvdnd_i[42:42]),.I3(s_dvdnd_i[43:43]),.O(N_2664_1_4));
defparam desc2069.INIT=16'h0001;
  LUT4 desc2070(.I0(s_dvdnd_i[46:46]),.I1(s_dvdnd_i[47:47]),.I2(s_dvdnd_i[48:48]),.I3(s_dvdnd_i[49:49]),.O(N_2664_2_4));
defparam desc2070.INIT=16'h0001;
  LUT4 desc2071(.I0(s_dvdnd_i[28:28]),.I1(s_dvdnd_i[29:29]),.I2(s_dvdnd_i[30:30]),.I3(s_dvdnd_i[31:31]),.O(N_2664_3_4));
defparam desc2071.INIT=16'h0001;
  LUT6 desc2072(.I0(s_dvsor_i[13:13]),.I1(s_dvsor_i[14:14]),.I2(s_dvsor_i[15:15]),.I3(s_dvsor_i[16:16]),.I4(s_dvsor_i[17:17]),.I5(s_dvsor_i[23:23]),.O(m112_i_3));
defparam desc2072.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2073(.I0(s_dvsor_i[7:7]),.I1(s_dvsor_i[8:8]),.I2(s_dvsor_i[9:9]),.I3(s_dvsor_i[10:10]),.I4(s_dvsor_i[11:11]),.I5(s_dvsor_i[12:12]),.O(m112_i_2));
defparam desc2073.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2074(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(fpu_op_i[2:2]),.I3(s_dvsor_i[1:1]),.I4(s_dvsor_i[2:2]),.I5(s_dvsor_i[0:0]),.O(m112_i_0));
defparam desc2074.INIT=64'hFFFFFFFFFFFFFFF7;
  LUT5_L desc2075(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[31:31]),.I3(post_norm_mul_output[31:31]),.I4(N_500),.LO(N_564));
defparam desc2075.INIT=32'hC480F7B3;
  LUT5_L desc2076(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[30:30]),.I3(post_norm_mul_output[30:30]),.I4(N_499),.LO(N_563));
defparam desc2076.INIT=32'hC480F7B3;
  LUT5_L desc2077(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[29:29]),.I3(post_norm_mul_output[29:29]),.I4(N_498),.LO(N_562));
defparam desc2077.INIT=32'hC480F7B3;
  LUT5_L desc2078(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[28:28]),.I3(post_norm_mul_output[28:28]),.I4(N_497),.LO(N_561));
defparam desc2078.INIT=32'hC480F7B3;
  LUT5_L desc2079(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[27:27]),.I3(post_norm_mul_output[27:27]),.I4(N_496),.LO(N_560));
defparam desc2079.INIT=32'hC480F7B3;
  LUT5_L desc2080(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[26:26]),.I3(post_norm_mul_output[26:26]),.I4(N_495),.LO(N_559));
defparam desc2080.INIT=32'hC480F7B3;
  LUT5_L desc2081(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[25:25]),.I3(post_norm_mul_output[25:25]),.I4(N_494),.LO(N_558));
defparam desc2081.INIT=32'hC480F7B3;
  LUT5_L desc2082(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[24:24]),.I3(post_norm_mul_output[24:24]),.I4(N_493),.LO(N_557));
defparam desc2082.INIT=32'hC480F7B3;
  LUT5_L desc2083(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[23:23]),.I3(post_norm_mul_output[23:23]),.I4(N_492),.LO(N_556));
defparam desc2083.INIT=32'hC480F7B3;
  LUT5_L desc2084(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[22:22]),.I3(post_norm_mul_output[22:22]),.I4(N_491),.LO(N_555));
defparam desc2084.INIT=32'hC480F7B3;
  LUT5_L desc2085(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[21:21]),.I3(post_norm_mul_output[21:21]),.I4(N_490),.LO(N_554));
defparam desc2085.INIT=32'hC480F7B3;
  LUT5_L desc2086(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[20:20]),.I3(post_norm_mul_output[20:20]),.I4(N_489),.LO(N_553));
defparam desc2086.INIT=32'hC480F7B3;
  LUT5_L desc2087(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[19:19]),.I3(post_norm_mul_output[19:19]),.I4(N_488),.LO(N_552));
defparam desc2087.INIT=32'hC480F7B3;
  LUT5_L desc2088(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[18:18]),.I3(post_norm_mul_output[18:18]),.I4(N_487),.LO(N_551));
defparam desc2088.INIT=32'hC480F7B3;
  LUT5_L desc2089(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[17:17]),.I3(post_norm_mul_output[17:17]),.I4(N_486),.LO(N_550));
defparam desc2089.INIT=32'hC480F7B3;
  LUT5_L desc2090(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[16:16]),.I3(post_norm_mul_output[16:16]),.I4(N_485),.LO(N_549));
defparam desc2090.INIT=32'hC480F7B3;
  LUT5_L desc2091(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[15:15]),.I3(post_norm_mul_output[15:15]),.I4(N_484),.LO(N_548));
defparam desc2091.INIT=32'hC480F7B3;
  LUT5_L desc2092(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[14:14]),.I3(post_norm_mul_output[14:14]),.I4(N_483),.LO(N_547));
defparam desc2092.INIT=32'hC480F7B3;
  LUT5_L desc2093(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[13:13]),.I3(post_norm_mul_output[13:13]),.I4(N_482),.LO(N_546));
defparam desc2093.INIT=32'hC480F7B3;
  LUT5_L desc2094(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[12:12]),.I3(post_norm_mul_output[12:12]),.I4(N_481),.LO(N_545));
defparam desc2094.INIT=32'hC480F7B3;
  LUT5_L desc2095(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[11:11]),.I3(post_norm_mul_output[11:11]),.I4(m69_i_m2_lut6_2_O6),.LO(N_544));
defparam desc2095.INIT=32'hC480F7B3;
  LUT5_L desc2096(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[10:10]),.I3(post_norm_mul_output[10:10]),.I4(m57_i_m2_lut6_2_O5),.LO(N_543));
defparam desc2096.INIT=32'hC480F7B3;
  LUT5_L desc2097(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[9:9]),.I3(post_norm_mul_output[9:9]),.I4(N_2637_i_lut6_2_O5),.LO(N_542));
defparam desc2097.INIT=32'hC480F7B3;
  LUT5_L desc2098(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[8:8]),.I3(post_norm_mul_output[8:8]),.I4(m36_i_m2_lut6_2_O5),.LO(N_541));
defparam desc2098.INIT=32'hC480F7B3;
  LUT5_L desc2099(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[7:7]),.I3(post_norm_mul_output[7:7]),.I4(m57_i_m2_lut6_2_O6),.LO(s_output1_6_2_i_m2[7:7]));
defparam desc2099.INIT=32'hC480F7B3;
  LUT5_L desc2100(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[6:6]),.I3(post_norm_mul_output[6:6]),.I4(m54_i_m2_lut6_2_O6),.LO(s_output1_6_2_i_m2[6:6]));
defparam desc2100.INIT=32'hC480F7B3;
  LUT5_L desc2101(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[5:5]),.I3(post_norm_mul_output[5:5]),.I4(m51_i_m2_lut6_2_O6),.LO(N_538));
defparam desc2101.INIT=32'hC480F7B3;
  LUT5_L desc2102(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[4:4]),.I3(post_norm_mul_output[4:4]),.I4(m48_i_m2_lut6_2_O6),.LO(N_537));
defparam desc2102.INIT=32'hC480F7B3;
  LUT5_L desc2103(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[3:3]),.I3(post_norm_mul_output[3:3]),.I4(m45_i_m2_lut6_2_O6),.LO(N_536));
defparam desc2103.INIT=32'hC480F7B3;
  LUT5_L N_503_i_c(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[2:2]),.I3(post_norm_mul_output[2:2]),.I4(m42_i_m2_lut6_2_O6),.LO(N_503_i));
defparam N_503_i_c.INIT=32'hC480F7B3;
  LUT5_L N_502_i_c(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[1:1]),.I3(post_norm_mul_output[1:1]),.I4(m39_i_m2),.LO(N_502_i));
defparam N_502_i_c.INIT=32'hC480F7B3;
  LUT5_L N_501_i_c(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(post_norm_div_output[0:0]),.I3(post_norm_mul_output[0:0]),.I4(m36_i_m2_lut6_2_O6),.LO(N_501_i));
defparam N_501_i_c.INIT=32'hC480F7B3;
  LUT6_L desc2104(.I0(serial_div_qutnt[4:4]),.I1(s_count[0:0]),.I2(s_state),.I3(N_447),.I4(N_449),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[4:4]));
defparam desc2104.INIT=64'hAAAAAA8AAAAAAABA;
  LUT6_L desc2105(.I0(serial_div_qutnt[5:5]),.I1(s_count[0:0]),.I2(s_state),.I3(N_447),.I4(N_449),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[5:5]));
defparam desc2105.INIT=64'hAAAAAA2AAAAAAAEA;
  LUT6 desc2106(.I0(s_dvd[23:23]),.I1(s_dvdnd_i[49:49]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_616));
defparam desc2106.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2107(.I0(s_dvd[22:22]),.I1(s_dvdnd_i[48:48]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_615));
defparam desc2107.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2108(.I0(s_dvd[21:21]),.I1(s_dvdnd_i[47:47]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_614));
defparam desc2108.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2109(.I0(s_dvd[20:20]),.I1(s_dvdnd_i[46:46]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_613));
defparam desc2109.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2110(.I0(s_dvd[19:19]),.I1(s_dvdnd_i[45:45]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_612));
defparam desc2110.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2111(.I0(s_dvd[18:18]),.I1(s_dvdnd_i[44:44]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_611));
defparam desc2111.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2112(.I0(s_dvd[17:17]),.I1(s_dvdnd_i[43:43]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_610));
defparam desc2112.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2113(.I0(s_dvd[16:16]),.I1(s_dvdnd_i[42:42]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_609));
defparam desc2113.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2114(.I0(s_dvd[15:15]),.I1(s_dvdnd_i[41:41]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_608));
defparam desc2114.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2115(.I0(s_dvd[14:14]),.I1(s_dvdnd_i[40:40]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_607));
defparam desc2115.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2116(.I0(s_dvd[13:13]),.I1(s_dvdnd_i[39:39]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_606));
defparam desc2116.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2117(.I0(s_dvd[12:12]),.I1(s_dvdnd_i[38:38]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_605));
defparam desc2117.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2118(.I0(s_dvd[11:11]),.I1(s_dvdnd_i[37:37]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_604));
defparam desc2118.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2119(.I0(s_dvd[10:10]),.I1(s_dvdnd_i[36:36]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_603));
defparam desc2119.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2120(.I0(s_dvd[9:9]),.I1(s_dvdnd_i[35:35]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_602));
defparam desc2120.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2121(.I0(s_dvd[8:8]),.I1(s_dvdnd_i[34:34]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_601));
defparam desc2121.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2122(.I0(s_dvd[7:7]),.I1(s_dvdnd_i[33:33]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_600));
defparam desc2122.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2123(.I0(s_dvd[6:6]),.I1(s_dvdnd_i[32:32]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_599));
defparam desc2123.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2124(.I0(s_dvd[5:5]),.I1(s_dvdnd_i[31:31]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_598));
defparam desc2124.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2125(.I0(s_dvd[4:4]),.I1(s_dvdnd_i[30:30]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_597));
defparam desc2125.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2126(.I0(s_dvd[3:3]),.I1(s_dvdnd_i[29:29]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_596));
defparam desc2126.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2127(.I0(s_dvd[2:2]),.I1(s_dvdnd_i[28:28]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_595));
defparam desc2127.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 desc2128(.I0(s_dvd[1:1]),.I1(s_dvdnd_i[27:27]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_594));
defparam desc2128.INIT=64'hAAAAAAAAAAAAAACA;
  LUT6 un17_s_state_df25_RNO(.I0(s_dvd[26:26]),.I1(s_count[3:3]),.I2(s_count[1:1]),.I3(s_count[4:4]),.I4(s_count[2:2]),.I5(s_count[0:0]),.O(N_151_i));
defparam un17_s_state_df25_RNO.INIT=64'hAAAAAAAAAAAA2AAA;
  LUT6 desc2129(.I0(s_dvdnd_i[26:26]),.I1(s_dvsor_i[0:0]),.I2(s_count[4:4]),.I3(s_count[2:2]),.I4(s_count[0:0]),.I5(s_count_RNIQN9Q_O6[3:3]),.O(N_468_i));
defparam desc2129.INIT=64'h3333333333333393;
  LUT6_L desc2130(.I0(serial_div_qutnt[3:3]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_448),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o_5_iv_i_i[3:3]));
defparam desc2130.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2131(.I0(serial_div_qutnt[19:19]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_448),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o_5_iv_i_i[19:19]));
defparam desc2131.INIT=64'hAAAAA2AAAAAAAEAA;
  LUT6_L desc2132(.I0(serial_div_qutnt[21:21]),.I1(s_count[0:0]),.I2(s_state),.I3(N_447),.I4(N_453),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[21:21]));
defparam desc2132.INIT=64'hAAAAAA2AAAAAAAEA;
  LUT6_L desc2133(.I0(serial_div_qutnt[22:22]),.I1(s_count[0:0]),.I2(s_state),.I3(N_448),.I4(N_453),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[22:22]));
defparam desc2133.INIT=64'hAAAAAA8AAAAAAABA;
  LUT6_L desc2134(.I0(serial_div_qutnt[23:23]),.I1(s_count[0:0]),.I2(s_state),.I3(N_448),.I4(N_453),.I5(un17_s_state_cry[25:25]),.LO(s_qutnt_o[23:23]));
defparam desc2134.INIT=64'hAAAAAA2AAAAAAAEA;
  LUT6_L s_ine_o_5_0_i_m2_RNI9KOC1(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(fpu_op_i[2:2]),.I3(post_norm_sqrt_ine_o),.I4(postnorm_addsub_ine_o),.I5(N_504),.LO(s_ine_o_5));
defparam s_ine_o_5_0_i_m2_RNI9KOC1.INIT=64'h1F0F1C0C13031000;
  LUT6_L desc2135(.I0(serial_div_qutnt[17:17]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_447),.I5(un17_s_state_cry[25:25]),.LO(N_587_i));
defparam desc2135.INIT=64'hAAAAA2AAAAAAAEAA;
  LUT6_L desc2136(.I0(serial_div_qutnt[1:1]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_447),.I5(un17_s_state_cry[25:25]),.LO(N_584_i));
defparam desc2136.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2137(.I0(serial_div_qutnt[25:25]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_451),.I5(un17_s_state_cry[25:25]),.LO(i30_mux_i));
defparam desc2137.INIT=64'hAAAAA2AAAAAAAEAA;
  LUT6_L desc2138(.I0(serial_div_qutnt[11:11]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(s_count_RNIQN9Q_O6[3:3]),.I5(un17_s_state_cry[25:25]),.LO(N_2633_i));
defparam desc2138.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2139(.I0(serial_div_qutnt[9:9]),.I1(s_count[4:4]),.I2(s_count[2:2]),.I3(s_count[0:0]),.I4(N_451),.I5(un17_s_state_cry[25:25]),.LO(N_2631_i));
defparam desc2139.INIT=64'hAAAAA8AAAAAAABAA;
  LUT6_L desc2140(.I0(s_dvsor_i[3:3]),.I1(s_dvsor_i[4:4]),.I2(s_dvsor_i[5:5]),.I3(s_dvsor_i[6:6]),.I4(N_2664_1_0),.I5(N_2664_2_0),.LO(m112_i_1));
defparam desc2140.INIT=64'hFFFFFFFEFFFEFFFE;
  LUT6 desc2141(.I0(s_dvsor_i[22:22]),.I1(m112_i_0),.I2(m112_i_4),.I3(m112_i_2),.I4(m112_i_3),.I5(m112_i_1),.O(div_zero_o_0));
defparam desc2141.INIT=64'h0000000000000001;
  LUT2 v_div_5_cry_0_RNO_cZ(.I0(s_dvsor_i[0:0]),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_0_RNO));
defparam v_div_5_cry_0_RNO_cZ.INIT=4'h1;
  LUT2 v_div_5_cry_1_RNO_cZ(.I0(N_594),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_1_RNO));
defparam v_div_5_cry_1_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_2_RNO_cZ(.I0(N_595),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_2_RNO));
defparam v_div_5_cry_2_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_3_RNO_cZ(.I0(N_596),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_3_RNO));
defparam v_div_5_cry_3_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_4_RNO_cZ(.I0(N_597),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_4_RNO));
defparam v_div_5_cry_4_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_5_RNO_cZ(.I0(N_598),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_5_RNO));
defparam v_div_5_cry_5_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_6_RNO_cZ(.I0(N_599),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_6_RNO));
defparam v_div_5_cry_6_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_7_RNO_cZ(.I0(N_600),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_7_RNO));
defparam v_div_5_cry_7_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_8_RNO_cZ(.I0(N_601),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_8_RNO));
defparam v_div_5_cry_8_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_9_RNO_cZ(.I0(N_602),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_9_RNO));
defparam v_div_5_cry_9_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_10_RNO_cZ(.I0(N_603),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_10_RNO));
defparam v_div_5_cry_10_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_11_RNO_cZ(.I0(N_604),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_11_RNO));
defparam v_div_5_cry_11_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_12_RNO_cZ(.I0(N_605),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_12_RNO));
defparam v_div_5_cry_12_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_13_RNO_cZ(.I0(N_606),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_13_RNO));
defparam v_div_5_cry_13_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_14_RNO_cZ(.I0(N_607),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_14_RNO));
defparam v_div_5_cry_14_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_15_RNO_cZ(.I0(N_608),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_15_RNO));
defparam v_div_5_cry_15_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_16_RNO_cZ(.I0(N_609),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_16_RNO));
defparam v_div_5_cry_16_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_17_RNO_cZ(.I0(N_610),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_17_RNO));
defparam v_div_5_cry_17_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_18_RNO_cZ(.I0(N_611),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_18_RNO));
defparam v_div_5_cry_18_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_19_RNO_cZ(.I0(N_612),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_19_RNO));
defparam v_div_5_cry_19_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_20_RNO_cZ(.I0(N_613),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_20_RNO));
defparam v_div_5_cry_20_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_21_RNO_cZ(.I0(N_614),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_21_RNO));
defparam v_div_5_cry_21_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_22_RNO_cZ(.I0(N_615),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_22_RNO));
defparam v_div_5_cry_22_RNO_cZ.INIT=4'h2;
  LUT2 v_div_5_cry_23_RNO_cZ(.I0(N_616),.I1(un17_s_state_cry[25:25]),.O(v_div_5_cry_23_RNO));
defparam v_div_5_cry_23_RNO_cZ.INIT=4'h2;
  XORCY v_div_5_s_26(.LI(v_div_5_axb_26),.CI(v_div_5_cry_25),.O(v_div_5[26:26]));
  XORCY v_div_5_s_25(.LI(v_div_5_axb_25),.CI(v_div_5_cry_24),.O(v_div_5[25:25]));
  MUXCY_L v_div_5_cry_25_cZ(.DI(N_2621_i),.CI(v_div_5_cry_24),.S(v_div_5_axb_25),.LO(v_div_5_cry_25));
  XORCY v_div_5_s_24(.LI(v_div_5_axb_24),.CI(v_div_5_cry_23),.O(v_div_5[24:24]));
  MUXCY_L v_div_5_cry_24_cZ(.DI(N_2620_i),.CI(v_div_5_cry_23),.S(v_div_5_axb_24),.LO(v_div_5_cry_24));
  XORCY v_div_5_s_23(.LI(v_div_5_axb_23),.CI(v_div_5_cry_22),.O(v_div_5[23:23]));
  MUXCY_L v_div_5_cry_23_cZ(.DI(v_div_5_cry_23_RNO),.CI(v_div_5_cry_22),.S(v_div_5_axb_23),.LO(v_div_5_cry_23));
  XORCY v_div_5_s_22(.LI(v_div_5_axb_22),.CI(v_div_5_cry_21),.O(v_div_5[22:22]));
  MUXCY_L v_div_5_cry_22_cZ(.DI(v_div_5_cry_22_RNO),.CI(v_div_5_cry_21),.S(v_div_5_axb_22),.LO(v_div_5_cry_22));
  XORCY v_div_5_s_21(.LI(v_div_5_axb_21),.CI(v_div_5_cry_20),.O(v_div_5[21:21]));
  MUXCY_L v_div_5_cry_21_cZ(.DI(v_div_5_cry_21_RNO),.CI(v_div_5_cry_20),.S(v_div_5_axb_21),.LO(v_div_5_cry_21));
  XORCY v_div_5_s_20(.LI(v_div_5_axb_20),.CI(v_div_5_cry_19),.O(v_div_5[20:20]));
  MUXCY_L v_div_5_cry_20_cZ(.DI(v_div_5_cry_20_RNO),.CI(v_div_5_cry_19),.S(v_div_5_axb_20),.LO(v_div_5_cry_20));
  XORCY v_div_5_s_19(.LI(v_div_5_axb_19),.CI(v_div_5_cry_18),.O(v_div_5[19:19]));
  MUXCY_L v_div_5_cry_19_cZ(.DI(v_div_5_cry_19_RNO),.CI(v_div_5_cry_18),.S(v_div_5_axb_19),.LO(v_div_5_cry_19));
  XORCY v_div_5_s_18(.LI(v_div_5_axb_18),.CI(v_div_5_cry_17),.O(v_div_5[18:18]));
  MUXCY_L v_div_5_cry_18_cZ(.DI(v_div_5_cry_18_RNO),.CI(v_div_5_cry_17),.S(v_div_5_axb_18),.LO(v_div_5_cry_18));
  XORCY v_div_5_s_17(.LI(v_div_5_axb_17),.CI(v_div_5_cry_16),.O(v_div_5[17:17]));
  MUXCY_L v_div_5_cry_17_cZ(.DI(v_div_5_cry_17_RNO),.CI(v_div_5_cry_16),.S(v_div_5_axb_17),.LO(v_div_5_cry_17));
  XORCY v_div_5_s_16(.LI(v_div_5_axb_16),.CI(v_div_5_cry_15),.O(v_div_5[16:16]));
  MUXCY_L v_div_5_cry_16_cZ(.DI(v_div_5_cry_16_RNO),.CI(v_div_5_cry_15),.S(v_div_5_axb_16),.LO(v_div_5_cry_16));
  XORCY v_div_5_s_15(.LI(v_div_5_axb_15),.CI(v_div_5_cry_14),.O(v_div_5[15:15]));
  MUXCY_L v_div_5_cry_15_cZ(.DI(v_div_5_cry_15_RNO),.CI(v_div_5_cry_14),.S(v_div_5_axb_15),.LO(v_div_5_cry_15));
  XORCY v_div_5_s_14(.LI(v_div_5_axb_14),.CI(v_div_5_cry_13),.O(v_div_5[14:14]));
  MUXCY_L v_div_5_cry_14_cZ(.DI(v_div_5_cry_14_RNO),.CI(v_div_5_cry_13),.S(v_div_5_axb_14),.LO(v_div_5_cry_14));
  XORCY v_div_5_s_13(.LI(v_div_5_axb_13),.CI(v_div_5_cry_12),.O(v_div_5[13:13]));
  MUXCY_L v_div_5_cry_13_cZ(.DI(v_div_5_cry_13_RNO),.CI(v_div_5_cry_12),.S(v_div_5_axb_13),.LO(v_div_5_cry_13));
  XORCY v_div_5_s_12(.LI(v_div_5_axb_12),.CI(v_div_5_cry_11),.O(v_div_5[12:12]));
  MUXCY_L v_div_5_cry_12_cZ(.DI(v_div_5_cry_12_RNO),.CI(v_div_5_cry_11),.S(v_div_5_axb_12),.LO(v_div_5_cry_12));
  XORCY v_div_5_s_11(.LI(v_div_5_axb_11),.CI(v_div_5_cry_10),.O(v_div_5[11:11]));
  MUXCY_L v_div_5_cry_11_cZ(.DI(v_div_5_cry_11_RNO),.CI(v_div_5_cry_10),.S(v_div_5_axb_11),.LO(v_div_5_cry_11));
  XORCY v_div_5_s_10(.LI(v_div_5_axb_10),.CI(v_div_5_cry_9),.O(v_div_5[10:10]));
  MUXCY_L v_div_5_cry_10_cZ(.DI(v_div_5_cry_10_RNO),.CI(v_div_5_cry_9),.S(v_div_5_axb_10),.LO(v_div_5_cry_10));
  XORCY v_div_5_s_9(.LI(v_div_5_axb_9),.CI(v_div_5_cry_8),.O(v_div_5[9:9]));
  MUXCY_L v_div_5_cry_9_cZ(.DI(v_div_5_cry_9_RNO),.CI(v_div_5_cry_8),.S(v_div_5_axb_9),.LO(v_div_5_cry_9));
  XORCY v_div_5_s_8(.LI(v_div_5_axb_8),.CI(v_div_5_cry_7),.O(v_div_5[8:8]));
  MUXCY_L v_div_5_cry_8_cZ(.DI(v_div_5_cry_8_RNO),.CI(v_div_5_cry_7),.S(v_div_5_axb_8),.LO(v_div_5_cry_8));
  XORCY v_div_5_s_7(.LI(v_div_5_axb_7),.CI(v_div_5_cry_6),.O(v_div_5[7:7]));
  MUXCY_L v_div_5_cry_7_cZ(.DI(v_div_5_cry_7_RNO),.CI(v_div_5_cry_6),.S(v_div_5_axb_7),.LO(v_div_5_cry_7));
  XORCY v_div_5_s_6(.LI(v_div_5_axb_6),.CI(v_div_5_cry_5),.O(v_div_5[6:6]));
  MUXCY_L v_div_5_cry_6_cZ(.DI(v_div_5_cry_6_RNO),.CI(v_div_5_cry_5),.S(v_div_5_axb_6),.LO(v_div_5_cry_6));
  XORCY v_div_5_s_5(.LI(v_div_5_axb_5),.CI(v_div_5_cry_4),.O(v_div_5[5:5]));
  MUXCY_L v_div_5_cry_5_cZ(.DI(v_div_5_cry_5_RNO),.CI(v_div_5_cry_4),.S(v_div_5_axb_5),.LO(v_div_5_cry_5));
  XORCY v_div_5_s_4(.LI(v_div_5_axb_4),.CI(v_div_5_cry_3),.O(v_div_5[4:4]));
  MUXCY_L v_div_5_cry_4_cZ(.DI(v_div_5_cry_4_RNO),.CI(v_div_5_cry_3),.S(v_div_5_axb_4),.LO(v_div_5_cry_4));
  XORCY v_div_5_s_3(.LI(v_div_5_axb_3),.CI(v_div_5_cry_2),.O(v_div_5[3:3]));
  MUXCY_L v_div_5_cry_3_cZ(.DI(v_div_5_cry_3_RNO),.CI(v_div_5_cry_2),.S(v_div_5_axb_3),.LO(v_div_5_cry_3));
  XORCY v_div_5_s_2(.LI(v_div_5_axb_2),.CI(v_div_5_cry_1),.O(v_div_5[2:2]));
  MUXCY_L v_div_5_cry_2_cZ(.DI(v_div_5_cry_2_RNO),.CI(v_div_5_cry_1),.S(v_div_5_axb_2),.LO(v_div_5_cry_2));
  XORCY v_div_5_s_1(.LI(v_div_5_axb_1),.CI(v_div_5_cry_0),.O(v_div_5[1:1]));
  MUXCY_L v_div_5_cry_1_cZ(.DI(v_div_5_cry_1_RNO),.CI(v_div_5_cry_0),.S(v_div_5_axb_1),.LO(v_div_5_cry_1));
  XORCY v_div_5_s_0(.LI(v_div_5_axb_0),.CI(v_div_5_cry_0_cy),.O(v_div_5[0:0]));
  MUXCY_L v_div_5_cry_0_cZ(.DI(v_div_5_cry_0_RNO),.CI(v_div_5_cry_0_cy),.S(v_div_5_axb_0),.LO(v_div_5_cry_0));
  FDRE desc2142(.Q(serial_div_rmndr[7:7]),.D(v_div_5[7:7]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2143(.Q(serial_div_rmndr[6:6]),.D(v_div_5[6:6]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2144(.Q(serial_div_rmndr[5:5]),.D(v_div_5[5:5]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2145(.Q(serial_div_rmndr[4:4]),.D(v_div_5[4:4]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2146(.Q(serial_div_rmndr[3:3]),.D(v_div_5[3:3]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2147(.Q(serial_div_rmndr[2:2]),.D(v_div_5[2:2]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2148(.Q(serial_div_rmndr[1:1]),.D(v_div_5[1:1]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2149(.Q(serial_div_rmndr[0:0]),.D(v_div_5[0:0]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2150(.Q(serial_div_rmndr[22:22]),.D(v_div_5[22:22]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2151(.Q(serial_div_rmndr[21:21]),.D(v_div_5[21:21]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2152(.Q(serial_div_rmndr[20:20]),.D(v_div_5[20:20]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2153(.Q(serial_div_rmndr[19:19]),.D(v_div_5[19:19]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2154(.Q(serial_div_rmndr[18:18]),.D(v_div_5[18:18]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2155(.Q(serial_div_rmndr[17:17]),.D(v_div_5[17:17]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2156(.Q(serial_div_rmndr[16:16]),.D(v_div_5[16:16]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2157(.Q(serial_div_rmndr[15:15]),.D(v_div_5[15:15]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2158(.Q(serial_div_rmndr[14:14]),.D(v_div_5[14:14]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2159(.Q(serial_div_rmndr[13:13]),.D(v_div_5[13:13]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2160(.Q(serial_div_rmndr[12:12]),.D(v_div_5[12:12]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2161(.Q(serial_div_rmndr[11:11]),.D(v_div_5[11:11]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2162(.Q(serial_div_rmndr[10:10]),.D(v_div_5[10:10]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2163(.Q(serial_div_rmndr[9:9]),.D(v_div_5[9:9]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2164(.Q(serial_div_rmndr[8:8]),.D(v_div_5[8:8]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2165(.Q(serial_div_rmndr[26:26]),.D(v_div_5[26:26]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2166(.Q(serial_div_rmndr[25:25]),.D(v_div_5[25:25]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2167(.Q(serial_div_rmndr[24:24]),.D(v_div_5[24:24]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2168(.Q(serial_div_rmndr[23:23]),.D(v_div_5[23:23]),.C(clk_i),.R(s_start_i),.CE(s_state));
  MUXCY_L desc2169(.DI(un17_s_state_lt23),.CI(un17_s_state_cry[21:21]),.S(un17_s_state_df23),.LO(un17_s_state_cry[23:23]));
  MUXCY_L desc2170(.DI(un17_s_state_lt21),.CI(un17_s_state_cry[19:19]),.S(un17_s_state_df21),.LO(un17_s_state_cry[21:21]));
  MUXCY_L desc2171(.DI(un17_s_state_lt19),.CI(un17_s_state_cry[17:17]),.S(un17_s_state_df19),.LO(un17_s_state_cry[19:19]));
  MUXCY_L desc2172(.DI(un17_s_state_lt17),.CI(un17_s_state_cry[15:15]),.S(un17_s_state_df17),.LO(un17_s_state_cry[17:17]));
  MUXCY_L desc2173(.DI(un17_s_state_lt15),.CI(un17_s_state_cry[13:13]),.S(un17_s_state_df15),.LO(un17_s_state_cry[15:15]));
  MUXCY_L desc2174(.DI(un17_s_state_lt13),.CI(un17_s_state_cry[11:11]),.S(un17_s_state_df13),.LO(un17_s_state_cry[13:13]));
  MUXCY_L desc2175(.DI(un17_s_state_lt11),.CI(un17_s_state_cry[9:9]),.S(un17_s_state_df11),.LO(un17_s_state_cry[11:11]));
  MUXCY_L desc2176(.DI(un17_s_state_lt9),.CI(un17_s_state_cry[7:7]),.S(un17_s_state_df9),.LO(un17_s_state_cry[9:9]));
  MUXCY_L desc2177(.DI(un17_s_state_lt7),.CI(un17_s_state_cry[5:5]),.S(un17_s_state_df7),.LO(un17_s_state_cry[7:7]));
  MUXCY_L desc2178(.DI(un17_s_state_lt5),.CI(un17_s_state_cry[3:3]),.S(un17_s_state_df5),.LO(un17_s_state_cry[5:5]));
  MUXCY_L desc2179(.DI(un17_s_state_lt3),.CI(un17_s_state_cry[1:1]),.S(un17_s_state_df3),.LO(un17_s_state_cry[3:3]));
  MUXCY_L desc2180(.DI(un17_s_state_lt1),.CI(un17_s_state_cry[0:0]),.S(un17_s_state_df1),.LO(un17_s_state_cry[1:1]));
  MUXCY_L desc2181(.DI(s_dvsor_i[0:0]),.CI(GND),.S(N_468_i),.LO(un17_s_state_cry[0:0]));
  FDRE desc2182(.Q(serial_div_qutnt[25:25]),.D(i30_mux_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2183(.Q(serial_div_qutnt[24:24]),.D(N_2630_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2184(.Q(serial_div_qutnt[20:20]),.D(N_589_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2185(.Q(serial_div_qutnt[19:19]),.D(s_qutnt_o_5_iv_i_i[19:19]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2186(.Q(serial_div_qutnt[17:17]),.D(N_587_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2187(.Q(serial_div_qutnt[15:15]),.D(N_2629_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2188(.Q(serial_div_qutnt[14:14]),.D(N_2635_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2189(.Q(serial_div_qutnt[13:13]),.D(N_2634_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2190(.Q(serial_div_qutnt[12:12]),.D(N_2628_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2191(.Q(serial_div_qutnt[11:11]),.D(N_2633_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2192(.Q(serial_div_qutnt[10:10]),.D(N_2632_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2193(.Q(serial_div_qutnt[9:9]),.D(N_2631_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2194(.Q(serial_div_qutnt[8:8]),.D(N_2627_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2195(.Q(serial_div_qutnt[7:7]),.D(s_qutnt_o_5_iv_i_i[7:7]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2196(.Q(serial_div_qutnt[6:6]),.D(s_qutnt_o_5_iv_i_i[6:6]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2197(.Q(serial_div_qutnt[3:3]),.D(s_qutnt_o_5_iv_i_i[3:3]),.C(clk_i),.R(s_start_i),.CE(s_state));
  FDRE desc2198(.Q(serial_div_qutnt[1:1]),.D(N_584_i),.C(clk_i),.R(s_start_i),.CE(s_state));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT5 desc2199(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_1491_i));
defparam desc2199.INIT=32'hE1E1E1E0;
  LUT4 desc2200(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.O(N_237_i));
defparam desc2200.INIT=16'hFE01;
  LUT5 desc2201(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_1490_i));
defparam desc2201.INIT=32'h55555554;
  LUT5 desc2202(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_239_i));
defparam desc2202.INIT=32'hFFFE0001;
  LUT2 desc2203(.I0(s_count[4:4]),.I1(s_count[2:2]),.O(N_449));
defparam desc2203.INIT=4'hB;
  LUT5 desc2204(.I0(N_447),.I1(s_count[0:0]),.I2(s_state),.I3(s_count[4:4]),.I4(s_count[2:2]),.O(N_1489_i_0));
defparam desc2204.INIT=32'hF0F0F0E0;
  LUT2 desc2205(.I0(s_count[3:3]),.I1(s_count[1:1]),.O(N_447));
defparam desc2205.INIT=4'hE;
  LUT2 desc2206(.I0(s_count[3:3]),.I1(s_count[1:1]),.O(N_448));
defparam desc2206.INIT=4'hB;
  LUT2 desc2207(.I0(s_count[3:3]),.I1(s_count[1:1]),.O(s_count_RNIQN9Q_O6[3:3]));
defparam desc2207.INIT=4'h7;
  LUT2 desc2208(.I0(s_count[3:3]),.I1(s_count[1:1]),.O(N_451));
defparam desc2208.INIT=4'hD;
  LUT3 m117_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[27:27]),.I2(post_norm_sqrt_output[27:27]),.O(N_496));
defparam m117_i_m2_lut6_2_o6.INIT=8'h1B;
  LUT3 m117_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[31:31]),.I2(postnorm_addsub_output_o[31:31]),.O(N_500));
defparam m117_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m99_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[21:21]),.I2(postnorm_addsub_output_o[21:21]),.O(N_490));
defparam m99_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m99_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[24:24]),.I2(post_norm_sqrt_output[24:24]),.O(N_493));
defparam m99_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m96_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[20:20]),.I2(postnorm_addsub_output_o[20:20]),.O(N_489));
defparam m96_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m96_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[26:26]),.I2(post_norm_sqrt_output[26:26]),.O(N_495));
defparam m96_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m93_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[19:19]),.I2(postnorm_addsub_output_o[19:19]),.O(N_488));
defparam m93_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m93_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[29:29]),.I2(post_norm_sqrt_output[29:29]),.O(N_498));
defparam m93_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m78_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[14:14]),.I2(postnorm_addsub_output_o[14:14]),.O(N_483));
defparam m78_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m78_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[17:17]),.I2(postnorm_addsub_output_o[17:17]),.O(N_486));
defparam m78_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m75_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[13:13]),.I2(postnorm_addsub_output_o[13:13]),.O(N_482));
defparam m75_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m75_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[18:18]),.I2(postnorm_addsub_output_o[18:18]),.O(N_487));
defparam m75_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m72_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[12:12]),.I2(postnorm_addsub_output_o[12:12]),.O(N_481));
defparam m72_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m72_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[22:22]),.I2(postnorm_addsub_output_o[22:22]),.O(N_491));
defparam m72_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m69_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[11:11]),.I2(postnorm_addsub_output_o[11:11]),.O(m69_i_m2_lut6_2_O6));
defparam m69_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m69_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[30:30]),.I2(post_norm_sqrt_output[30:30]),.O(N_499));
defparam m69_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m57_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[7:7]),.I2(postnorm_addsub_output_o[7:7]),.O(m57_i_m2_lut6_2_O6));
defparam m57_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m57_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[10:10]),.I2(postnorm_addsub_output_o[10:10]),.O(m57_i_m2_lut6_2_O5));
defparam m57_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m54_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[6:6]),.I2(postnorm_addsub_output_o[6:6]),.O(m54_i_m2_lut6_2_O6));
defparam m54_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m54_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[15:15]),.I2(postnorm_addsub_output_o[15:15]),.O(N_484));
defparam m54_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m51_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[5:5]),.I2(postnorm_addsub_output_o[5:5]),.O(m51_i_m2_lut6_2_O6));
defparam m51_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m51_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[16:16]),.I2(postnorm_addsub_output_o[16:16]),.O(N_485));
defparam m51_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 m48_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[4:4]),.I2(postnorm_addsub_output_o[4:4]),.O(m48_i_m2_lut6_2_O6));
defparam m48_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m48_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[23:23]),.I2(post_norm_sqrt_output[23:23]),.O(N_492));
defparam m48_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m45_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[3:3]),.I2(postnorm_addsub_output_o[3:3]),.O(m45_i_m2_lut6_2_O6));
defparam m45_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m45_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[25:25]),.I2(post_norm_sqrt_output[25:25]),.O(N_494));
defparam m45_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m42_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[2:2]),.I2(postnorm_addsub_output_o[2:2]),.O(m42_i_m2_lut6_2_O6));
defparam m42_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m42_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(postnorm_addsub_output_o[28:28]),.I2(post_norm_sqrt_output[28:28]),.O(N_497));
defparam m42_i_m2_lut6_2_o5.INIT=8'h1B;
  LUT3 m36_i_m2_lut6_2_o6(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[0:0]),.I2(postnorm_addsub_output_o[0:0]),.O(m36_i_m2_lut6_2_O6));
defparam m36_i_m2_lut6_2_o6.INIT=8'h27;
  LUT3 m36_i_m2_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[8:8]),.I2(postnorm_addsub_output_o[8:8]),.O(m36_i_m2_lut6_2_O5));
defparam m36_i_m2_lut6_2_o5.INIT=8'h27;
  LUT3 desc2209(.I0(s_count[4:4]),.I1(s_count[2:2]),.I2(s_count[0:0]),.O(N_452));
defparam desc2209.INIT=8'hFE;
  LUT2 desc2210(.I0(s_count[1:1]),.I1(s_count[0:0]),.O(N_466_i_i));
defparam desc2210.INIT=4'h9;
  LUT3 desc2211(.I0(s_count[4:4]),.I1(s_count[2:2]),.I2(s_count[0:0]),.O(N_445));
defparam desc2211.INIT=8'hFD;
  LUT2 desc2212(.I0(s_count[4:4]),.I1(s_count[2:2]),.O(N_453));
defparam desc2212.INIT=4'h7;
  LUT3 N_2637_i_lut6_2_o6(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(fpu_op_i[2:2]),.O(N_2637_i));
defparam N_2637_i_lut6_2_o6.INIT=8'hE0;
  LUT3 N_2637_i_lut6_2_o5(.I0(fpu_op_i[2:2]),.I1(post_norm_sqrt_output[9:9]),.I2(postnorm_addsub_output_o[9:9]),.O(N_2637_i_lut6_2_O5));
defparam N_2637_i_lut6_2_o5.INIT=8'h27;
  LUT3 un17_s_state_df23_lut6_2_o6(.I0(s_dvsor_i[23:23]),.I1(N_2620_i),.I2(N_616),.O(un17_s_state_df23));
defparam un17_s_state_df23_lut6_2_o6.INIT=8'h21;
  LUT3 un17_s_state_df23_lut6_2_o5(.I0(s_dvsor_i[23:23]),.I1(N_2620_i),.I2(N_616),.O(un17_s_state_lt23));
defparam un17_s_state_df23_lut6_2_o5.INIT=8'h02;
  LUT4 un17_s_state_df21_lut6_2_o6(.I0(s_dvsor_i[21:21]),.I1(s_dvsor_i[22:22]),.I2(N_614),.I3(N_615),.O(un17_s_state_df21));
defparam un17_s_state_df21_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df21_lut6_2_o5(.I0(s_dvsor_i[21:21]),.I1(s_dvsor_i[22:22]),.I2(N_614),.I3(N_615),.O(un17_s_state_lt21));
defparam un17_s_state_df21_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df19_lut6_2_o6(.I0(s_dvsor_i[19:19]),.I1(s_dvsor_i[20:20]),.I2(N_612),.I3(N_613),.O(un17_s_state_df19));
defparam un17_s_state_df19_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df19_lut6_2_o5(.I0(s_dvsor_i[19:19]),.I1(s_dvsor_i[20:20]),.I2(N_612),.I3(N_613),.O(un17_s_state_lt19));
defparam un17_s_state_df19_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df17_lut6_2_o6(.I0(s_dvsor_i[17:17]),.I1(s_dvsor_i[18:18]),.I2(N_610),.I3(N_611),.O(un17_s_state_df17));
defparam un17_s_state_df17_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df17_lut6_2_o5(.I0(s_dvsor_i[17:17]),.I1(s_dvsor_i[18:18]),.I2(N_610),.I3(N_611),.O(un17_s_state_lt17));
defparam un17_s_state_df17_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df15_lut6_2_o6(.I0(s_dvsor_i[15:15]),.I1(s_dvsor_i[16:16]),.I2(N_608),.I3(N_609),.O(un17_s_state_df15));
defparam un17_s_state_df15_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df15_lut6_2_o5(.I0(s_dvsor_i[15:15]),.I1(s_dvsor_i[16:16]),.I2(N_608),.I3(N_609),.O(un17_s_state_lt15));
defparam un17_s_state_df15_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df13_lut6_2_o6(.I0(s_dvsor_i[13:13]),.I1(s_dvsor_i[14:14]),.I2(N_606),.I3(N_607),.O(un17_s_state_df13));
defparam un17_s_state_df13_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df13_lut6_2_o5(.I0(s_dvsor_i[13:13]),.I1(s_dvsor_i[14:14]),.I2(N_606),.I3(N_607),.O(un17_s_state_lt13));
defparam un17_s_state_df13_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df11_lut6_2_o6(.I0(s_dvsor_i[11:11]),.I1(s_dvsor_i[12:12]),.I2(N_604),.I3(N_605),.O(un17_s_state_df11));
defparam un17_s_state_df11_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df11_lut6_2_o5(.I0(s_dvsor_i[11:11]),.I1(s_dvsor_i[12:12]),.I2(N_604),.I3(N_605),.O(un17_s_state_lt11));
defparam un17_s_state_df11_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df9_lut6_2_o6(.I0(s_dvsor_i[9:9]),.I1(s_dvsor_i[10:10]),.I2(N_602),.I3(N_603),.O(un17_s_state_df9));
defparam un17_s_state_df9_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df9_lut6_2_o5(.I0(s_dvsor_i[9:9]),.I1(s_dvsor_i[10:10]),.I2(N_602),.I3(N_603),.O(un17_s_state_lt9));
defparam un17_s_state_df9_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df7_lut6_2_o6(.I0(s_dvsor_i[7:7]),.I1(s_dvsor_i[8:8]),.I2(N_600),.I3(N_601),.O(un17_s_state_df7));
defparam un17_s_state_df7_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df7_lut6_2_o5(.I0(s_dvsor_i[7:7]),.I1(s_dvsor_i[8:8]),.I2(N_600),.I3(N_601),.O(un17_s_state_lt7));
defparam un17_s_state_df7_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df5_lut6_2_o6(.I0(s_dvsor_i[6:6]),.I1(s_dvsor_i[5:5]),.I2(N_598),.I3(N_599),.O(un17_s_state_df5));
defparam un17_s_state_df5_lut6_2_o6.INIT=16'h8241;
  LUT4 un17_s_state_df5_lut6_2_o5(.I0(s_dvsor_i[6:6]),.I1(s_dvsor_i[5:5]),.I2(N_598),.I3(N_599),.O(un17_s_state_lt5));
defparam un17_s_state_df5_lut6_2_o5.INIT=16'h08AE;
  LUT4 un17_s_state_df3_lut6_2_o6(.I0(s_dvsor_i[3:3]),.I1(s_dvsor_i[4:4]),.I2(N_596),.I3(N_597),.O(un17_s_state_df3));
defparam un17_s_state_df3_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df3_lut6_2_o5(.I0(s_dvsor_i[3:3]),.I1(s_dvsor_i[4:4]),.I2(N_596),.I3(N_597),.O(un17_s_state_lt3));
defparam un17_s_state_df3_lut6_2_o5.INIT=16'h08CE;
  LUT4 un17_s_state_df1_lut6_2_o6(.I0(s_dvsor_i[1:1]),.I1(s_dvsor_i[2:2]),.I2(N_594),.I3(N_595),.O(un17_s_state_df1));
defparam un17_s_state_df1_lut6_2_o6.INIT=16'h8421;
  LUT4 un17_s_state_df1_lut6_2_o5(.I0(s_dvsor_i[1:1]),.I1(s_dvsor_i[2:2]),.I2(N_594),.I3(N_595),.O(un17_s_state_lt1));
defparam un17_s_state_df1_lut6_2_o5.INIT=16'h08CE;
endmodule
module post_norm_div_inj (un11_s_exp_10_o_0,s_opb_i_4,s_opb_i_5,s_opb_i_6,s_opb_i_7,s_opb_i_1,s_opb_i_2,s_opb_i_3,s_opb_i_0,s_opa_i_1,s_opa_i_2,s_opa_i_3,s_opa_i_4,s_opa_i_5,s_opa_i_6,s_opa_i_7,s_opa_i_0,serial_div_rmndr,serial_div_qutnt,s_rmode_i,s_rmode_i_0,s_fractb_i,s_fracta_i,post_norm_div_output,clk_i,un11_s_exp_10_o_axb_0_i,s_infb,un1_s_infa,result_4,N_1942_i,post_norm_div_ine,result_5,result_3_21_1,result_3_21_3,result_11,un1_s_nan_a,un1_s_nan_b,un3_s_op_0);
input [9:1] un11_s_exp_10_o_0 ;
output s_opb_i_4 ;
output s_opb_i_5 ;
output s_opb_i_6 ;
output s_opb_i_7 ;
output s_opb_i_1 ;
output s_opb_i_2 ;
output s_opb_i_3 ;
input [30:23] s_opb_i_0 ;
output s_opa_i_1 ;
output s_opa_i_2 ;
output s_opa_i_3 ;
output s_opa_i_4 ;
output s_opa_i_5 ;
output s_opa_i_6 ;
output s_opa_i_7 ;
input [30:23] s_opa_i_0 ;
input [26:0] serial_div_rmndr ;
input [26:0] serial_div_qutnt ;
output [1:0] s_rmode_i ;
input [1:0] s_rmode_i_0 ;
input [22:0] s_fractb_i ;
input [22:16] s_fracta_i ;
output [31:0] post_norm_div_output ;
input clk_i ;
input un11_s_exp_10_o_axb_0_i ;
output s_infb ;
output un1_s_infa ;
output result_4 ;
input N_1942_i ;
output post_norm_div_ine ;
output result_5 ;
input result_3_21_1 ;
input result_3_21_3 ;
input result_11 ;
output un1_s_nan_a ;
output un1_s_nan_b ;
output un3_s_op_0 ;
wire s_opb_i_4 ;
wire s_opb_i_5 ;
wire s_opb_i_6 ;
wire s_opb_i_7 ;
wire s_opb_i_1 ;
wire s_opb_i_2 ;
wire s_opb_i_3 ;
wire s_opa_i_1 ;
wire s_opa_i_2 ;
wire s_opa_i_3 ;
wire s_opa_i_4 ;
wire s_opa_i_5 ;
wire s_opa_i_6 ;
wire s_opa_i_7 ;
wire clk_i ;
wire un11_s_exp_10_o_axb_0_i ;
wire s_infb ;
wire un1_s_infa ;
wire result_4 ;
wire N_1942_i ;
wire post_norm_div_ine ;
wire result_5 ;
wire result_3_21_1 ;
wire result_3_21_3 ;
wire result_11 ;
wire un1_s_nan_a ;
wire un1_s_nan_b ;
wire un3_s_op_0 ;
wire s_exp_10_i_8_tmp_d_array_0 ;
wire s_exp_10_i_7_tmp_d_array_0 ;
wire s_exp_10_i_6_tmp_d_array_0 ;
wire s_exp_10_i_5_tmp_d_array_0 ;
wire s_exp_10_i_4_tmp_d_array_0 ;
wire s_exp_10_i_3_tmp_d_array_0 ;
wire s_exp_10_i_2_tmp_d_array_0 ;
wire s_exp_10_i_1_tmp_d_array_0 ;
wire s_exp_10_i_0_tmp_d_array_0 ;
wire s_exp_10_i_tmp_d_array_0 ;
wire [9:0] s_exp_10_i ;
wire [6:0] v_shr_2 ;
wire [9:1] s_exp_10b ;
wire [26:0] s_fraco1 ;
wire [22:1] un6_s_frac_rnd1 ;
wire [22:0] s_frac_rnd ;
wire [8:0] s_expo3_30 ;
wire [8:0] s_expo3_31 ;
wire [8:0] s_expo3_3 ;
wire [5:0] s_shr1 ;
wire [26:0] s_qutnt_i ;
wire [8:0] s_expo3 ;
wire [30:22] s_output_o ;
wire [23:23] s_opa_i ;
wire s_shl1 ;
wire [26:0] s_fraco1_3 ;
wire [5:5] s_expo3_RNISDPK1_O6 ;
wire [8:0] s_expo1 ;
wire [6:6] s_expo1_3 ;
wire s_shl1_0_0 ;
wire [23:23] s_opb_i ;
wire [26:0] s_rmndr_i ;
wire [22:0] s_fraco2 ;
wire [3:3] v_count_1 ;
wire [3:1] v_count ;
wire [2:1] un2_s_lost ;
wire s_exp_10_i_1Q_Q31 ;
wire VCC ;
wire GND ;
wire s_exp_10_i_1Q_Q31_0 ;
wire s_exp_10_i_1Q_Q31_1 ;
wire s_exp_10_i_1Q_Q31_2 ;
wire s_exp_10_i_1Q_Q31_3 ;
wire s_exp_10_i_1Q_Q31_4 ;
wire s_exp_10_i_1Q_Q31_5 ;
wire s_exp_10_i_1Q_Q31_6 ;
wire s_exp_10_i_1Q_Q31_7 ;
wire s_exp_10_i_1Q_Q31_8 ;
wire un6_s_frac_rnd_1_axb_25 ;
wire s_exp_10b_axbxc8_RNIGLJC4 ;
wire v_shr_1_c4 ;
wire s_exp_10b_c5 ;
wire s_roundup ;
wire result_3_2_4 ;
wire result_3_3_4 ;
wire un18_s_roundup ;
wire un4_s_ine_o_1 ;
wire N_83 ;
wire N_84 ;
wire N_99 ;
wire N_100 ;
wire N_110 ;
wire N_111 ;
wire N_107 ;
wire N_82 ;
wire N_91 ;
wire N_98 ;
wire N_118 ;
wire N_109 ;
wire N_52 ;
wire N_44 ;
wire N_48 ;
wire N_102 ;
wire N_51 ;
wire N_89 ;
wire N_105 ;
wire N_116 ;
wire N_90 ;
wire N_106 ;
wire N_117 ;
wire un6_s_inf_result ;
wire un6_s_infa ;
wire N_33 ;
wire N_37 ;
wire N_41 ;
wire N_45 ;
wire N_60 ;
wire N_68 ;
wire N_123 ;
wire N_1424 ;
wire N_54 ;
wire un1_s_infa_0 ;
wire result_4_0_3 ;
wire N_1419 ;
wire N_1426 ;
wire N_1422 ;
wire N_1480 ;
wire N_1423 ;
wire N_1433 ;
wire N_108 ;
wire un1_s_shr1_1 ;
wire N_114 ;
wire un2_s_lost_0_c2 ;
wire N_271 ;
wire N_27 ;
wire s_exp_10b_axbxc7_lut6_2_RNIQA981 ;
wire un6_s_frac_rnd_0_axb_27 ;
wire un6_s_frac_rnd_0_axb_28 ;
wire un6_s_frac_rnd_0_axb_29 ;
wire un6_s_frac_rnd_0_axb_30 ;
wire un6_s_frac_rnd_0_axb_31 ;
wire un6_s_frac_rnd_0_axb_32 ;
wire un6_s_frac_rnd_0_axb_33 ;
wire un6_s_frac_rnd_1_cry_0_sf ;
wire un6_s_frac_rnd_1_axb_1 ;
wire un6_s_frac_rnd_1_axb_2 ;
wire un6_s_frac_rnd_1_axb_3 ;
wire un6_s_frac_rnd_1_axb_4 ;
wire un6_s_frac_rnd_1_axb_5 ;
wire un6_s_frac_rnd_1_axb_6 ;
wire un6_s_frac_rnd_1_axb_7 ;
wire un6_s_frac_rnd_1_axb_8 ;
wire un6_s_frac_rnd_1_axb_9 ;
wire un6_s_frac_rnd_1_axb_10 ;
wire un6_s_frac_rnd_1_axb_11 ;
wire un6_s_frac_rnd_1_axb_12 ;
wire un6_s_frac_rnd_1_axb_13 ;
wire un6_s_frac_rnd_1_axb_14 ;
wire un6_s_frac_rnd_1_axb_15 ;
wire un6_s_frac_rnd_1_axb_16 ;
wire un6_s_frac_rnd_1_axb_17 ;
wire un6_s_frac_rnd_1_axb_18 ;
wire un6_s_frac_rnd_1_axb_19 ;
wire un6_s_frac_rnd_1_axb_20 ;
wire un6_s_frac_rnd_1_axb_21 ;
wire un6_s_frac_rnd_1_axb_22 ;
wire un6_s_frac_rnd_1_axb_23 ;
wire un6_s_frac_rnd_1_axb_26 ;
wire un6_s_frac_rnd_1_axb_27 ;
wire un6_s_frac_rnd_1_axb_28 ;
wire un6_s_frac_rnd_1_axb_29 ;
wire un6_s_frac_rnd_1_axb_30 ;
wire un6_s_frac_rnd_1_axb_31 ;
wire un6_s_frac_rnd_1_axb_32 ;
wire un6_s_frac_rnd_1_axb_33 ;
wire N_1357_i ;
wire s_sign_i ;
wire un1_s_ine_o_0 ;
wire N_1479 ;
wire N_1488 ;
wire N_55 ;
wire N_50 ;
wire N_104 ;
wire N_93 ;
wire N_101 ;
wire N_95 ;
wire N_97 ;
wire N_103 ;
wire N_96 ;
wire N_94 ;
wire result_16 ;
wire result_4_2 ;
wire N_88 ;
wire N_115 ;
wire N_86 ;
wire N_113 ;
wire N_47 ;
wire N_85 ;
wire N_112 ;
wire m26_i ;
wire un4_s_lost_ac0_1 ;
wire un4_s_lost_ac0_2 ;
wire N_119 ;
wire N_114_0 ;
wire result_3_1_2 ;
wire N_1461_1 ;
wire un6_s_frac_rnd_1_axb_34 ;
wire un6_s_frac_rnd_0_axb_34 ;
wire N_1428 ;
wire N_1429 ;
wire N_1421 ;
wire N_1420 ;
wire N_1487 ;
wire N_26 ;
wire s_infb_0 ;
wire result_5_20 ;
wire result_5_1_0 ;
wire result_5_0 ;
wire result_3_3 ;
wire result_3_2 ;
wire result_3_0 ;
wire result_1_21_1 ;
wire result_1_21_0 ;
wire result_3 ;
wire N_28 ;
wire N_31 ;
wire N_46 ;
wire N_43 ;
wire N_42 ;
wire N_40 ;
wire N_39 ;
wire N_38 ;
wire N_36 ;
wire N_35 ;
wire N_34 ;
wire N_32 ;
wire N_30 ;
wire N_29 ;
wire N_49 ;
wire m26_i_1 ;
wire N_1416_2 ;
wire result_5_28 ;
wire m73_i ;
wire N_1437 ;
wire N_1431 ;
wire N_92 ;
wire un16_s_roundup ;
wire N_148 ;
wire un7_s_nan_in ;
wire N_1483 ;
wire N_1455 ;
wire un4_s_lost_c3 ;
wire un4_s_lost_c4 ;
wire un4_s_lost_c5 ;
wire un6_s_frac_rnd_1_cry_33 ;
wire un6_s_frac_rnd_1_cry_32 ;
wire un6_s_frac_rnd_1_cry_31 ;
wire un6_s_frac_rnd_1_cry_30 ;
wire un6_s_frac_rnd_1_cry_29 ;
wire un6_s_frac_rnd_1_cry_28 ;
wire un6_s_frac_rnd_1_cry_27 ;
wire un6_s_frac_rnd_1_cry_26 ;
wire un6_s_frac_rnd_1_cry_25 ;
wire un6_s_frac_rnd_1_cry_24 ;
wire un6_s_frac_rnd_1_cry_22 ;
wire un6_s_frac_rnd_1_cry_21 ;
wire un6_s_frac_rnd_1_cry_20 ;
wire un6_s_frac_rnd_1_cry_19 ;
wire un6_s_frac_rnd_1_cry_18 ;
wire un6_s_frac_rnd_1_cry_17 ;
wire un6_s_frac_rnd_1_cry_16 ;
wire un6_s_frac_rnd_1_cry_15 ;
wire un6_s_frac_rnd_1_cry_14 ;
wire un6_s_frac_rnd_1_cry_13 ;
wire un6_s_frac_rnd_1_cry_12 ;
wire un6_s_frac_rnd_1_cry_11 ;
wire un6_s_frac_rnd_1_cry_10 ;
wire un6_s_frac_rnd_1_cry_9 ;
wire un6_s_frac_rnd_1_cry_8 ;
wire un6_s_frac_rnd_1_cry_7 ;
wire un6_s_frac_rnd_1_cry_6 ;
wire un6_s_frac_rnd_1_cry_5 ;
wire un6_s_frac_rnd_1_cry_4 ;
wire un6_s_frac_rnd_1_cry_3 ;
wire un6_s_frac_rnd_1_cry_2 ;
wire un6_s_frac_rnd_1_cry_1 ;
wire un6_s_frac_rnd_1_cry_0 ;
wire un6_s_frac_rnd_0_cry_33 ;
wire un6_s_frac_rnd_0_cry_32 ;
wire un6_s_frac_rnd_0_cry_31 ;
wire un6_s_frac_rnd_0_cry_30 ;
wire un6_s_frac_rnd_0_cry_29 ;
wire un6_s_frac_rnd_0_cry_28 ;
wire un6_s_frac_rnd_0_cry_27 ;
wire un6_s_frac_rnd_0_cry_26 ;
// instances
  SRLC32E desc2213(.Q(s_exp_10_i_8_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[1:1]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2214(.Q(s_exp_10_i_7_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_0),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_axb_0_i),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2215(.Q(s_exp_10_i_6_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_1),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[9:9]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2216(.Q(s_exp_10_i_5_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_2),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[8:8]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2217(.Q(s_exp_10_i_4_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_3),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[7:7]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2218(.Q(s_exp_10_i_3_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_4),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[6:6]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2219(.Q(s_exp_10_i_2_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_5),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[5:5]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2220(.Q(s_exp_10_i_1_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_6),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[4:4]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2221(.Q(s_exp_10_i_0_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_7),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[3:3]),.CLK(clk_i),.CE(VCC));
  SRLC32E desc2222(.Q(s_exp_10_i_tmp_d_array_0),.Q31(s_exp_10_i_1Q_Q31_8),.A({GND,GND,GND,GND,VCC}),.D(un11_s_exp_10_o_0[2:2]),.CLK(clk_i),.CE(VCC));
  LUT1 un6_s_frac_rnd_1_axb_25_cZ(.I0(GND),.O(un6_s_frac_rnd_1_axb_25));
defparam un6_s_frac_rnd_1_axb_25_cZ.INIT=2'h3;
  LUT6 desc2223(.I0(s_exp_10b_axbxc7_lut6_2_RNIQA981),.I1(s_exp_10_i[0:0]),.I2(s_exp_10b[8:8]),.I3(s_exp_10b[9:9]),.I4(s_expo1_3[6:6]),.I5(s_qutnt_i[26:26]),.O(s_shl1_0_0));
defparam desc2223.INIT=64'h00000000080F0007;
  LUT2 un6_s_frac_rnd_0_cry_26_RNO(.I0(s_expo1[0:0]),.I1(s_fraco1[26:26]),.O(s_expo3_30[0:0]));
defparam un6_s_frac_rnd_0_cry_26_RNO.INIT=4'h9;
  LUT2 desc2224(.I0(s_expo1[1:1]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_27));
defparam desc2224.INIT=4'h9;
  LUT2 desc2225(.I0(s_expo1[2:2]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_28));
defparam desc2225.INIT=4'h9;
  LUT2 desc2226(.I0(s_expo1[3:3]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_29));
defparam desc2226.INIT=4'h9;
  LUT2 desc2227(.I0(s_expo1[4:4]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_30));
defparam desc2227.INIT=4'h9;
  LUT2 desc2228(.I0(s_expo1[5:5]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_31));
defparam desc2228.INIT=4'h9;
  LUT2 desc2229(.I0(s_expo1[6:6]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_32));
defparam desc2229.INIT=4'h9;
  LUT2 desc2230(.I0(s_expo1[7:7]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_33));
defparam desc2230.INIT=4'h9;
  LUT1 un6_s_frac_rnd_1_cry_0_RNO(.I0(s_fraco1[3:3]),.O(un6_s_frac_rnd_1_cry_0_sf));
defparam un6_s_frac_rnd_1_cry_0_RNO.INIT=2'h1;
  LUT1 desc2231(.I0(s_fraco1[4:4]),.O(un6_s_frac_rnd_1_axb_1));
defparam desc2231.INIT=2'h2;
  LUT1 desc2232(.I0(s_fraco1[5:5]),.O(un6_s_frac_rnd_1_axb_2));
defparam desc2232.INIT=2'h2;
  LUT1 desc2233(.I0(s_fraco1[6:6]),.O(un6_s_frac_rnd_1_axb_3));
defparam desc2233.INIT=2'h2;
  LUT1 desc2234(.I0(s_fraco1[7:7]),.O(un6_s_frac_rnd_1_axb_4));
defparam desc2234.INIT=2'h2;
  LUT1 desc2235(.I0(s_fraco1[8:8]),.O(un6_s_frac_rnd_1_axb_5));
defparam desc2235.INIT=2'h2;
  LUT1 desc2236(.I0(s_fraco1[9:9]),.O(un6_s_frac_rnd_1_axb_6));
defparam desc2236.INIT=2'h2;
  LUT1 desc2237(.I0(s_fraco1[10:10]),.O(un6_s_frac_rnd_1_axb_7));
defparam desc2237.INIT=2'h2;
  LUT1 desc2238(.I0(s_fraco1[11:11]),.O(un6_s_frac_rnd_1_axb_8));
defparam desc2238.INIT=2'h2;
  LUT1 desc2239(.I0(s_fraco1[12:12]),.O(un6_s_frac_rnd_1_axb_9));
defparam desc2239.INIT=2'h2;
  LUT1 desc2240(.I0(s_fraco1[13:13]),.O(un6_s_frac_rnd_1_axb_10));
defparam desc2240.INIT=2'h2;
  LUT1 desc2241(.I0(s_fraco1[14:14]),.O(un6_s_frac_rnd_1_axb_11));
defparam desc2241.INIT=2'h2;
  LUT1 desc2242(.I0(s_fraco1[15:15]),.O(un6_s_frac_rnd_1_axb_12));
defparam desc2242.INIT=2'h2;
  LUT1 desc2243(.I0(s_fraco1[16:16]),.O(un6_s_frac_rnd_1_axb_13));
defparam desc2243.INIT=2'h2;
  LUT1 desc2244(.I0(s_fraco1[17:17]),.O(un6_s_frac_rnd_1_axb_14));
defparam desc2244.INIT=2'h2;
  LUT1 desc2245(.I0(s_fraco1[18:18]),.O(un6_s_frac_rnd_1_axb_15));
defparam desc2245.INIT=2'h2;
  LUT1 desc2246(.I0(s_fraco1[19:19]),.O(un6_s_frac_rnd_1_axb_16));
defparam desc2246.INIT=2'h2;
  LUT1 desc2247(.I0(s_fraco1[20:20]),.O(un6_s_frac_rnd_1_axb_17));
defparam desc2247.INIT=2'h2;
  LUT1 desc2248(.I0(s_fraco1[21:21]),.O(un6_s_frac_rnd_1_axb_18));
defparam desc2248.INIT=2'h2;
  LUT1 desc2249(.I0(s_fraco1[22:22]),.O(un6_s_frac_rnd_1_axb_19));
defparam desc2249.INIT=2'h2;
  LUT1 desc2250(.I0(s_fraco1[23:23]),.O(un6_s_frac_rnd_1_axb_20));
defparam desc2250.INIT=2'h2;
  LUT1 desc2251(.I0(s_fraco1[24:24]),.O(un6_s_frac_rnd_1_axb_21));
defparam desc2251.INIT=2'h2;
  LUT1 desc2252(.I0(s_fraco1[25:25]),.O(un6_s_frac_rnd_1_axb_22));
defparam desc2252.INIT=2'h2;
  LUT1 un6_s_frac_rnd_1_cry_23_RNO(.I0(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_23));
defparam un6_s_frac_rnd_1_cry_23_RNO.INIT=2'h2;
  LUT2 desc2253(.I0(s_expo1[0:0]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_26));
defparam desc2253.INIT=4'h9;
  LUT2 desc2254(.I0(s_expo1[1:1]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_27));
defparam desc2254.INIT=4'h9;
  LUT2 desc2255(.I0(s_expo1[2:2]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_28));
defparam desc2255.INIT=4'h9;
  LUT2 desc2256(.I0(s_expo1[3:3]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_29));
defparam desc2256.INIT=4'h9;
  LUT2 desc2257(.I0(s_expo1[4:4]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_30));
defparam desc2257.INIT=4'h9;
  LUT2 desc2258(.I0(s_expo1[5:5]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_31));
defparam desc2258.INIT=4'h9;
  LUT2 desc2259(.I0(s_expo1[6:6]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_32));
defparam desc2259.INIT=4'h9;
  LUT2 desc2260(.I0(s_expo1[7:7]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_33));
defparam desc2260.INIT=4'h9;
  FD desc2261(.Q(s_opb_i_4),.D(s_opb_i_0[27:27]),.C(clk_i));
  FD desc2262(.Q(s_opb_i_5),.D(s_opb_i_0[28:28]),.C(clk_i));
  FD desc2263(.Q(s_opb_i_6),.D(s_opb_i_0[29:29]),.C(clk_i));
  FD desc2264(.Q(s_opb_i_7),.D(s_opb_i_0[30:30]),.C(clk_i));
  FD desc2265(.Q(s_opb_i[23:23]),.D(s_opb_i_0[23:23]),.C(clk_i));
  FD desc2266(.Q(s_opb_i_1),.D(s_opb_i_0[24:24]),.C(clk_i));
  FD desc2267(.Q(s_opb_i_2),.D(s_opb_i_0[25:25]),.C(clk_i));
  FD desc2268(.Q(s_opb_i_3),.D(s_opb_i_0[26:26]),.C(clk_i));
  FD desc2269(.Q(s_opa_i_5),.D(s_opa_i_0[28:28]),.C(clk_i));
  FD desc2270(.Q(s_opa_i_6),.D(s_opa_i_0[29:29]),.C(clk_i));
  FD desc2271(.Q(s_opa_i_7),.D(s_opa_i_0[30:30]),.C(clk_i));
  FD desc2272(.Q(s_opa_i[23:23]),.D(s_opa_i_0[23:23]),.C(clk_i));
  FD desc2273(.Q(s_opa_i_1),.D(s_opa_i_0[24:24]),.C(clk_i));
  FD desc2274(.Q(s_opa_i_2),.D(s_opa_i_0[25:25]),.C(clk_i));
  FD desc2275(.Q(s_opa_i_3),.D(s_opa_i_0[26:26]),.C(clk_i));
  FD desc2276(.Q(s_opa_i_4),.D(s_opa_i_0[27:27]),.C(clk_i));
  FD desc2277(.Q(s_rmndr_i[25:25]),.D(serial_div_rmndr[25:25]),.C(clk_i));
  FD desc2278(.Q(s_rmndr_i[26:26]),.D(serial_div_rmndr[26:26]),.C(clk_i));
  FD desc2279(.Q(s_rmndr_i[10:10]),.D(serial_div_rmndr[10:10]),.C(clk_i));
  FD desc2280(.Q(s_rmndr_i[11:11]),.D(serial_div_rmndr[11:11]),.C(clk_i));
  FD desc2281(.Q(s_rmndr_i[12:12]),.D(serial_div_rmndr[12:12]),.C(clk_i));
  FD desc2282(.Q(s_rmndr_i[13:13]),.D(serial_div_rmndr[13:13]),.C(clk_i));
  FD desc2283(.Q(s_rmndr_i[14:14]),.D(serial_div_rmndr[14:14]),.C(clk_i));
  FD desc2284(.Q(s_rmndr_i[15:15]),.D(serial_div_rmndr[15:15]),.C(clk_i));
  FD desc2285(.Q(s_rmndr_i[16:16]),.D(serial_div_rmndr[16:16]),.C(clk_i));
  FD desc2286(.Q(s_rmndr_i[17:17]),.D(serial_div_rmndr[17:17]),.C(clk_i));
  FD desc2287(.Q(s_rmndr_i[18:18]),.D(serial_div_rmndr[18:18]),.C(clk_i));
  FD desc2288(.Q(s_rmndr_i[19:19]),.D(serial_div_rmndr[19:19]),.C(clk_i));
  FD desc2289(.Q(s_rmndr_i[20:20]),.D(serial_div_rmndr[20:20]),.C(clk_i));
  FD desc2290(.Q(s_rmndr_i[21:21]),.D(serial_div_rmndr[21:21]),.C(clk_i));
  FD desc2291(.Q(s_rmndr_i[22:22]),.D(serial_div_rmndr[22:22]),.C(clk_i));
  FD desc2292(.Q(s_rmndr_i[23:23]),.D(serial_div_rmndr[23:23]),.C(clk_i));
  FD desc2293(.Q(s_rmndr_i[24:24]),.D(serial_div_rmndr[24:24]),.C(clk_i));
  FD desc2294(.Q(s_qutnt_i[22:22]),.D(serial_div_qutnt[22:22]),.C(clk_i));
  FD desc2295(.Q(s_qutnt_i[23:23]),.D(serial_div_qutnt[23:23]),.C(clk_i));
  FD desc2296(.Q(s_qutnt_i[24:24]),.D(serial_div_qutnt[24:24]),.C(clk_i));
  FD desc2297(.Q(s_qutnt_i[25:25]),.D(serial_div_qutnt[25:25]),.C(clk_i));
  FD desc2298(.Q(s_qutnt_i[26:26]),.D(serial_div_qutnt[26:26]),.C(clk_i));
  FD desc2299(.Q(s_rmndr_i[0:0]),.D(serial_div_rmndr[0:0]),.C(clk_i));
  FD desc2300(.Q(s_rmndr_i[1:1]),.D(serial_div_rmndr[1:1]),.C(clk_i));
  FD desc2301(.Q(s_rmndr_i[2:2]),.D(serial_div_rmndr[2:2]),.C(clk_i));
  FD desc2302(.Q(s_rmndr_i[3:3]),.D(serial_div_rmndr[3:3]),.C(clk_i));
  FD desc2303(.Q(s_rmndr_i[4:4]),.D(serial_div_rmndr[4:4]),.C(clk_i));
  FD desc2304(.Q(s_rmndr_i[5:5]),.D(serial_div_rmndr[5:5]),.C(clk_i));
  FD desc2305(.Q(s_rmndr_i[6:6]),.D(serial_div_rmndr[6:6]),.C(clk_i));
  FD desc2306(.Q(s_rmndr_i[7:7]),.D(serial_div_rmndr[7:7]),.C(clk_i));
  FD desc2307(.Q(s_rmndr_i[8:8]),.D(serial_div_rmndr[8:8]),.C(clk_i));
  FD desc2308(.Q(s_rmndr_i[9:9]),.D(serial_div_rmndr[9:9]),.C(clk_i));
  FD desc2309(.Q(s_qutnt_i[7:7]),.D(serial_div_qutnt[7:7]),.C(clk_i));
  FD desc2310(.Q(s_qutnt_i[8:8]),.D(serial_div_qutnt[8:8]),.C(clk_i));
  FD desc2311(.Q(s_qutnt_i[9:9]),.D(serial_div_qutnt[9:9]),.C(clk_i));
  FD desc2312(.Q(s_qutnt_i[10:10]),.D(serial_div_qutnt[10:10]),.C(clk_i));
  FD desc2313(.Q(s_qutnt_i[11:11]),.D(serial_div_qutnt[11:11]),.C(clk_i));
  FD desc2314(.Q(s_qutnt_i[12:12]),.D(serial_div_qutnt[12:12]),.C(clk_i));
  FD desc2315(.Q(s_qutnt_i[13:13]),.D(serial_div_qutnt[13:13]),.C(clk_i));
  FD desc2316(.Q(s_qutnt_i[14:14]),.D(serial_div_qutnt[14:14]),.C(clk_i));
  FD desc2317(.Q(s_qutnt_i[15:15]),.D(serial_div_qutnt[15:15]),.C(clk_i));
  FD desc2318(.Q(s_qutnt_i[16:16]),.D(serial_div_qutnt[16:16]),.C(clk_i));
  FD desc2319(.Q(s_qutnt_i[17:17]),.D(serial_div_qutnt[17:17]),.C(clk_i));
  FD desc2320(.Q(s_qutnt_i[18:18]),.D(serial_div_qutnt[18:18]),.C(clk_i));
  FD desc2321(.Q(s_qutnt_i[19:19]),.D(serial_div_qutnt[19:19]),.C(clk_i));
  FD desc2322(.Q(s_qutnt_i[20:20]),.D(serial_div_qutnt[20:20]),.C(clk_i));
  FD desc2323(.Q(s_qutnt_i[21:21]),.D(serial_div_qutnt[21:21]),.C(clk_i));
  FD desc2324(.Q(s_qutnt_i[0:0]),.D(serial_div_qutnt[0:0]),.C(clk_i));
  FD desc2325(.Q(s_qutnt_i[1:1]),.D(serial_div_qutnt[1:1]),.C(clk_i));
  FD desc2326(.Q(s_qutnt_i[2:2]),.D(serial_div_qutnt[2:2]),.C(clk_i));
  FD desc2327(.Q(s_qutnt_i[3:3]),.D(serial_div_qutnt[3:3]),.C(clk_i));
  FD desc2328(.Q(s_qutnt_i[4:4]),.D(serial_div_qutnt[4:4]),.C(clk_i));
  FD desc2329(.Q(s_qutnt_i[5:5]),.D(serial_div_qutnt[5:5]),.C(clk_i));
  FD desc2330(.Q(s_qutnt_i[6:6]),.D(serial_div_qutnt[6:6]),.C(clk_i));
  FD desc2331(.Q(s_fraco2[12:12]),.D(s_frac_rnd[12:12]),.C(clk_i));
  FD desc2332(.Q(s_fraco2[13:13]),.D(s_frac_rnd[13:13]),.C(clk_i));
  FD desc2333(.Q(s_fraco2[14:14]),.D(s_frac_rnd[14:14]),.C(clk_i));
  FD desc2334(.Q(s_fraco2[15:15]),.D(s_frac_rnd[15:15]),.C(clk_i));
  FD desc2335(.Q(s_fraco2[16:16]),.D(s_frac_rnd[16:16]),.C(clk_i));
  FD desc2336(.Q(s_fraco2[17:17]),.D(s_frac_rnd[17:17]),.C(clk_i));
  FD desc2337(.Q(s_fraco2[18:18]),.D(s_frac_rnd[18:18]),.C(clk_i));
  FD desc2338(.Q(s_fraco2[19:19]),.D(s_frac_rnd[19:19]),.C(clk_i));
  FD desc2339(.Q(s_fraco2[20:20]),.D(s_frac_rnd[20:20]),.C(clk_i));
  FD desc2340(.Q(s_fraco2[21:21]),.D(s_frac_rnd[21:21]),.C(clk_i));
  FD desc2341(.Q(s_fraco2[22:22]),.D(s_frac_rnd[22:22]),.C(clk_i));
  FD desc2342(.Q(s_rmode_i[0:0]),.D(s_rmode_i_0[0:0]),.C(clk_i));
  FD desc2343(.Q(s_rmode_i[1:1]),.D(s_rmode_i_0[1:1]),.C(clk_i));
  FD desc2344(.Q(s_fraco2[0:0]),.D(s_frac_rnd[0:0]),.C(clk_i));
  FD desc2345(.Q(s_fraco2[1:1]),.D(s_frac_rnd[1:1]),.C(clk_i));
  FD desc2346(.Q(s_fraco2[2:2]),.D(s_frac_rnd[2:2]),.C(clk_i));
  FD desc2347(.Q(s_fraco2[3:3]),.D(s_frac_rnd[3:3]),.C(clk_i));
  FD desc2348(.Q(s_fraco2[4:4]),.D(s_frac_rnd[4:4]),.C(clk_i));
  FD desc2349(.Q(s_fraco2[5:5]),.D(s_frac_rnd[5:5]),.C(clk_i));
  FD desc2350(.Q(s_fraco2[6:6]),.D(s_frac_rnd[6:6]),.C(clk_i));
  FD desc2351(.Q(s_fraco2[7:7]),.D(s_frac_rnd[7:7]),.C(clk_i));
  FD desc2352(.Q(s_fraco2[8:8]),.D(s_frac_rnd[8:8]),.C(clk_i));
  FD desc2353(.Q(s_fraco2[9:9]),.D(s_frac_rnd[9:9]),.C(clk_i));
  FD desc2354(.Q(s_fraco2[10:10]),.D(s_frac_rnd[10:10]),.C(clk_i));
  FD desc2355(.Q(s_fraco2[11:11]),.D(s_frac_rnd[11:11]),.C(clk_i));
  FD desc2356(.Q(s_fraco1[26:26]),.D(s_fraco1_3[26:26]),.C(clk_i));
  FD desc2357(.Q(s_expo1[0:0]),.D(N_1357_i),.C(clk_i));
  FD desc2358(.Q(s_expo1[6:6]),.D(s_expo1_3[6:6]),.C(clk_i));
  FD desc2359(.Q(s_fraco1[11:11]),.D(s_fraco1_3[11:11]),.C(clk_i));
  FD desc2360(.Q(s_fraco1[12:12]),.D(s_fraco1_3[12:12]),.C(clk_i));
  FD desc2361(.Q(s_fraco1[13:13]),.D(s_fraco1_3[13:13]),.C(clk_i));
  FD desc2362(.Q(s_fraco1[14:14]),.D(s_fraco1_3[14:14]),.C(clk_i));
  FD desc2363(.Q(s_fraco1[15:15]),.D(s_fraco1_3[15:15]),.C(clk_i));
  FD desc2364(.Q(s_fraco1[16:16]),.D(s_fraco1_3[16:16]),.C(clk_i));
  FD desc2365(.Q(s_fraco1[17:17]),.D(s_fraco1_3[17:17]),.C(clk_i));
  FD desc2366(.Q(s_fraco1[18:18]),.D(s_fraco1_3[18:18]),.C(clk_i));
  FD desc2367(.Q(s_fraco1[19:19]),.D(s_fraco1_3[19:19]),.C(clk_i));
  FD desc2368(.Q(s_fraco1[20:20]),.D(s_fraco1_3[20:20]),.C(clk_i));
  FD desc2369(.Q(s_fraco1[21:21]),.D(s_fraco1_3[21:21]),.C(clk_i));
  FD desc2370(.Q(s_fraco1[22:22]),.D(s_fraco1_3[22:22]),.C(clk_i));
  FD desc2371(.Q(s_fraco1[23:23]),.D(s_fraco1_3[23:23]),.C(clk_i));
  FD desc2372(.Q(s_fraco1[24:24]),.D(s_fraco1_3[24:24]),.C(clk_i));
  FD desc2373(.Q(s_fraco1[25:25]),.D(s_fraco1_3[25:25]),.C(clk_i));
  FD desc2374(.Q(s_fraco1[0:0]),.D(s_fraco1_3[0:0]),.C(clk_i));
  FD desc2375(.Q(s_fraco1[1:1]),.D(s_fraco1_3[1:1]),.C(clk_i));
  FD desc2376(.Q(s_fraco1[2:2]),.D(s_fraco1_3[2:2]),.C(clk_i));
  FD desc2377(.Q(s_fraco1[3:3]),.D(s_fraco1_3[3:3]),.C(clk_i));
  FD desc2378(.Q(s_fraco1[4:4]),.D(s_fraco1_3[4:4]),.C(clk_i));
  FD desc2379(.Q(s_fraco1[5:5]),.D(s_fraco1_3[5:5]),.C(clk_i));
  FD desc2380(.Q(s_fraco1[6:6]),.D(s_fraco1_3[6:6]),.C(clk_i));
  FD desc2381(.Q(s_fraco1[7:7]),.D(s_fraco1_3[7:7]),.C(clk_i));
  FD desc2382(.Q(s_fraco1[8:8]),.D(s_fraco1_3[8:8]),.C(clk_i));
  FD desc2383(.Q(s_fraco1[9:9]),.D(s_fraco1_3[9:9]),.C(clk_i));
  FD desc2384(.Q(s_fraco1[10:10]),.D(s_fraco1_3[10:10]),.C(clk_i));
  FD desc2385(.Q(s_expo3[2:2]),.D(s_expo3_3[2:2]),.C(clk_i));
  FD desc2386(.Q(s_expo3[3:3]),.D(s_expo3_3[3:3]),.C(clk_i));
  FD desc2387(.Q(s_expo3[4:4]),.D(s_expo3_3[4:4]),.C(clk_i));
  FD desc2388(.Q(s_expo3[5:5]),.D(s_expo3_3[5:5]),.C(clk_i));
  FD desc2389(.Q(s_expo3[6:6]),.D(s_expo3_3[6:6]),.C(clk_i));
  FD desc2390(.Q(s_expo3[7:7]),.D(s_expo3_3[7:7]),.C(clk_i));
  FD desc2391(.Q(s_expo3[8:8]),.D(s_expo3_3[8:8]),.C(clk_i));
  FD desc2392(.Q(s_expo3[0:0]),.D(s_expo3_3[0:0]),.C(clk_i));
  FD desc2393(.Q(s_expo3[1:1]),.D(s_expo3_3[1:1]),.C(clk_i));
  FD s_sign_i_Z(.Q(s_sign_i),.D(N_1942_i),.C(clk_i));
  FD ine_o_Z(.Q(post_norm_div_ine),.D(un1_s_ine_o_0),.C(clk_i));
  FDR desc2394(.Q(post_norm_div_output[0:0]),.D(s_fraco2[0:0]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2395(.Q(post_norm_div_output[1:1]),.D(s_fraco2[1:1]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2396(.Q(post_norm_div_output[2:2]),.D(s_fraco2[2:2]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2397(.Q(post_norm_div_output[3:3]),.D(s_fraco2[3:3]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2398(.Q(post_norm_div_output[4:4]),.D(s_fraco2[4:4]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2399(.Q(post_norm_div_output[5:5]),.D(s_fraco2[5:5]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2400(.Q(post_norm_div_output[6:6]),.D(s_fraco2[6:6]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2401(.Q(post_norm_div_output[7:7]),.D(s_fraco2[7:7]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2402(.Q(post_norm_div_output[8:8]),.D(s_fraco2[8:8]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2403(.Q(post_norm_div_output[9:9]),.D(s_fraco2[9:9]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2404(.Q(post_norm_div_output[10:10]),.D(s_fraco2[10:10]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2405(.Q(post_norm_div_output[11:11]),.D(s_fraco2[11:11]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2406(.Q(post_norm_div_output[12:12]),.D(s_fraco2[12:12]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2407(.Q(post_norm_div_output[13:13]),.D(s_fraco2[13:13]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2408(.Q(post_norm_div_output[14:14]),.D(s_fraco2[14:14]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2409(.Q(post_norm_div_output[15:15]),.D(s_fraco2[15:15]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2410(.Q(post_norm_div_output[16:16]),.D(s_fraco2[16:16]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2411(.Q(post_norm_div_output[17:17]),.D(s_fraco2[17:17]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2412(.Q(post_norm_div_output[18:18]),.D(s_fraco2[18:18]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2413(.Q(post_norm_div_output[19:19]),.D(s_fraco2[19:19]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2414(.Q(post_norm_div_output[20:20]),.D(s_fraco2[20:20]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2415(.Q(post_norm_div_output[21:21]),.D(s_fraco2[21:21]),.C(clk_i),.R(s_expo3_RNISDPK1_O6[5:5]));
  FDR desc2416(.Q(s_expo1[1:1]),.D(s_exp_10b[1:1]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2417(.Q(s_expo1[2:2]),.D(s_exp_10b[2:2]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2418(.Q(s_expo1[3:3]),.D(s_exp_10b[3:3]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2419(.Q(s_expo1[4:4]),.D(s_exp_10b[4:4]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2420(.Q(s_expo1[5:5]),.D(s_exp_10b[5:5]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2421(.Q(s_expo1[7:7]),.D(s_exp_10b[7:7]),.C(clk_i),.R(s_exp_10b[9:9]));
  FDR desc2422(.Q(s_expo1[8:8]),.D(s_exp_10b[8:8]),.C(clk_i),.R(s_exp_10b[9:9]));
  FD desc2423(.Q(s_exp_10_i[2:2]),.D(s_exp_10_i_tmp_d_array_0),.C(clk_i));
  FD desc2424(.Q(s_exp_10_i[3:3]),.D(s_exp_10_i_0_tmp_d_array_0),.C(clk_i));
  FD desc2425(.Q(s_exp_10_i[4:4]),.D(s_exp_10_i_1_tmp_d_array_0),.C(clk_i));
  FD desc2426(.Q(s_exp_10_i[5:5]),.D(s_exp_10_i_2_tmp_d_array_0),.C(clk_i));
  FD desc2427(.Q(s_exp_10_i[6:6]),.D(s_exp_10_i_3_tmp_d_array_0),.C(clk_i));
  FD desc2428(.Q(s_exp_10_i[7:7]),.D(s_exp_10_i_4_tmp_d_array_0),.C(clk_i));
  FD desc2429(.Q(s_exp_10_i[8:8]),.D(s_exp_10_i_5_tmp_d_array_0),.C(clk_i));
  FD desc2430(.Q(s_exp_10_i[9:9]),.D(s_exp_10_i_6_tmp_d_array_0),.C(clk_i));
  FD desc2431(.Q(s_exp_10_i[0:0]),.D(s_exp_10_i_7_tmp_d_array_0),.C(clk_i));
  FD desc2432(.Q(s_exp_10_i[1:1]),.D(s_exp_10_i_8_tmp_d_array_0),.C(clk_i));
  LUT5_L desc2433(.I0(s_expo3[4:4]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[27:27]));
defparam desc2433.INIT=32'hFFFFFEFC;
  LUT5_L desc2434(.I0(s_expo3[6:6]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[29:29]));
defparam desc2434.INIT=32'hFFFFFEFC;
  LUT5_L desc2435(.I0(s_expo3[7:7]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[30:30]));
defparam desc2435.INIT=32'hFFFFFEFC;
  LUT5_L desc2436(.I0(s_expo3[3:3]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[26:26]));
defparam desc2436.INIT=32'hFFFFFEFC;
  LUT5_L desc2437(.I0(s_expo3[2:2]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[25:25]));
defparam desc2437.INIT=32'hFFFFFEFC;
  LUT5_L desc2438(.I0(s_fraco2[22:22]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[22:22]));
defparam desc2438.INIT=32'h00000200;
  LUT5_L desc2439(.I0(s_expo3[1:1]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.LO(s_output_o[24:24]));
defparam desc2439.INIT=32'hFFFFFEFC;
  LUT6 desc2440(.I0(s_qutnt_i[0:0]),.I1(s_qutnt_i[1:1]),.I2(s_qutnt_i[2:2]),.I3(s_qutnt_i[3:3]),.I4(N_1422),.I5(N_1479),.O(N_1488));
defparam desc2440.INIT=64'h0000000100000000;
  LUT6_L desc2441(.I0(s_qutnt_i[8:8]),.I1(s_qutnt_i[9:9]),.I2(N_55),.I3(N_1433),.I4(N_1480),.I5(N_1426),.LO(v_count_1[3:3]));
defparam desc2441.INIT=64'h00FF000000FE0000;
  LUT6 desc2442(.I0(s_qutnt_i[26:26]),.I1(s_shr1[0:0]),.I2(s_shr1[1:1]),.I3(s_shr1[3:3]),.I4(s_shr1[2:2]),.I5(N_50),.O(N_104));
defparam desc2442.INIT=64'h000200FF00020000;
  LUT6_L desc2443(.I0(s_qutnt_i[10:10]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_93),.LO(s_fraco1_3[11:11]));
defparam desc2443.INIT=64'h888B000F88880000;
  LUT6_L desc2444(.I0(s_qutnt_i[18:18]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_101),.LO(s_fraco1_3[19:19]));
defparam desc2444.INIT=64'h888B000F88880000;
  LUT6_L desc2445(.I0(s_qutnt_i[12:12]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_95),.LO(s_fraco1_3[13:13]));
defparam desc2445.INIT=64'h888B000F88880000;
  LUT6_L desc2446(.I0(s_qutnt_i[14:14]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_97),.LO(s_fraco1_3[15:15]));
defparam desc2446.INIT=64'h888B000F88880000;
  LUT6_L desc2447(.I0(s_qutnt_i[22:22]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_105),.LO(s_fraco1_3[23:23]));
defparam desc2447.INIT=64'h888B000F88880000;
  LUT6_L desc2448(.I0(s_qutnt_i[15:15]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_98),.LO(s_fraco1_3[16:16]));
defparam desc2448.INIT=64'h888B000F88880000;
  LUT6_L desc2449(.I0(s_qutnt_i[21:21]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_104),.LO(s_fraco1_3[22:22]));
defparam desc2449.INIT=64'h888B000F88880000;
  LUT6_L desc2450(.I0(s_qutnt_i[23:23]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_106),.LO(s_fraco1_3[24:24]));
defparam desc2450.INIT=64'h888B000F88880000;
  LUT6_L desc2451(.I0(s_qutnt_i[17:17]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_100),.LO(s_fraco1_3[18:18]));
defparam desc2451.INIT=64'h888B000F88880000;
  LUT6_L desc2452(.I0(s_qutnt_i[20:20]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_103),.LO(s_fraco1_3[21:21]));
defparam desc2452.INIT=64'h888B000F88880000;
  LUT6_L desc2453(.I0(s_qutnt_i[24:24]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(N_107),.I5(un1_s_shr1_1),.LO(s_fraco1_3[25:25]));
defparam desc2453.INIT=64'h888B8888000F0000;
  LUT6_L desc2454(.I0(s_qutnt_i[19:19]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_102),.LO(s_fraco1_3[20:20]));
defparam desc2454.INIT=64'h888B000F88880000;
  LUT6_L desc2455(.I0(s_qutnt_i[16:16]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_99),.LO(s_fraco1_3[17:17]));
defparam desc2455.INIT=64'h888B000F88880000;
  LUT6_L desc2456(.I0(s_qutnt_i[13:13]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_96),.LO(s_fraco1_3[14:14]));
defparam desc2456.INIT=64'h888B000F88880000;
  LUT6_L desc2457(.I0(s_qutnt_i[11:11]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(s_shr1[4:4]),.I4(un1_s_shr1_1),.I5(N_94),.LO(s_fraco1_3[12:12]));
defparam desc2457.INIT=64'h888B000F88880000;
  LUT6 desc2458(.I0(s_fracta_i[20:20]),.I1(s_fracta_i[21:21]),.I2(s_opa_i_5),.I3(s_opa_i_6),.I4(s_opa_i_7),.I5(result_16),.O(result_4_2));
defparam desc2458.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2459(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_54),.I4(N_50),.I5(N_88),.O(N_115));
defparam desc2459.INIT=64'h7757755522022000;
  LUT6 desc2460(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_52),.I4(N_48),.I5(N_86),.O(N_113));
defparam desc2460.INIT=64'h7757755522022000;
  LUT6 desc2461(.I0(s_qutnt_i[25:25]),.I1(s_qutnt_i[26:26]),.I2(s_shr1[0:0]),.I3(s_shr1[1:1]),.I4(s_shr1[3:3]),.I5(s_shr1[2:2]),.O(N_107));
defparam desc2461.INIT=64'h00000000000000CA;
  LUT6 un1_s_shr1_1_cZ(.I0(s_shr1[5:5]),.I1(s_shr1[4:4]),.I2(s_shr1[0:0]),.I3(s_shr1[1:1]),.I4(s_shr1[3:3]),.I5(s_shr1[2:2]),.O(un1_s_shr1_1));
defparam un1_s_shr1_1_cZ.INIT=64'h0000000000000001;
  LUT6 desc2462(.I0(s_qutnt_i[23:23]),.I1(s_qutnt_i[24:24]),.I2(s_qutnt_i[25:25]),.I3(s_qutnt_i[26:26]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_51));
defparam desc2462.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2463(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_47),.I4(N_51),.I5(N_85),.O(N_112));
defparam desc2463.INIT=64'h7775575522200200;
  LUT6 un4_s_lost_ac0_1_cZ(.I0(s_shr1[0:0]),.I1(s_shr1[1:1]),.I2(N_271),.I3(v_count[1:1]),.I4(m26_i),.I5(s_roundup),.O(un4_s_lost_ac0_1));
defparam un4_s_lost_ac0_1_cZ.INIT=64'h8421000088220000;
  LUT6 un4_s_lost_c5_RNO(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(un2_s_lost_0_c2),.I4(N_271),.I5(s_roundup),.O(un2_s_lost[2:2]));
defparam un4_s_lost_c5_RNO.INIT=64'hAAAA6AAAAAAAAAAA;
  LUT5 un4_s_lost_ac0_2_cZ(.I0(s_shr1[0:0]),.I1(s_shr1[1:1]),.I2(N_271),.I3(v_count[1:1]),.I4(s_roundup),.O(un4_s_lost_ac0_2));
defparam un4_s_lost_ac0_2_cZ.INIT=32'h00C600CC;
  FD desc2464(.Q(s_shl1),.D(s_shl1_0_0),.C(clk_i));
  LUT5_L desc2465(.I0(s_qutnt_i[7:7]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_117),.LO(s_fraco1_3[8:8]));
defparam desc2465.INIT=32'h8B0F8800;
  LUT5_L desc2466(.I0(s_qutnt_i[8:8]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_118),.LO(s_fraco1_3[9:9]));
defparam desc2466.INIT=32'h8B0F8800;
  LUT5_L desc2467(.I0(s_qutnt_i[9:9]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_119),.LO(s_fraco1_3[10:10]));
defparam desc2467.INIT=32'h8B0F8800;
  LUT5_L desc2468(.I0(s_qutnt_i[0:0]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_110),.LO(s_fraco1_3[1:1]));
defparam desc2468.INIT=32'h8B0F8800;
  LUT5_L desc2469(.I0(s_qutnt_i[1:1]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_111),.LO(s_fraco1_3[2:2]));
defparam desc2469.INIT=32'h8B0F8800;
  LUT5_L desc2470(.I0(s_qutnt_i[2:2]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_112),.LO(s_fraco1_3[3:3]));
defparam desc2470.INIT=32'h8B0F8800;
  LUT5_L desc2471(.I0(s_qutnt_i[6:6]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_116),.LO(s_fraco1_3[7:7]));
defparam desc2471.INIT=32'h8B0F8800;
  LUT5_L desc2472(.I0(s_qutnt_i[5:5]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_115),.LO(s_fraco1_3[6:6]));
defparam desc2472.INIT=32'h8B0F8800;
  LUT5_L desc2473(.I0(s_qutnt_i[4:4]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_114_0),.LO(s_fraco1_3[5:5]));
defparam desc2473.INIT=32'h8B0F8800;
  LUT5_L desc2474(.I0(s_qutnt_i[3:3]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_113),.LO(s_fraco1_3[4:4]));
defparam desc2474.INIT=32'h8B0F8800;
  LUT2 desc2475(.I0(s_rmndr_i[0:0]),.I1(s_rmndr_i[1:1]),.O(result_3_1_2));
defparam desc2475.INIT=4'hE;
  LUT2 desc2476(.I0(s_qutnt_i[0:0]),.I1(s_qutnt_i[1:1]),.O(N_1461_1));
defparam desc2476.INIT=4'h1;
  LUT2 un6_s_frac_rnd_1_s_34_RNO(.I0(s_expo1[8:8]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_1_axb_34));
defparam un6_s_frac_rnd_1_s_34_RNO.INIT=4'h9;
  LUT2 un6_s_frac_rnd_0_s_34_RNO(.I0(s_expo1[8:8]),.I1(s_fraco1[26:26]),.O(un6_s_frac_rnd_0_axb_34));
defparam un6_s_frac_rnd_0_s_34_RNO.INIT=4'h9;
  LUT2 desc2477(.I0(s_qutnt_i[8:8]),.I1(s_qutnt_i[9:9]),.O(N_1428));
defparam desc2477.INIT=4'hE;
  LUT2 desc2478(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[17:17]),.O(N_1429));
defparam desc2478.INIT=4'hE;
  LUT2 desc2479(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[11:11]),.O(N_55));
defparam desc2479.INIT=4'hE;
  LUT2 desc2480(.I0(s_qutnt_i[18:18]),.I1(s_qutnt_i[19:19]),.O(N_1421));
defparam desc2480.INIT=4'hE;
  LUT2 desc2481(.I0(s_qutnt_i[12:12]),.I1(s_qutnt_i[13:13]),.O(N_1420));
defparam desc2481.INIT=4'hE;
  LUT2 desc2482(.I0(s_qutnt_i[20:20]),.I1(s_qutnt_i[21:21]),.O(N_1487));
defparam desc2482.INIT=4'h1;
  LUT2 desc2483(.I0(s_qutnt_i[4:4]),.I1(s_qutnt_i[5:5]),.O(N_1479));
defparam desc2483.INIT=4'h1;
  LUT3 desc2484(.I0(s_qutnt_i[25:25]),.I1(s_qutnt_i[26:26]),.I2(s_shr1[0:0]),.O(N_26));
defparam desc2484.INIT=8'hCA;
  LUT3_L s_infb_0_cZ(.I0(s_opb_i[23:23]),.I1(s_opb_i_1),.I2(s_opb_i_2),.LO(s_infb_0));
defparam s_infb_0_cZ.INIT=8'h80;
  LUT4 desc2485(.I0(s_fractb_i[16:16]),.I1(s_fractb_i[17:17]),.I2(s_fractb_i[18:18]),.I3(s_fractb_i[19:19]),.O(result_5_20));
defparam desc2485.INIT=16'hFFFE;
  LUT4 desc2486(.I0(s_fracta_i[18:18]),.I1(s_fracta_i[19:19]),.I2(s_fracta_i[16:16]),.I3(s_fracta_i[17:17]),.O(result_16));
defparam desc2486.INIT=16'hFFFE;
  LUT6 desc2487(.I0(s_fractb_i[16:16]),.I1(s_fractb_i[17:17]),.I2(s_fractb_i[18:18]),.I3(s_fractb_i[19:19]),.I4(s_opb_i_5),.I5(s_opb_i_6),.O(result_5_1_0));
defparam desc2487.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2488(.I0(s_opb_i[23:23]),.I1(s_fractb_i[22:22]),.I2(s_opb_i_1),.I3(s_opb_i_2),.I4(s_opb_i_3),.I5(s_opb_i_4),.O(result_5_0));
defparam desc2488.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2489(.I0(s_rmndr_i[12:12]),.I1(s_rmndr_i[13:13]),.I2(s_rmndr_i[14:14]),.I3(s_rmndr_i[15:15]),.I4(s_rmndr_i[24:24]),.I5(s_rmndr_i[26:26]),.O(result_3_3));
defparam desc2489.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc2490(.I0(s_rmndr_i[6:6]),.I1(s_rmndr_i[7:7]),.I2(s_rmndr_i[8:8]),.I3(s_rmndr_i[9:9]),.I4(s_rmndr_i[10:10]),.I5(s_rmndr_i[11:11]),.LO(result_3_2));
defparam desc2490.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2491(.I0(s_rmndr_i[18:18]),.I1(s_rmndr_i[19:19]),.I2(s_rmndr_i[20:20]),.I3(s_rmndr_i[21:21]),.I4(s_rmndr_i[22:22]),.I5(s_rmndr_i[23:23]),.O(result_3_0));
defparam desc2491.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2492(.I0(s_fractb_i[6:6]),.I1(s_fractb_i[7:7]),.I2(s_fractb_i[8:8]),.I3(s_fractb_i[9:9]),.I4(s_fractb_i[10:10]),.I5(s_fractb_i[11:11]),.O(result_1_21_1));
defparam desc2492.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2493(.I0(s_fractb_i[0:0]),.I1(s_fractb_i[1:1]),.I2(s_fractb_i[2:2]),.I3(s_fractb_i[3:3]),.I4(s_fractb_i[4:4]),.I5(s_fractb_i[5:5]),.O(result_1_21_0));
defparam desc2493.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT5 desc2494(.I0(s_expo3[1:1]),.I1(s_expo3[2:2]),.I2(s_expo3[4:4]),.I3(s_expo3[5:5]),.I4(s_expo3[6:6]),.O(result_3));
defparam desc2494.INIT=32'h80000000;
  LUT5 desc2495(.I0(s_qutnt_i[1:1]),.I1(s_qutnt_i[2:2]),.I2(s_qutnt_i[3:3]),.I3(s_shr1[0:0]),.I4(s_shr1[1:1]),.O(N_28));
defparam desc2495.INIT=32'hF0CCAAAA;
  LUT6 desc2496(.I0(s_qutnt_i[4:4]),.I1(s_qutnt_i[6:6]),.I2(s_qutnt_i[5:5]),.I3(s_qutnt_i[3:3]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_31));
defparam desc2496.INIT=64'hCCCCF0F0AAAAFF00;
  LUT6 desc2497(.I0(s_qutnt_i[19:19]),.I1(s_qutnt_i[20:20]),.I2(s_qutnt_i[21:21]),.I3(s_qutnt_i[22:22]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_47));
defparam desc2497.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2498(.I0(s_qutnt_i[18:18]),.I1(s_qutnt_i[19:19]),.I2(s_qutnt_i[20:20]),.I3(s_qutnt_i[21:21]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_46));
defparam desc2498.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2499(.I0(s_qutnt_i[17:17]),.I1(s_qutnt_i[18:18]),.I2(s_qutnt_i[19:19]),.I3(s_qutnt_i[20:20]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_45));
defparam desc2499.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2500(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[17:17]),.I2(s_qutnt_i[18:18]),.I3(s_qutnt_i[19:19]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_44));
defparam desc2500.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2501(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[17:17]),.I2(s_qutnt_i[18:18]),.I3(s_qutnt_i[15:15]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_43));
defparam desc2501.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc2502(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[17:17]),.I2(s_qutnt_i[14:14]),.I3(s_qutnt_i[15:15]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_42));
defparam desc2502.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc2503(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[13:13]),.I2(s_qutnt_i[14:14]),.I3(s_qutnt_i[15:15]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_41));
defparam desc2503.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc2504(.I0(s_qutnt_i[12:12]),.I1(s_qutnt_i[13:13]),.I2(s_qutnt_i[14:14]),.I3(s_qutnt_i[15:15]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_40));
defparam desc2504.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2505(.I0(s_qutnt_i[11:11]),.I1(s_qutnt_i[12:12]),.I2(s_qutnt_i[13:13]),.I3(s_qutnt_i[14:14]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_39));
defparam desc2505.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2506(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[11:11]),.I2(s_qutnt_i[12:12]),.I3(s_qutnt_i[13:13]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_38));
defparam desc2506.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2507(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[11:11]),.I2(s_qutnt_i[9:9]),.I3(s_qutnt_i[12:12]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_37));
defparam desc2507.INIT=64'hFF00CCCCAAAAF0F0;
  LUT6 desc2508(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[11:11]),.I2(s_qutnt_i[8:8]),.I3(s_qutnt_i[9:9]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_36));
defparam desc2508.INIT=64'hCCCCAAAAFF00F0F0;
  LUT6 desc2509(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[7:7]),.I2(s_qutnt_i[8:8]),.I3(s_qutnt_i[9:9]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_35));
defparam desc2509.INIT=64'hAAAAFF00F0F0CCCC;
  LUT6 desc2510(.I0(s_qutnt_i[6:6]),.I1(s_qutnt_i[7:7]),.I2(s_qutnt_i[8:8]),.I3(s_qutnt_i[9:9]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_34));
defparam desc2510.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2511(.I0(s_qutnt_i[6:6]),.I1(s_qutnt_i[7:7]),.I2(s_qutnt_i[8:8]),.I3(s_qutnt_i[5:5]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_33));
defparam desc2511.INIT=64'hF0F0CCCCAAAAFF00;
  LUT6 desc2512(.I0(s_qutnt_i[4:4]),.I1(s_qutnt_i[6:6]),.I2(s_qutnt_i[7:7]),.I3(s_qutnt_i[5:5]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_32));
defparam desc2512.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc2513(.I0(s_qutnt_i[2:2]),.I1(s_qutnt_i[4:4]),.I2(s_qutnt_i[5:5]),.I3(s_qutnt_i[3:3]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_30));
defparam desc2513.INIT=64'hF0F0CCCCFF00AAAA;
  LUT6 desc2514(.I0(s_qutnt_i[1:1]),.I1(s_qutnt_i[2:2]),.I2(s_qutnt_i[4:4]),.I3(s_qutnt_i[3:3]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_29));
defparam desc2514.INIT=64'hF0F0FF00CCCCAAAA;
  LUT6 desc2515(.I0(s_qutnt_i[22:22]),.I1(s_qutnt_i[23:23]),.I2(s_qutnt_i[24:24]),.I3(s_qutnt_i[25:25]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_50));
defparam desc2515.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2516(.I0(s_qutnt_i[21:21]),.I1(s_qutnt_i[22:22]),.I2(s_qutnt_i[23:23]),.I3(s_qutnt_i[24:24]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_49));
defparam desc2516.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2517(.I0(s_qutnt_i[20:20]),.I1(s_qutnt_i[21:21]),.I2(s_qutnt_i[22:22]),.I3(s_qutnt_i[23:23]),.I4(s_shr1[0:0]),.I5(s_shr1[1:1]),.O(N_48));
defparam desc2517.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 desc2518(.I0(s_rmndr_i[2:2]),.I1(s_rmndr_i[3:3]),.I2(s_rmndr_i[4:4]),.I3(s_rmndr_i[5:5]),.I4(result_3_1_2),.I5(result_3_2),.O(result_3_2_4));
defparam desc2518.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 s_infb_c(.I0(s_opb_i_3),.I1(s_opb_i_4),.I2(s_opb_i_5),.I3(s_opb_i_6),.I4(s_opb_i_7),.I5(s_infb_0),.O(s_infb));
defparam s_infb_c.INIT=64'h8000000000000000;
  LUT6 un1_s_infa_c(.I0(s_opa_i_3),.I1(s_opa_i_4),.I2(s_opa_i_5),.I3(s_opa_i_6),.I4(s_opa_i_7),.I5(un1_s_infa_0),.O(un1_s_infa));
defparam un1_s_infa_c.INIT=64'h8000000000000000;
  LUT6 desc2519(.I0(s_qutnt_i[0:0]),.I1(s_qutnt_i[1:1]),.I2(s_qutnt_i[2:2]),.I3(s_qutnt_i[6:6]),.I4(s_qutnt_i[5:5]),.I5(s_qutnt_i[3:3]),.O(m26_i_1));
defparam desc2519.INIT=64'hBABABABABABABBBA;
  LUT6_L desc2520(.I0(N_1424),.I1(N_1487),.I2(N_55),.I3(N_1428),.I4(N_1480),.I5(N_1426),.LO(N_1416_2));
defparam desc2520.INIT=64'hFFF00000FFF40000;
  LUT5 desc2521(.I0(s_rmndr_i[16:16]),.I1(s_rmndr_i[17:17]),.I2(s_rmndr_i[25:25]),.I3(result_3_0),.I4(result_3_3),.O(result_3_3_4));
defparam desc2521.INIT=32'hFFFFFFFE;
  LUT6 desc2522(.I0(s_fractb_i[12:12]),.I1(s_fractb_i[13:13]),.I2(s_fractb_i[14:14]),.I3(s_fractb_i[15:15]),.I4(result_1_21_0),.I5(result_1_21_1),.O(result_5_28));
defparam desc2522.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT5 desc2523(.I0(s_shr1[1:1]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_26),.I4(N_49),.O(N_103));
defparam desc2523.INIT=32'h13031000;
  LUT4 desc2524(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_47),.I3(N_51),.O(N_101));
defparam desc2524.INIT=16'h5410;
  LUT6 desc2525(.I0(N_1421),.I1(N_1429),.I2(N_1433),.I3(N_1480),.I4(N_1426),.I5(N_1416_2),.O(m73_i));
defparam desc2525.INIT=64'hFFFFFFFFF0F0FEF0;
  LUT6 desc2526(.I0(s_qutnt_i[2:2]),.I1(s_qutnt_i[3:3]),.I2(N_1422),.I3(N_1479),.I4(N_55),.I5(N_1428),.O(N_1437));
defparam desc2526.INIT=64'hFEEEFEEEFFEEFEEE;
  LUT6 desc2527(.I0(s_fractb_i[20:20]),.I1(s_fractb_i[21:21]),.I2(s_opb_i_7),.I3(result_5_0),.I4(result_5_1_0),.I5(result_5_28),.O(result_5));
defparam desc2527.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 desc2528(.I0(s_fracta_i[22:22]),.I1(s_opa_i[23:23]),.I2(result_4_0_3),.I3(result_3_21_1),.I4(result_4_2),.I5(result_3_21_3),.O(result_4));
defparam desc2528.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L desc2529(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_36),.I3(N_44),.I4(N_40),.I5(N_48),.LO(N_90));
defparam desc2529.INIT=64'hFEDCBA9876543210;
  LUT6_L desc2530(.I0(N_114),.I1(N_1419),.I2(N_1421),.I3(N_1424),.I4(N_1429),.I5(N_1487),.LO(N_1431));
defparam desc2530.INIT=64'hCCCCFFFECCCCFCFC;
  LUT6 desc2531(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_28),.I3(N_32),.I4(N_36),.I5(N_40),.O(N_82));
defparam desc2531.INIT=64'hFEBADC9876325410;
  LUT6 desc2532(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_30),.I3(N_34),.I4(N_38),.I5(N_42),.O(N_84));
defparam desc2532.INIT=64'hFEBADC9876325410;
  LUT6_L desc2533(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_31),.I3(N_35),.I4(N_39),.I5(N_43),.LO(N_85));
defparam desc2533.INIT=64'hFEBADC9876325410;
  LUT6_L desc2534(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_38),.I3(N_42),.I4(N_46),.I5(N_50),.LO(N_92));
defparam desc2534.INIT=64'hFEBADC9876325410;
  LUT6_L desc2535(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_37),.I3(N_41),.I4(N_45),.I5(N_49),.LO(N_91));
defparam desc2535.INIT=64'hFEBADC9876325410;
  LUT6_L desc2536(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_35),.I3(N_39),.I4(N_43),.I5(N_47),.LO(N_89));
defparam desc2536.INIT=64'hFEBADC9876325410;
  LUT6_L desc2537(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_34),.I3(N_38),.I4(N_42),.I5(N_46),.LO(N_88));
defparam desc2537.INIT=64'hFEBADC9876325410;
  LUT6_L desc2538(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_32),.I3(N_36),.I4(N_44),.I5(N_40),.LO(N_86));
defparam desc2538.INIT=64'hFEBA7632DC985410;
  LUT6 desc2539(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_29),.I3(N_33),.I4(N_37),.I5(N_41),.O(N_83));
defparam desc2539.INIT=64'hFEBADC9876325410;
  LUT5 desc2540(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_54),.I3(N_46),.I4(N_50),.O(N_100));
defparam desc2540.INIT=32'h75643120;
  LUT6 desc2541(.I0(s_shr1[1:1]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_26),.I4(N_45),.I5(N_49),.O(N_99));
defparam desc2541.INIT=64'h3733343007030400;
  LUT5 desc2542(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_43),.I3(N_47),.I4(N_51),.O(N_97));
defparam desc2542.INIT=32'h76325410;
  LUT6 desc2543(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_54),.I3(N_42),.I4(N_46),.I5(N_50),.O(N_96));
defparam desc2543.INIT=64'hF7E6B3A2D5C49180;
  LUT6 desc2544(.I0(s_shr1[1:1]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_26),.I4(N_49),.I5(N_68),.O(N_95));
defparam desc2544.INIT=64'h7F3F73334C0C4000;
  LUT6 desc2545(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_52),.I3(N_44),.I4(N_40),.I5(N_48),.O(N_94));
defparam desc2545.INIT=64'hF7B3E6A2D591C480;
  LUT6 desc2546(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_39),.I3(N_43),.I4(N_47),.I5(N_51),.O(N_93));
defparam desc2546.INIT=64'hFEBADC9876325410;
  LUT6 desc2547(.I0(N_1421),.I1(N_1424),.I2(N_1429),.I3(N_1487),.I4(N_1488),.I5(v_count_1[3:3]),.O(v_count[3:3]));
defparam desc2547.INIT=64'hFFFFFFFF01000000;
  LUT6 un6_s_inf_result_cZ(.I0(s_expo3[8:8]),.I1(s_expo3[0:0]),.I2(s_expo3[3:3]),.I3(s_expo3[7:7]),.I4(result_3),.I5(result_5),.O(un6_s_inf_result));
defparam un6_s_inf_result_cZ.INIT=64'hEAAAAAAAFFFFFFFF;
  LUT6 un1_s_nan_a_c(.I0(s_fracta_i[22:22]),.I1(result_11),.I2(result_16),.I3(result_3_21_1),.I4(result_3_21_3),.I5(un1_s_infa),.O(un1_s_nan_a));
defparam un1_s_nan_a_c.INIT=64'hFFFFFFFE00000000;
  LUT6 un1_s_nan_b_c(.I0(s_fractb_i[20:20]),.I1(s_fractb_i[21:21]),.I2(s_fractb_i[22:22]),.I3(result_5_20),.I4(result_5_28),.I5(s_infb),.O(un1_s_nan_b));
defparam un1_s_nan_b_c.INIT=64'hFFFFFFFE00000000;
  LUT2 un6_s_op_0(.I0(result_5),.I1(result_4),.O(un3_s_op_0));
defparam un6_s_op_0.INIT=4'h8;
  LUT3 desc2548(.I0(s_shr1[4:4]),.I1(N_108),.I2(N_92),.O(N_119));
defparam desc2548.INIT=8'hD8;
  LUT5 desc2549(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(N_60),.I3(N_103),.I4(N_68),.O(N_114_0));
defparam desc2549.INIT=32'hFE54BA10;
  LUT5 un16_s_roundup_cZ(.I0(s_fraco1[0:0]),.I1(s_fraco1[1:1]),.I2(s_fraco1[3:3]),.I3(result_3_2_4),.I4(result_3_3_4),.O(un16_s_roundup));
defparam un16_s_roundup_cZ.INIT=32'hFFFFFFFE;
  LUT6 desc2550(.I0(N_1461_1),.I1(N_1420),.I2(N_1479),.I3(N_1428),.I4(N_1437),.I5(N_1431),.O(v_count[1:1]));
defparam desc2550.INIT=64'hAAAA0020AAAA0000;
  LUT6_L desc2551(.I0(s_qutnt_i[18:18]),.I1(s_qutnt_i[19:19]),.I2(s_qutnt_i[20:20]),.I3(s_qutnt_i[21:21]),.I4(s_qutnt_i[22:22]),.I5(N_123),.LO(N_148));
defparam desc2551.INIT=64'h4544454445444545;
  LUT6 un7_s_nan_in_cZ(.I0(s_infb),.I1(un1_s_infa),.I2(result_5),.I3(un1_s_nan_b),.I4(result_4),.I5(un1_s_nan_a),.O(un7_s_nan_in));
defparam un7_s_nan_in_cZ.INIT=64'hFFFFFFFFFF88FF8F;
  LUT6 s_exp_10b_axbxc4(.I0(s_exp_10_i[4:4]),.I1(s_exp_10_i[3:3]),.I2(s_exp_10_i[2:2]),.I3(s_exp_10_i[1:1]),.I4(s_exp_10_i[0:0]),.I5(s_qutnt_i[26:26]),.O(s_exp_10b[4:4]));
defparam s_exp_10b_axbxc4.INIT=64'hAAAAAAAAAAAAAAA9;
  LUT5 v_shr_1_c4_cZ(.I0(s_exp_10_i[3:3]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_qutnt_i[26:26]),.O(v_shr_1_c4));
defparam v_shr_1_c4_cZ.INIT=32'hFEFEFEFF;
  LUT6 s_exp_10b_c5_cZ(.I0(s_exp_10_i[4:4]),.I1(s_exp_10_i[3:3]),.I2(s_exp_10_i[2:2]),.I3(s_exp_10_i[1:1]),.I4(s_exp_10_i[0:0]),.I5(s_qutnt_i[26:26]),.O(s_exp_10b_c5));
defparam s_exp_10b_c5_cZ.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT5_L desc2552(.I0(s_qutnt_i[0:0]),.I1(s_shl1),.I2(s_shr1[5:5]),.I3(un1_s_shr1_1),.I4(N_109),.LO(s_fraco1_3[0:0]));
defparam desc2552.INIT=32'h220F2200;
  LUT6 s_roundup_3(.I0(s_sign_i),.I1(s_fraco1[2:2]),.I2(s_rmode_i[0:0]),.I3(s_rmode_i[1:1]),.I4(un16_s_roundup),.I5(un18_s_roundup),.O(s_roundup));
defparam s_roundup_3.INIT=64'hA50CA500000C0000;
  LUT6_L desc2553(.I0(s_qutnt_i[16:16]),.I1(s_qutnt_i[17:17]),.I2(s_qutnt_i[13:13]),.I3(s_qutnt_i[14:14]),.I4(s_qutnt_i[15:15]),.I5(N_148),.LO(N_1483));
defparam desc2553.INIT=64'h0F000F0A0F000F0B;
  LUT3_L desc2554(.I0(s_fraco1[21:21]),.I1(un6_s_frac_rnd1[18:18]),.I2(s_roundup),.LO(s_frac_rnd[18:18]));
defparam desc2554.INIT=8'hCA;
  LUT6 un1_s_ine_o_RNO(.I0(s_shr1[5:5]),.I1(s_shr1[4:4]),.I2(s_shr1[3:3]),.I3(s_shr1[2:2]),.I4(un2_s_lost_0_c2),.I5(N_27),.O(un2_s_lost[1:1]));
defparam un1_s_ine_o_RNO.INIT=64'hAAAAAAAA6AAAAAAA;
  LUT6 s_exp_10b_axbxc7_lut6_2_RNIQA981_cZ(.I0(s_exp_10b[1:1]),.I1(s_exp_10b[2:2]),.I2(s_exp_10b[3:3]),.I3(s_exp_10b[4:4]),.I4(s_exp_10b[5:5]),.I5(s_exp_10b[7:7]),.O(s_exp_10b_axbxc7_lut6_2_RNIQA981));
defparam s_exp_10b_axbxc7_lut6_2_RNIQA981_cZ.INIT=64'h0000000000000001;
  LUT5 s_exp_10b_axbxc8(.I0(s_exp_10_i[8:8]),.I1(s_exp_10_i[7:7]),.I2(s_exp_10_i[6:6]),.I3(s_exp_10_i[5:5]),.I4(s_exp_10b_c5),.O(s_exp_10b[8:8]));
defparam s_exp_10b_axbxc8.INIT=32'hAAAAAAA9;
  LUT6_L desc2555(.I0(s_qutnt_i[10:10]),.I1(s_qutnt_i[11:11]),.I2(s_qutnt_i[8:8]),.I3(s_qutnt_i[9:9]),.I4(s_qutnt_i[12:12]),.I5(N_1483),.LO(N_1455));
defparam desc2555.INIT=64'hF0FBF0FBF0FBF0FA;
  LUT6 s_exp_10b_axbxc9(.I0(s_exp_10_i[9:9]),.I1(s_exp_10_i[8:8]),.I2(s_exp_10_i[7:7]),.I3(s_exp_10_i[6:6]),.I4(s_exp_10_i[5:5]),.I5(s_exp_10b_c5),.O(s_exp_10b[9:9]));
defparam s_exp_10b_axbxc9.INIT=64'hAAAAAAAAAAAAAAA9;
  LUT6 desc2556(.I0(s_qutnt_i[4:4]),.I1(s_qutnt_i[7:7]),.I2(s_qutnt_i[5:5]),.I3(N_1423),.I4(m26_i_1),.I5(N_1455),.O(m26_i));
defparam desc2556.INIT=64'hFFFF00ABFFFF00AA;
  LUT6 desc2557(.I0(s_exp_10_i[9:9]),.I1(s_exp_10_i[8:8]),.I2(s_exp_10_i[7:7]),.I3(s_exp_10_i[6:6]),.I4(s_exp_10_i[5:5]),.I5(s_exp_10b_c5),.O(s_expo1_3[6:6]));
defparam desc2557.INIT=64'h5500550055000056;
  LUT6 s_exp_10b_axbxc8_RNIGLJC4_cZ(.I0(s_exp_10_i[0:0]),.I1(s_qutnt_i[26:26]),.I2(s_exp_10b[8:8]),.I3(s_expo1_3[6:6]),.I4(s_exp_10b[9:9]),.I5(s_exp_10b_axbxc7_lut6_2_RNIQA981),.O(s_exp_10b_axbxc8_RNIGLJC4));
defparam s_exp_10b_axbxc8_RNIGLJC4_cZ.INIT=64'h0600FFF90000FFFF;
  LUT6_L un4_s_lost_c3_cZ(.I0(s_shr1[2:2]),.I1(un2_s_lost_0_c2),.I2(m73_i),.I3(un4_s_lost_ac0_1),.I4(un4_s_lost_ac0_2),.I5(N_27),.LO(un4_s_lost_c3));
defparam un4_s_lost_c3_cZ.INIT=64'hFAFAFAA0F6F6F660;
  LUT6_L desc2558(.I0(s_exp_10_i[0:0]),.I1(s_qutnt_i[26:26]),.I2(s_exp_10b[8:8]),.I3(s_expo1_3[6:6]),.I4(s_exp_10b[9:9]),.I5(s_exp_10b_axbxc7_lut6_2_RNIQA981),.LO(N_1357_i));
defparam desc2558.INIT=64'hF9FF999FFFFF9999;
  LUT6 v_shr_1_c4_RNIEPFK5(.I0(s_exp_10_i[6:6]),.I1(s_exp_10_i[5:5]),.I2(v_shr_1_c4),.I3(s_exp_10b[4:4]),.I4(s_exp_10b_c5),.I5(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[6:6]));
defparam v_shr_1_c4_RNIEPFK5.INIT=64'h000000005556666A;
  LUT6_L desc2559(.I0(s_exp_10_i[0:0]),.I1(s_qutnt_i[26:26]),.I2(s_exp_10b[8:8]),.I3(s_expo1_3[6:6]),.I4(s_exp_10b[9:9]),.I5(s_exp_10b_axbxc7_lut6_2_RNIQA981),.LO(v_shr_2[0:0]));
defparam desc2559.INIT=64'h5155000455550000;
  LUT6_L un4_s_lost_c4_cZ(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(un2_s_lost_0_c2),.I3(v_count[3:3]),.I4(N_27),.I5(un4_s_lost_c3),.LO(un4_s_lost_c4));
defparam un4_s_lost_c4_cZ.INIT=64'hAAFF6AFF00AA006A;
  LUT6_L un4_s_lost_c5_cZ(.I0(N_55),.I1(N_1428),.I2(N_1426),.I3(N_1488),.I4(un2_s_lost[2:2]),.I5(un4_s_lost_c4),.LO(un4_s_lost_c5));
defparam un4_s_lost_c5_cZ.INIT=64'hFFFFFEFFFEFF0000;
  LUT6_L un1_s_ine_o(.I0(un4_s_ine_o_1),.I1(un6_s_infa),.I2(un3_s_op_0),.I3(un6_s_inf_result),.I4(un2_s_lost[1:1]),.I5(un4_s_lost_c5),.LO(un1_s_ine_o_0));
defparam un1_s_ine_o.INIT=64'hF0F0F0F0F0F0B0A0;
  XORCY un6_s_frac_rnd_1_s_34(.LI(un6_s_frac_rnd_1_axb_34),.CI(un6_s_frac_rnd_1_cry_33),.O(s_expo3_31[8:8]));
  XORCY un6_s_frac_rnd_1_s_33(.LI(un6_s_frac_rnd_1_axb_33),.CI(un6_s_frac_rnd_1_cry_32),.O(s_expo3_31[7:7]));
  MUXCY_L un6_s_frac_rnd_1_cry_33_cZ(.DI(s_expo1[7:7]),.CI(un6_s_frac_rnd_1_cry_32),.S(un6_s_frac_rnd_1_axb_33),.LO(un6_s_frac_rnd_1_cry_33));
  XORCY un6_s_frac_rnd_1_s_32(.LI(un6_s_frac_rnd_1_axb_32),.CI(un6_s_frac_rnd_1_cry_31),.O(s_expo3_31[6:6]));
  MUXCY_L un6_s_frac_rnd_1_cry_32_cZ(.DI(s_expo1[6:6]),.CI(un6_s_frac_rnd_1_cry_31),.S(un6_s_frac_rnd_1_axb_32),.LO(un6_s_frac_rnd_1_cry_32));
  XORCY un6_s_frac_rnd_1_s_31(.LI(un6_s_frac_rnd_1_axb_31),.CI(un6_s_frac_rnd_1_cry_30),.O(s_expo3_31[5:5]));
  MUXCY_L un6_s_frac_rnd_1_cry_31_cZ(.DI(s_expo1[5:5]),.CI(un6_s_frac_rnd_1_cry_30),.S(un6_s_frac_rnd_1_axb_31),.LO(un6_s_frac_rnd_1_cry_31));
  XORCY un6_s_frac_rnd_1_s_30(.LI(un6_s_frac_rnd_1_axb_30),.CI(un6_s_frac_rnd_1_cry_29),.O(s_expo3_31[4:4]));
  MUXCY_L un6_s_frac_rnd_1_cry_30_cZ(.DI(s_expo1[4:4]),.CI(un6_s_frac_rnd_1_cry_29),.S(un6_s_frac_rnd_1_axb_30),.LO(un6_s_frac_rnd_1_cry_30));
  XORCY un6_s_frac_rnd_1_s_29(.LI(un6_s_frac_rnd_1_axb_29),.CI(un6_s_frac_rnd_1_cry_28),.O(s_expo3_31[3:3]));
  MUXCY_L un6_s_frac_rnd_1_cry_29_cZ(.DI(s_expo1[3:3]),.CI(un6_s_frac_rnd_1_cry_28),.S(un6_s_frac_rnd_1_axb_29),.LO(un6_s_frac_rnd_1_cry_29));
  XORCY un6_s_frac_rnd_1_s_28(.LI(un6_s_frac_rnd_1_axb_28),.CI(un6_s_frac_rnd_1_cry_27),.O(s_expo3_31[2:2]));
  MUXCY_L un6_s_frac_rnd_1_cry_28_cZ(.DI(s_expo1[2:2]),.CI(un6_s_frac_rnd_1_cry_27),.S(un6_s_frac_rnd_1_axb_28),.LO(un6_s_frac_rnd_1_cry_28));
  XORCY un6_s_frac_rnd_1_s_27(.LI(un6_s_frac_rnd_1_axb_27),.CI(un6_s_frac_rnd_1_cry_26),.O(s_expo3_31[1:1]));
  MUXCY_L un6_s_frac_rnd_1_cry_27_cZ(.DI(s_expo1[1:1]),.CI(un6_s_frac_rnd_1_cry_26),.S(un6_s_frac_rnd_1_axb_27),.LO(un6_s_frac_rnd_1_cry_27));
  XORCY un6_s_frac_rnd_1_s_26(.LI(un6_s_frac_rnd_1_axb_26),.CI(un6_s_frac_rnd_1_cry_25),.O(s_expo3_31[0:0]));
  MUXCY_L un6_s_frac_rnd_1_cry_26_cZ(.DI(s_expo1[0:0]),.CI(un6_s_frac_rnd_1_cry_25),.S(un6_s_frac_rnd_1_axb_26),.LO(un6_s_frac_rnd_1_cry_26));
  XORCY un6_s_frac_rnd_1_s_25(.LI(un6_s_frac_rnd_1_axb_25),.CI(un6_s_frac_rnd_1_cry_24),.O(N_271));
  MUXCY_L un6_s_frac_rnd_1_cry_25_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_24),.S(un6_s_frac_rnd_1_axb_25),.LO(un6_s_frac_rnd_1_cry_25));
  MUXCY_L un6_s_frac_rnd_1_cry_23(.DI(GND),.CI(un6_s_frac_rnd_1_cry_22),.S(un6_s_frac_rnd_1_axb_23),.LO(un6_s_frac_rnd_1_cry_24));
  XORCY un6_s_frac_rnd_1_s_22(.LI(un6_s_frac_rnd_1_axb_22),.CI(un6_s_frac_rnd_1_cry_21),.O(un6_s_frac_rnd1[22:22]));
  MUXCY_L un6_s_frac_rnd_1_cry_22_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_21),.S(un6_s_frac_rnd_1_axb_22),.LO(un6_s_frac_rnd_1_cry_22));
  XORCY un6_s_frac_rnd_1_s_21(.LI(un6_s_frac_rnd_1_axb_21),.CI(un6_s_frac_rnd_1_cry_20),.O(un6_s_frac_rnd1[21:21]));
  MUXCY_L un6_s_frac_rnd_1_cry_21_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_20),.S(un6_s_frac_rnd_1_axb_21),.LO(un6_s_frac_rnd_1_cry_21));
  XORCY un6_s_frac_rnd_1_s_20(.LI(un6_s_frac_rnd_1_axb_20),.CI(un6_s_frac_rnd_1_cry_19),.O(un6_s_frac_rnd1[20:20]));
  MUXCY_L un6_s_frac_rnd_1_cry_20_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_19),.S(un6_s_frac_rnd_1_axb_20),.LO(un6_s_frac_rnd_1_cry_20));
  XORCY un6_s_frac_rnd_1_s_19(.LI(un6_s_frac_rnd_1_axb_19),.CI(un6_s_frac_rnd_1_cry_18),.O(un6_s_frac_rnd1[19:19]));
  MUXCY_L un6_s_frac_rnd_1_cry_19_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_18),.S(un6_s_frac_rnd_1_axb_19),.LO(un6_s_frac_rnd_1_cry_19));
  XORCY un6_s_frac_rnd_1_s_18(.LI(un6_s_frac_rnd_1_axb_18),.CI(un6_s_frac_rnd_1_cry_17),.O(un6_s_frac_rnd1[18:18]));
  MUXCY_L un6_s_frac_rnd_1_cry_18_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_17),.S(un6_s_frac_rnd_1_axb_18),.LO(un6_s_frac_rnd_1_cry_18));
  XORCY un6_s_frac_rnd_1_s_17(.LI(un6_s_frac_rnd_1_axb_17),.CI(un6_s_frac_rnd_1_cry_16),.O(un6_s_frac_rnd1[17:17]));
  MUXCY_L un6_s_frac_rnd_1_cry_17_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_16),.S(un6_s_frac_rnd_1_axb_17),.LO(un6_s_frac_rnd_1_cry_17));
  XORCY un6_s_frac_rnd_1_s_16(.LI(un6_s_frac_rnd_1_axb_16),.CI(un6_s_frac_rnd_1_cry_15),.O(un6_s_frac_rnd1[16:16]));
  MUXCY_L un6_s_frac_rnd_1_cry_16_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_15),.S(un6_s_frac_rnd_1_axb_16),.LO(un6_s_frac_rnd_1_cry_16));
  XORCY un6_s_frac_rnd_1_s_15(.LI(un6_s_frac_rnd_1_axb_15),.CI(un6_s_frac_rnd_1_cry_14),.O(un6_s_frac_rnd1[15:15]));
  MUXCY_L un6_s_frac_rnd_1_cry_15_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_14),.S(un6_s_frac_rnd_1_axb_15),.LO(un6_s_frac_rnd_1_cry_15));
  XORCY un6_s_frac_rnd_1_s_14(.LI(un6_s_frac_rnd_1_axb_14),.CI(un6_s_frac_rnd_1_cry_13),.O(un6_s_frac_rnd1[14:14]));
  MUXCY_L un6_s_frac_rnd_1_cry_14_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_13),.S(un6_s_frac_rnd_1_axb_14),.LO(un6_s_frac_rnd_1_cry_14));
  XORCY un6_s_frac_rnd_1_s_13(.LI(un6_s_frac_rnd_1_axb_13),.CI(un6_s_frac_rnd_1_cry_12),.O(un6_s_frac_rnd1[13:13]));
  MUXCY_L un6_s_frac_rnd_1_cry_13_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_12),.S(un6_s_frac_rnd_1_axb_13),.LO(un6_s_frac_rnd_1_cry_13));
  XORCY un6_s_frac_rnd_1_s_12(.LI(un6_s_frac_rnd_1_axb_12),.CI(un6_s_frac_rnd_1_cry_11),.O(un6_s_frac_rnd1[12:12]));
  MUXCY_L un6_s_frac_rnd_1_cry_12_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_11),.S(un6_s_frac_rnd_1_axb_12),.LO(un6_s_frac_rnd_1_cry_12));
  XORCY un6_s_frac_rnd_1_s_11(.LI(un6_s_frac_rnd_1_axb_11),.CI(un6_s_frac_rnd_1_cry_10),.O(un6_s_frac_rnd1[11:11]));
  MUXCY_L un6_s_frac_rnd_1_cry_11_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_10),.S(un6_s_frac_rnd_1_axb_11),.LO(un6_s_frac_rnd_1_cry_11));
  XORCY un6_s_frac_rnd_1_s_10(.LI(un6_s_frac_rnd_1_axb_10),.CI(un6_s_frac_rnd_1_cry_9),.O(un6_s_frac_rnd1[10:10]));
  MUXCY_L un6_s_frac_rnd_1_cry_10_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_9),.S(un6_s_frac_rnd_1_axb_10),.LO(un6_s_frac_rnd_1_cry_10));
  XORCY un6_s_frac_rnd_1_s_9(.LI(un6_s_frac_rnd_1_axb_9),.CI(un6_s_frac_rnd_1_cry_8),.O(un6_s_frac_rnd1[9:9]));
  MUXCY_L un6_s_frac_rnd_1_cry_9_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_8),.S(un6_s_frac_rnd_1_axb_9),.LO(un6_s_frac_rnd_1_cry_9));
  XORCY un6_s_frac_rnd_1_s_8(.LI(un6_s_frac_rnd_1_axb_8),.CI(un6_s_frac_rnd_1_cry_7),.O(un6_s_frac_rnd1[8:8]));
  MUXCY_L un6_s_frac_rnd_1_cry_8_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_7),.S(un6_s_frac_rnd_1_axb_8),.LO(un6_s_frac_rnd_1_cry_8));
  XORCY un6_s_frac_rnd_1_s_7(.LI(un6_s_frac_rnd_1_axb_7),.CI(un6_s_frac_rnd_1_cry_6),.O(un6_s_frac_rnd1[7:7]));
  MUXCY_L un6_s_frac_rnd_1_cry_7_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_6),.S(un6_s_frac_rnd_1_axb_7),.LO(un6_s_frac_rnd_1_cry_7));
  XORCY un6_s_frac_rnd_1_s_6(.LI(un6_s_frac_rnd_1_axb_6),.CI(un6_s_frac_rnd_1_cry_5),.O(un6_s_frac_rnd1[6:6]));
  MUXCY_L un6_s_frac_rnd_1_cry_6_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_5),.S(un6_s_frac_rnd_1_axb_6),.LO(un6_s_frac_rnd_1_cry_6));
  XORCY un6_s_frac_rnd_1_s_5(.LI(un6_s_frac_rnd_1_axb_5),.CI(un6_s_frac_rnd_1_cry_4),.O(un6_s_frac_rnd1[5:5]));
  MUXCY_L un6_s_frac_rnd_1_cry_5_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_4),.S(un6_s_frac_rnd_1_axb_5),.LO(un6_s_frac_rnd_1_cry_5));
  XORCY un6_s_frac_rnd_1_s_4(.LI(un6_s_frac_rnd_1_axb_4),.CI(un6_s_frac_rnd_1_cry_3),.O(un6_s_frac_rnd1[4:4]));
  MUXCY_L un6_s_frac_rnd_1_cry_4_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_3),.S(un6_s_frac_rnd_1_axb_4),.LO(un6_s_frac_rnd_1_cry_4));
  XORCY un6_s_frac_rnd_1_s_3(.LI(un6_s_frac_rnd_1_axb_3),.CI(un6_s_frac_rnd_1_cry_2),.O(un6_s_frac_rnd1[3:3]));
  MUXCY_L un6_s_frac_rnd_1_cry_3_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_2),.S(un6_s_frac_rnd_1_axb_3),.LO(un6_s_frac_rnd_1_cry_3));
  XORCY un6_s_frac_rnd_1_s_2(.LI(un6_s_frac_rnd_1_axb_2),.CI(un6_s_frac_rnd_1_cry_1),.O(un6_s_frac_rnd1[2:2]));
  MUXCY_L un6_s_frac_rnd_1_cry_2_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_1),.S(un6_s_frac_rnd_1_axb_2),.LO(un6_s_frac_rnd_1_cry_2));
  XORCY un6_s_frac_rnd_1_s_1(.LI(un6_s_frac_rnd_1_axb_1),.CI(un6_s_frac_rnd_1_cry_0),.O(un6_s_frac_rnd1[1:1]));
  MUXCY_L un6_s_frac_rnd_1_cry_1_cZ(.DI(GND),.CI(un6_s_frac_rnd_1_cry_0),.S(un6_s_frac_rnd_1_axb_1),.LO(un6_s_frac_rnd_1_cry_1));
  MUXCY_L un6_s_frac_rnd_1_cry_0_cZ(.DI(VCC),.CI(GND),.S(un6_s_frac_rnd_1_cry_0_sf),.LO(un6_s_frac_rnd_1_cry_0));
  XORCY un6_s_frac_rnd_0_s_34(.LI(un6_s_frac_rnd_0_axb_34),.CI(un6_s_frac_rnd_0_cry_33),.O(s_expo3_30[8:8]));
  XORCY un6_s_frac_rnd_0_s_33(.LI(un6_s_frac_rnd_0_axb_33),.CI(un6_s_frac_rnd_0_cry_32),.O(s_expo3_30[7:7]));
  MUXCY_L un6_s_frac_rnd_0_cry_33_cZ(.DI(s_expo1[7:7]),.CI(un6_s_frac_rnd_0_cry_32),.S(un6_s_frac_rnd_0_axb_33),.LO(un6_s_frac_rnd_0_cry_33));
  XORCY un6_s_frac_rnd_0_s_32(.LI(un6_s_frac_rnd_0_axb_32),.CI(un6_s_frac_rnd_0_cry_31),.O(s_expo3_30[6:6]));
  MUXCY_L un6_s_frac_rnd_0_cry_32_cZ(.DI(s_expo1[6:6]),.CI(un6_s_frac_rnd_0_cry_31),.S(un6_s_frac_rnd_0_axb_32),.LO(un6_s_frac_rnd_0_cry_32));
  XORCY un6_s_frac_rnd_0_s_31(.LI(un6_s_frac_rnd_0_axb_31),.CI(un6_s_frac_rnd_0_cry_30),.O(s_expo3_30[5:5]));
  MUXCY_L un6_s_frac_rnd_0_cry_31_cZ(.DI(s_expo1[5:5]),.CI(un6_s_frac_rnd_0_cry_30),.S(un6_s_frac_rnd_0_axb_31),.LO(un6_s_frac_rnd_0_cry_31));
  XORCY un6_s_frac_rnd_0_s_30(.LI(un6_s_frac_rnd_0_axb_30),.CI(un6_s_frac_rnd_0_cry_29),.O(s_expo3_30[4:4]));
  MUXCY_L un6_s_frac_rnd_0_cry_30_cZ(.DI(s_expo1[4:4]),.CI(un6_s_frac_rnd_0_cry_29),.S(un6_s_frac_rnd_0_axb_30),.LO(un6_s_frac_rnd_0_cry_30));
  XORCY un6_s_frac_rnd_0_s_29(.LI(un6_s_frac_rnd_0_axb_29),.CI(un6_s_frac_rnd_0_cry_28),.O(s_expo3_30[3:3]));
  MUXCY_L un6_s_frac_rnd_0_cry_29_cZ(.DI(s_expo1[3:3]),.CI(un6_s_frac_rnd_0_cry_28),.S(un6_s_frac_rnd_0_axb_29),.LO(un6_s_frac_rnd_0_cry_29));
  XORCY un6_s_frac_rnd_0_s_28(.LI(un6_s_frac_rnd_0_axb_28),.CI(un6_s_frac_rnd_0_cry_27),.O(s_expo3_30[2:2]));
  MUXCY_L un6_s_frac_rnd_0_cry_28_cZ(.DI(s_expo1[2:2]),.CI(un6_s_frac_rnd_0_cry_27),.S(un6_s_frac_rnd_0_axb_28),.LO(un6_s_frac_rnd_0_cry_28));
  XORCY un6_s_frac_rnd_0_s_27(.LI(un6_s_frac_rnd_0_axb_27),.CI(un6_s_frac_rnd_0_cry_26),.O(s_expo3_30[1:1]));
  MUXCY_L un6_s_frac_rnd_0_cry_27_cZ(.DI(s_expo1[1:1]),.CI(un6_s_frac_rnd_0_cry_26),.S(un6_s_frac_rnd_0_axb_27),.LO(un6_s_frac_rnd_0_cry_27));
  MUXCY_L un6_s_frac_rnd_0_cry_26_cZ(.DI(s_expo1[0:0]),.CI(GND),.S(s_expo3_30[0:0]),.LO(un6_s_frac_rnd_0_cry_26));
  FDS desc2560(.Q(s_shr1[5:5]),.D(v_shr_2[5:5]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2561(.Q(s_shr1[4:4]),.D(v_shr_2[4:4]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2562(.Q(s_shr1[3:3]),.D(v_shr_2[3:3]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2563(.Q(s_shr1[2:2]),.D(v_shr_2[2:2]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2564(.Q(s_shr1[1:1]),.D(v_shr_2[1:1]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2565(.Q(s_shr1[0:0]),.D(v_shr_2[0:0]),.C(clk_i),.S(v_shr_2[6:6]));
  FDS desc2566(.Q(post_norm_div_output[31:31]),.D(s_sign_i),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2567(.Q(post_norm_div_output[30:30]),.D(s_output_o[30:30]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2568(.Q(post_norm_div_output[29:29]),.D(s_output_o[29:29]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2569(.Q(post_norm_div_output[28:28]),.D(s_output_o[28:28]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2570(.Q(post_norm_div_output[27:27]),.D(s_output_o[27:27]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2571(.Q(post_norm_div_output[26:26]),.D(s_output_o[26:26]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2572(.Q(post_norm_div_output[25:25]),.D(s_output_o[25:25]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2573(.Q(post_norm_div_output[24:24]),.D(s_output_o[24:24]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2574(.Q(post_norm_div_output[23:23]),.D(s_output_o[23:23]),.C(clk_i),.S(un7_s_nan_in));
  FDS desc2575(.Q(post_norm_div_output[22:22]),.D(s_output_o[22:22]),.C(clk_i),.S(un7_s_nan_in));
  VCC VCC_cZ(.P(VCC));
  GND GND_cZ(.G(GND));
  LUT2 un6_s_frac_rnd_1_s_26_RNI6NIC_o6(.I0(N_271),.I1(s_roundup),.O(N_27));
defparam un6_s_frac_rnd_1_s_26_RNI6NIC_o6.INIT=4'hB;
  LUT4 un6_s_frac_rnd_1_s_26_RNI6NIC_o5(.I0(s_expo1[0:0]),.I1(s_fraco1[26:26]),.I2(s_expo3_31[0:0]),.I3(s_roundup),.O(s_expo3_3[0:0]));
defparam un6_s_frac_rnd_1_s_26_RNI6NIC_o5.INIT=16'hF099;
  LUT4 desc2576(.I0(s_infb),.I1(un1_s_infa),.I2(result_4),.I3(un6_s_inf_result),.O(s_expo3_RNISDPK1_O6[5:5]));
defparam desc2576.INIT=16'hFFEF;
  LUT5 desc2577(.I0(s_expo3[5:5]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.O(s_output_o[28:28]));
defparam desc2577.INIT=32'hFFFFFEFC;
  LUT2 un2_s_lost_0_ac0_1_lut6_2_o6(.I0(s_shr1[0:0]),.I1(s_shr1[1:1]),.O(un2_s_lost_0_c2));
defparam un2_s_lost_0_ac0_1_lut6_2_o6.INIT=4'h8;
  LUT5 un2_s_lost_0_ac0_1_lut6_2_o5(.I0(s_qutnt_i[26:26]),.I1(s_shr1[0:0]),.I2(s_shr1[1:1]),.I3(s_shr1[3:3]),.I4(s_shr1[2:2]),.O(N_108));
defparam un2_s_lost_0_ac0_1_lut6_2_o5.INIT=32'h00000002;
  LUT2 desc2578(.I0(s_qutnt_i[24:24]),.I1(s_qutnt_i[25:25]),.O(N_114));
defparam desc2578.INIT=4'h1;
  LUT4 desc2579(.I0(s_qutnt_i[25:25]),.I1(s_shl1),.I2(N_108),.I3(un1_s_shr1_1),.O(s_fraco1_3[26:26]));
defparam desc2579.INIT=16'hB800;
  LUT2 desc2580(.I0(s_qutnt_i[1:1]),.I1(s_qutnt_i[3:3]),.O(N_1423));
defparam desc2580.INIT=4'hE;
  LUT4 desc2581(.I0(s_qutnt_i[0:0]),.I1(s_qutnt_i[1:1]),.I2(s_qutnt_i[2:2]),.I3(s_qutnt_i[3:3]),.O(N_1433));
defparam desc2581.INIT=16'hFFFE;
  LUT2 desc2582(.I0(s_qutnt_i[6:6]),.I1(s_qutnt_i[7:7]),.O(N_1422));
defparam desc2582.INIT=4'hE;
  LUT4 desc2583(.I0(s_qutnt_i[6:6]),.I1(s_qutnt_i[7:7]),.I2(s_qutnt_i[4:4]),.I3(s_qutnt_i[5:5]),.O(N_1480));
defparam desc2583.INIT=16'h0001;
  LUT2 desc2584(.I0(s_qutnt_i[14:14]),.I1(s_qutnt_i[15:15]),.O(N_1419));
defparam desc2584.INIT=4'hE;
  LUT4 desc2585(.I0(s_qutnt_i[14:14]),.I1(s_qutnt_i[15:15]),.I2(s_qutnt_i[12:12]),.I3(s_qutnt_i[13:13]),.O(N_1426));
defparam desc2585.INIT=16'hFFFE;
  LUT3 un1_s_infa_0_lut6_2_o6(.I0(s_opa_i[23:23]),.I1(s_opa_i_1),.I2(s_opa_i_2),.O(un1_s_infa_0));
defparam un1_s_infa_0_lut6_2_o6.INIT=8'h80;
  LUT4 un1_s_infa_0_lut6_2_o5(.I0(s_opa_i_1),.I1(s_opa_i_2),.I2(s_opa_i_3),.I3(s_opa_i_4),.O(result_4_0_3));
defparam un1_s_infa_0_lut6_2_o5.INIT=16'hFFFE;
  LUT3 s_exp_10b_axbxc1_lut6_2_o6(.I0(s_exp_10_i[1:1]),.I1(s_exp_10_i[0:0]),.I2(s_qutnt_i[26:26]),.O(s_exp_10b[1:1]));
defparam s_exp_10b_axbxc1_lut6_2_o6.INIT=8'hA9;
  LUT3 s_exp_10b_axbxc1_lut6_2_o5(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[2:2]));
defparam s_exp_10b_axbxc1_lut6_2_o5.INIT=8'h06;
  LUT5 desc2586(.I0(s_qutnt_i[24:24]),.I1(s_qutnt_i[25:25]),.I2(s_qutnt_i[26:26]),.I3(s_shr1[0:0]),.I4(s_shr1[1:1]),.O(N_52));
defparam desc2586.INIT=32'h00F0CCAA;
  LUT3 desc2587(.I0(s_qutnt_i[26:26]),.I1(s_shr1[0:0]),.I2(s_shr1[1:1]),.O(N_54));
defparam desc2587.INIT=8'h02;
  LUT4 desc2588(.I0(s_qutnt_i[23:23]),.I1(s_qutnt_i[24:24]),.I2(s_qutnt_i[25:25]),.I3(s_qutnt_i[26:26]),.O(N_123));
defparam desc2588.INIT=16'h4544;
  LUT2 desc2589(.I0(s_qutnt_i[23:23]),.I1(s_qutnt_i[22:22]),.O(N_1424));
defparam desc2589.INIT=4'hE;
  LUT3 desc2590(.I0(s_shr1[2:2]),.I1(N_33),.I2(N_37),.O(N_60));
defparam desc2590.INIT=8'hE4;
  LUT3 desc2591(.I0(s_shr1[2:2]),.I1(N_41),.I2(N_45),.O(N_68));
defparam desc2591.INIT=8'hE4;
  LUT2 un6_s_infa_lut6_2_o6(.I0(s_infb),.I1(un1_s_infa),.O(un6_s_infa));
defparam un6_s_infa_lut6_2_o6.INIT=4'hE;
  LUT5 un6_s_infa_lut6_2_o5(.I0(s_expo3[0:0]),.I1(s_infb),.I2(un1_s_infa),.I3(result_4),.I4(un6_s_inf_result),.O(s_output_o[23:23]));
defparam un6_s_infa_lut6_2_o5.INIT=32'hFFFFFEFC;
  LUT3 desc2592(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_52),.O(N_106));
defparam desc2592.INIT=8'h10;
  LUT5 desc2593(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_52),.I4(N_90),.O(N_117));
defparam desc2593.INIT=32'h57550200;
  LUT3 desc2594(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_51),.O(N_105));
defparam desc2594.INIT=8'h10;
  LUT5 desc2595(.I0(s_shr1[4:4]),.I1(s_shr1[3:3]),.I2(s_shr1[2:2]),.I3(N_51),.I4(N_89),.O(N_116));
defparam desc2595.INIT=32'h57550200;
  LUT5 desc2596(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_52),.I3(N_44),.I4(N_48),.O(N_98));
defparam desc2596.INIT=32'h75643120;
  LUT4 desc2597(.I0(s_shr1[3:3]),.I1(s_shr1[2:2]),.I2(N_52),.I3(N_48),.O(N_102));
defparam desc2597.INIT=16'h5140;
  LUT5 s_exp_10b_axbxc3_lut6_2_o6(.I0(s_exp_10_i[3:3]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10_i[0:0]),.I4(s_qutnt_i[26:26]),.O(s_exp_10b[3:3]));
defparam s_exp_10b_axbxc3_lut6_2_o6.INIT=32'hAAAAAAA9;
  LUT4 s_exp_10b_axbxc3_lut6_2_o5(.I0(s_exp_10_i[2:2]),.I1(s_exp_10_i[1:1]),.I2(s_exp_10_i[0:0]),.I3(s_qutnt_i[26:26]),.O(s_exp_10b[2:2]));
defparam s_exp_10b_axbxc3_lut6_2_o5.INIT=16'hAAA9;
  LUT3 desc2598(.I0(s_shr1[4:4]),.I1(N_107),.I2(N_91),.O(N_118));
defparam desc2598.INIT=8'hD8;
  LUT3 desc2599(.I0(s_shr1[4:4]),.I1(N_82),.I2(N_98),.O(N_109));
defparam desc2599.INIT=8'hE4;
  LUT3 desc2600(.I0(s_shr1[4:4]),.I1(N_83),.I2(N_99),.O(N_110));
defparam desc2600.INIT=8'hE4;
  LUT3 desc2601(.I0(s_shr1[4:4]),.I1(N_84),.I2(N_100),.O(N_111));
defparam desc2601.INIT=8'hE4;
  LUT5 un18_s_roundup_lut6_2_o6(.I0(s_fraco1[0:0]),.I1(s_fraco1[1:1]),.I2(s_fraco1[2:2]),.I3(result_3_2_4),.I4(result_3_3_4),.O(un18_s_roundup));
defparam un18_s_roundup_lut6_2_o6.INIT=32'hFFFFFFFE;
  LUT5 un18_s_roundup_lut6_2_o5(.I0(s_fraco1[0:0]),.I1(s_fraco1[1:1]),.I2(s_fraco1[2:2]),.I3(result_3_2_4),.I4(result_3_3_4),.O(un4_s_ine_o_1));
defparam un18_s_roundup_lut6_2_o5.INIT=32'hFFFFFFFE;
  LUT3 desc2602(.I0(s_fraco1[6:6]),.I1(un6_s_frac_rnd1[3:3]),.I2(s_roundup),.O(s_frac_rnd[3:3]));
defparam desc2602.INIT=8'hCA;
  LUT3 desc2603(.I0(s_fraco1[7:7]),.I1(un6_s_frac_rnd1[4:4]),.I2(s_roundup),.O(s_frac_rnd[4:4]));
defparam desc2603.INIT=8'hCA;
  LUT3 desc2604(.I0(s_fraco1[25:25]),.I1(un6_s_frac_rnd1[22:22]),.I2(s_roundup),.O(s_frac_rnd[22:22]));
defparam desc2604.INIT=8'hCA;
  LUT3 desc2605(.I0(s_fraco1[24:24]),.I1(un6_s_frac_rnd1[21:21]),.I2(s_roundup),.O(s_frac_rnd[21:21]));
defparam desc2605.INIT=8'hCA;
  LUT3 desc2606(.I0(s_fraco1[10:10]),.I1(un6_s_frac_rnd1[7:7]),.I2(s_roundup),.O(s_frac_rnd[7:7]));
defparam desc2606.INIT=8'hCA;
  LUT3 desc2607(.I0(s_fraco1[9:9]),.I1(un6_s_frac_rnd1[6:6]),.I2(s_roundup),.O(s_frac_rnd[6:6]));
defparam desc2607.INIT=8'hCA;
  LUT3 desc2608(.I0(s_fraco1[12:12]),.I1(un6_s_frac_rnd1[9:9]),.I2(s_roundup),.O(s_frac_rnd[9:9]));
defparam desc2608.INIT=8'hCA;
  LUT3 desc2609(.I0(s_fraco1[11:11]),.I1(un6_s_frac_rnd1[8:8]),.I2(s_roundup),.O(s_frac_rnd[8:8]));
defparam desc2609.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_27_RNIJUFE_o6(.I0(s_expo3_30[1:1]),.I1(s_expo3_31[1:1]),.I2(s_roundup),.O(s_expo3_3[1:1]));
defparam un6_s_frac_rnd_1_s_27_RNIJUFE_o6.INIT=8'hCA;
  LUT2 un6_s_frac_rnd_1_s_27_RNIJUFE_o5(.I0(s_fraco1[3:3]),.I1(s_roundup),.O(s_frac_rnd[0:0]));
defparam un6_s_frac_rnd_1_s_27_RNIJUFE_o5.INIT=4'h6;
  LUT3 desc2610(.I0(s_fraco1[23:23]),.I1(un6_s_frac_rnd1[20:20]),.I2(s_roundup),.O(s_frac_rnd[20:20]));
defparam desc2610.INIT=8'hCA;
  LUT3 desc2611(.I0(s_fraco1[22:22]),.I1(un6_s_frac_rnd1[19:19]),.I2(s_roundup),.O(s_frac_rnd[19:19]));
defparam desc2611.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_28_RNIUSMJ_o6(.I0(s_expo3_30[3:3]),.I1(s_expo3_31[3:3]),.I2(s_roundup),.O(s_expo3_3[3:3]));
defparam un6_s_frac_rnd_1_s_28_RNIUSMJ_o6.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_28_RNIUSMJ_o5(.I0(s_expo3_30[2:2]),.I1(s_expo3_31[2:2]),.I2(s_roundup),.O(s_expo3_3[2:2]));
defparam un6_s_frac_rnd_1_s_28_RNIUSMJ_o5.INIT=8'hCA;
  LUT3 desc2612(.I0(s_fraco1[20:20]),.I1(un6_s_frac_rnd1[17:17]),.I2(s_roundup),.O(s_frac_rnd[17:17]));
defparam desc2612.INIT=8'hCA;
  LUT3 desc2613(.I0(s_fraco1[19:19]),.I1(un6_s_frac_rnd1[16:16]),.I2(s_roundup),.O(s_frac_rnd[16:16]));
defparam desc2613.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_30_RNI20NJ_o6(.I0(s_expo3_30[5:5]),.I1(s_expo3_31[5:5]),.I2(s_roundup),.O(s_expo3_3[5:5]));
defparam un6_s_frac_rnd_1_s_30_RNI20NJ_o6.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_30_RNI20NJ_o5(.I0(s_expo3_30[4:4]),.I1(s_expo3_31[4:4]),.I2(s_roundup),.O(s_expo3_3[4:4]));
defparam un6_s_frac_rnd_1_s_30_RNI20NJ_o5.INIT=8'hCA;
  LUT3 desc2614(.I0(s_fraco1[18:18]),.I1(un6_s_frac_rnd1[15:15]),.I2(s_roundup),.O(s_frac_rnd[15:15]));
defparam desc2614.INIT=8'hCA;
  LUT3 desc2615(.I0(s_fraco1[17:17]),.I1(un6_s_frac_rnd1[14:14]),.I2(s_roundup),.O(s_frac_rnd[14:14]));
defparam desc2615.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_32_RNIA0NJ_o6(.I0(s_expo3_30[7:7]),.I1(s_expo3_31[7:7]),.I2(s_roundup),.O(s_expo3_3[7:7]));
defparam un6_s_frac_rnd_1_s_32_RNIA0NJ_o6.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_32_RNIA0NJ_o5(.I0(s_expo3_30[6:6]),.I1(s_expo3_31[6:6]),.I2(s_roundup),.O(s_expo3_3[6:6]));
defparam un6_s_frac_rnd_1_s_32_RNIA0NJ_o5.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_34_RNICTOL_o6(.I0(s_expo3_30[8:8]),.I1(s_expo3_31[8:8]),.I2(s_roundup),.O(s_expo3_3[8:8]));
defparam un6_s_frac_rnd_1_s_34_RNICTOL_o6.INIT=8'hCA;
  LUT3 un6_s_frac_rnd_1_s_34_RNICTOL_o5(.I0(s_fraco1[8:8]),.I1(un6_s_frac_rnd1[5:5]),.I2(s_roundup),.O(s_frac_rnd[5:5]));
defparam un6_s_frac_rnd_1_s_34_RNICTOL_o5.INIT=8'hCA;
  LUT3 desc2616(.I0(s_fraco1[5:5]),.I1(un6_s_frac_rnd1[2:2]),.I2(s_roundup),.O(s_frac_rnd[2:2]));
defparam desc2616.INIT=8'hCA;
  LUT3 desc2617(.I0(s_fraco1[4:4]),.I1(un6_s_frac_rnd1[1:1]),.I2(s_roundup),.O(s_frac_rnd[1:1]));
defparam desc2617.INIT=8'hCA;
  LUT3 desc2618(.I0(s_fraco1[13:13]),.I1(un6_s_frac_rnd1[10:10]),.I2(s_roundup),.O(s_frac_rnd[10:10]));
defparam desc2618.INIT=8'hCA;
  LUT3 desc2619(.I0(s_fraco1[14:14]),.I1(un6_s_frac_rnd1[11:11]),.I2(s_roundup),.O(s_frac_rnd[11:11]));
defparam desc2619.INIT=8'hCA;
  LUT3 desc2620(.I0(s_fraco1[15:15]),.I1(un6_s_frac_rnd1[12:12]),.I2(s_roundup),.O(s_frac_rnd[12:12]));
defparam desc2620.INIT=8'hCA;
  LUT3 desc2621(.I0(s_fraco1[16:16]),.I1(un6_s_frac_rnd1[13:13]),.I2(s_roundup),.O(s_frac_rnd[13:13]));
defparam desc2621.INIT=8'hCA;
  LUT4 s_exp_10b_axbxc7_lut6_2_o6(.I0(s_exp_10_i[7:7]),.I1(s_exp_10_i[6:6]),.I2(s_exp_10_i[5:5]),.I3(s_exp_10b_c5),.O(s_exp_10b[7:7]));
defparam s_exp_10b_axbxc7_lut6_2_o6.INIT=16'hAAA9;
  LUT2 s_exp_10b_axbxc7_lut6_2_o5(.I0(s_exp_10_i[5:5]),.I1(s_exp_10b_c5),.O(s_exp_10b[5:5]));
defparam s_exp_10b_axbxc7_lut6_2_o5.INIT=4'h9;
  LUT3 v_shr_1_c4_RNIPTMG5_o6(.I0(v_shr_1_c4),.I1(s_exp_10b[4:4]),.I2(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[4:4]));
defparam v_shr_1_c4_RNIPTMG5_o6.INIT=8'h06;
  LUT5 v_shr_1_c4_RNIPTMG5_o5(.I0(s_exp_10_i[5:5]),.I1(v_shr_1_c4),.I2(s_exp_10b[4:4]),.I3(s_exp_10b_c5),.I4(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[5:5]));
defparam v_shr_1_c4_RNIPTMG5_o5.INIT=32'h000056A9;
  LUT2 desc2622(.I0(s_exp_10_i[1:1]),.I1(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[1:1]));
defparam desc2622.INIT=4'h2;
  LUT4 desc2623(.I0(s_exp_10_i[3:3]),.I1(s_exp_10_i[2:2]),.I2(s_exp_10_i[1:1]),.I3(s_exp_10b_axbxc8_RNIGLJC4),.O(v_shr_2[3:3]));
defparam desc2623.INIT=16'h0056;
endmodule
module pre_norm_sqrt_inj (v_count,v_count_i,v_count_1_0_a2_7_i_0,v_count_56_0_2,pre_norm_sqrt_fracta_o_0,s_fracta_52_o_0_e,pre_norm_div_dvdnd_0,pre_norm_sqrt_exp_o,v_count_1_0_0_a2_0,v_count_1_0_1,v_count_1_0_2,pre_norm_div_dvdnd_17,pre_norm_div_dvdnd_16,pre_norm_div_dvdnd_9,pre_norm_div_dvdnd_10,pre_norm_div_dvdnd_11,pre_norm_div_dvdnd_8,pre_norm_div_dvdnd_21,pre_norm_div_dvdnd_22,pre_norm_div_dvdnd_18,pre_norm_div_dvdnd_20,pre_norm_div_dvdnd_19,s_opa_i_23,s_opa_i_0,s_opa_i_2,s_opa_i_3,s_opa_i_1,s_opa_i_8,s_opa_i_10,s_opa_i_11,s_opa_i_9,s_opa_i_6,s_opa_i_7,s_opa_i_5,s_opa_i_4,s_opa_i_14,s_opa_i_12,s_opa_i_13,s_opa_i_15,s_opa_i_21,s_opa_i_22,s_opa_i_20,s_opa_i_24,s_opa_i_30,s_opa_i_27,s_opa_i_25,s_opa_i_26,pre_norm_sqrt_fracta_o_15,pre_norm_sqrt_fracta_o_16,pre_norm_sqrt_fracta_o_6,pre_norm_sqrt_fracta_o_10,pre_norm_sqrt_fracta_o_9,pre_norm_sqrt_fracta_o_8,pre_norm_sqrt_fracta_o_7,pre_norm_sqrt_fracta_o_21,pre_norm_sqrt_fracta_o_0_d0,pre_norm_sqrt_fracta_o_18,pre_norm_sqrt_fracta_o_19,pre_norm_sqrt_fracta_o_22,pre_norm_sqrt_fracta_o_11,pre_norm_sqrt_fracta_o_12,pre_norm_sqrt_fracta_o_13,pre_norm_sqrt_fracta_o_14,pre_norm_sqrt_fracta_o_20,s_opa_i_i,N_88,N_55,s_dvdnd_50_o_108_0_e,N_38_0,N_1620,s_dvdnd_50_o_105_0_e,N_45,N_1619,N_41,N_1624,N_1087,N_1166,N_1174,un2_s_snan_o_8,N_95,N_1245,N_53,N_48_0,s_dvdnd_50_o_106_0_e,m49_0_e,s_dvdnd_50_o_102_0_e,s_dvdnd_50_o_109_0_e,N_1238,N_1227,clk_i,un2_s_snan_o_20,N_1077,N_399,N_396,N_44,N_1241,N_30_0,un2_s_snan_o_22,result_i_o3_lut6_2_O6,N_1242,N_27_0,N_63,N_1264);
inout [4:1] v_count ;
input v_count_i ;
output v_count_1_0_a2_7_i_0 ;
output [4:4] v_count_56_0_2 ;
output [51:51] pre_norm_sqrt_fracta_o_0 ;
output [33:30] s_fracta_52_o_0_e ;
output [49:49] pre_norm_div_dvdnd_0 ;
output [7:0] pre_norm_sqrt_exp_o ;
input [1:1] v_count_1_0_0_a2_0 ;
input v_count_1_0_1 ;
input v_count_1_0_2 ;
input pre_norm_div_dvdnd_17 ;
output pre_norm_div_dvdnd_16 ;
input pre_norm_div_dvdnd_9 ;
input pre_norm_div_dvdnd_10 ;
output pre_norm_div_dvdnd_11 ;
output pre_norm_div_dvdnd_8 ;
input pre_norm_div_dvdnd_21 ;
output pre_norm_div_dvdnd_22 ;
input pre_norm_div_dvdnd_18 ;
output pre_norm_div_dvdnd_20 ;
output pre_norm_div_dvdnd_19 ;
input s_opa_i_23 ;
input s_opa_i_0 ;
input s_opa_i_2 ;
input s_opa_i_3 ;
input s_opa_i_1 ;
input s_opa_i_8 ;
input s_opa_i_10 ;
input s_opa_i_11 ;
input s_opa_i_9 ;
input s_opa_i_6 ;
input s_opa_i_7 ;
input s_opa_i_5 ;
input s_opa_i_4 ;
input s_opa_i_14 ;
input s_opa_i_12 ;
input s_opa_i_13 ;
input s_opa_i_15 ;
input s_opa_i_21 ;
input s_opa_i_22 ;
input s_opa_i_20 ;
input s_opa_i_24 ;
input s_opa_i_30 ;
input s_opa_i_27 ;
input s_opa_i_25 ;
input s_opa_i_26 ;
output pre_norm_sqrt_fracta_o_15 ;
output pre_norm_sqrt_fracta_o_16 ;
output pre_norm_sqrt_fracta_o_6 ;
output pre_norm_sqrt_fracta_o_10 ;
output pre_norm_sqrt_fracta_o_9 ;
output pre_norm_sqrt_fracta_o_8 ;
output pre_norm_sqrt_fracta_o_7 ;
output pre_norm_sqrt_fracta_o_21 ;
output pre_norm_sqrt_fracta_o_0_d0 ;
output pre_norm_sqrt_fracta_o_18 ;
output pre_norm_sqrt_fracta_o_19 ;
output pre_norm_sqrt_fracta_o_22 ;
output pre_norm_sqrt_fracta_o_11 ;
output pre_norm_sqrt_fracta_o_12 ;
output pre_norm_sqrt_fracta_o_13 ;
output pre_norm_sqrt_fracta_o_14 ;
output pre_norm_sqrt_fracta_o_20 ;
input [29:28] s_opa_i_i ;
output N_88 ;
input N_55 ;
output s_dvdnd_50_o_108_0_e ;
input N_38_0 ;
input N_1620 ;
output s_dvdnd_50_o_105_0_e ;
input N_45 ;
input N_1619 ;
input N_41 ;
input N_1624 ;
output N_1087 ;
output N_1166 ;
output N_1174 ;
output un2_s_snan_o_8 ;
input N_95 ;
input N_1245 ;
output N_53 ;
input N_48_0 ;
output s_dvdnd_50_o_106_0_e ;
output m49_0_e ;
output s_dvdnd_50_o_102_0_e ;
output s_dvdnd_50_o_109_0_e ;
input N_1238 ;
input N_1227 ;
input clk_i ;
input un2_s_snan_o_20 ;
input N_1077 ;
input N_399 ;
input N_396 ;
input N_44 ;
input N_1241 ;
input N_30_0 ;
input un2_s_snan_o_22 ;
input result_i_o3_lut6_2_O6 ;
input N_1242 ;
input N_27_0 ;
input N_63 ;
input N_1264 ;
wire pre_norm_div_dvdnd_17 ;
wire pre_norm_div_dvdnd_16 ;
wire pre_norm_div_dvdnd_9 ;
wire pre_norm_div_dvdnd_10 ;
wire pre_norm_div_dvdnd_11 ;
wire pre_norm_div_dvdnd_8 ;
wire pre_norm_div_dvdnd_21 ;
wire pre_norm_div_dvdnd_22 ;
wire pre_norm_div_dvdnd_18 ;
wire pre_norm_div_dvdnd_20 ;
wire pre_norm_div_dvdnd_19 ;
wire s_opa_i_23 ;
wire s_opa_i_0 ;
wire s_opa_i_2 ;
wire s_opa_i_3 ;
wire s_opa_i_1 ;
wire s_opa_i_8 ;
wire s_opa_i_10 ;
wire s_opa_i_11 ;
wire s_opa_i_9 ;
wire s_opa_i_6 ;
wire s_opa_i_7 ;
wire s_opa_i_5 ;
wire s_opa_i_4 ;
wire s_opa_i_14 ;
wire s_opa_i_12 ;
wire s_opa_i_13 ;
wire s_opa_i_15 ;
wire s_opa_i_21 ;
wire s_opa_i_22 ;
wire s_opa_i_20 ;
wire s_opa_i_24 ;
wire s_opa_i_30 ;
wire s_opa_i_27 ;
wire s_opa_i_25 ;
wire s_opa_i_26 ;
wire pre_norm_sqrt_fracta_o_15 ;
wire pre_norm_sqrt_fracta_o_16 ;
wire pre_norm_sqrt_fracta_o_6 ;
wire pre_norm_sqrt_fracta_o_10 ;
wire pre_norm_sqrt_fracta_o_9 ;
wire pre_norm_sqrt_fracta_o_8 ;
wire pre_norm_sqrt_fracta_o_7 ;
wire pre_norm_sqrt_fracta_o_21 ;
wire pre_norm_sqrt_fracta_o_0_d0 ;
wire pre_norm_sqrt_fracta_o_18 ;
wire pre_norm_sqrt_fracta_o_19 ;
wire pre_norm_sqrt_fracta_o_22 ;
wire pre_norm_sqrt_fracta_o_11 ;
wire pre_norm_sqrt_fracta_o_12 ;
wire pre_norm_sqrt_fracta_o_13 ;
wire pre_norm_sqrt_fracta_o_14 ;
wire pre_norm_sqrt_fracta_o_20 ;
wire N_88 ;
wire N_55 ;
wire s_dvdnd_50_o_108_0_e ;
wire N_38_0 ;
wire N_1620 ;
wire s_dvdnd_50_o_105_0_e ;
wire N_45 ;
wire N_1619 ;
wire N_41 ;
wire N_1624 ;
wire N_1087 ;
wire N_1166 ;
wire N_1174 ;
wire un2_s_snan_o_8 ;
wire N_95 ;
wire N_1245 ;
wire N_53 ;
wire N_48_0 ;
wire s_dvdnd_50_o_106_0_e ;
wire m49_0_e ;
wire s_dvdnd_50_o_102_0_e ;
wire s_dvdnd_50_o_109_0_e ;
wire N_1238 ;
wire N_1227 ;
wire clk_i ;
wire un2_s_snan_o_20 ;
wire N_1077 ;
wire N_399 ;
wire N_396 ;
wire N_44 ;
wire N_1241 ;
wire N_30_0 ;
wire un2_s_snan_o_22 ;
wire result_i_o3_lut6_2_O6 ;
wire N_1242 ;
wire N_27_0 ;
wire N_63 ;
wire N_1264 ;
wire [49:26] pre_norm_div_dvdnd ;
wire [4:4] v_count_0_o3_i_o2_0 ;
wire [8:8] s_exp_tem_1 ;
wire [8:1] s_exp_tem ;
wire [49:49] pre_norm_div_dvdnd_i ;
wire [8:8] s_exp_tem_0 ;
wire [2:2] v_count_0_a2_1 ;
wire GND ;
wire VCC ;
wire N_73 ;
wire N_57 ;
wire N_69 ;
wire N_208 ;
wire s_exp_tem_axb_1 ;
wire s_exp_tem_axb_0 ;
wire N_92 ;
wire s_exp_tem_axb_7 ;
wire s_exp_tem_axb_4 ;
wire s_exp_tem_axb_2 ;
wire s_exp_tem_axb_3 ;
wire s_exp_tem_cry_6 ;
wire s_exp_tem_cry_5 ;
wire s_exp_tem_cry_4 ;
wire s_exp_tem_cry_3 ;
wire s_exp_tem_cry_2 ;
wire s_exp_tem_cry_1 ;
wire s_exp_tem_cry_0 ;
// instances
  LUT6_2 desc2624(.I0(s_opa_i_0),.I1(v_count[1:1]),.I2(v_count[3:3]),.I3(v_count[2:2]),.I4(v_count_i),.I5(v_count[4:4]),.O6(pre_norm_div_dvdnd[26:26]),.O5(N_73));
defparam desc2624.INIT=64'h0000000000020000;
  LUT5 desc2625(.I0(N_48_0),.I1(N_1620),.I2(v_count[3:3]),.I3(s_opa_i_23),.I4(v_count[4:4]),.O(s_fracta_52_o_0_e[30:30]));
defparam desc2625.INIT=32'h00000C0A;
  LUT6 desc2626(.I0(v_count[1:1]),.I1(v_count[2:2]),.I2(v_count[3:3]),.I3(v_count_i),.I4(s_opa_i_0),.I5(v_count[4:4]),.O(s_dvdnd_50_o_102_0_e));
defparam desc2626.INIT=64'h0000000001000000;
  LUT5 desc2627(.I0(N_38_0),.I1(N_1620),.I2(v_count[2:2]),.I3(v_count[3:3]),.I4(v_count[4:4]),.O(s_dvdnd_50_o_109_0_e));
defparam desc2627.INIT=32'h000000C5;
  LUT6 desc2628(.I0(N_1620),.I1(N_53),.I2(v_count[2:2]),.I3(v_count[3:3]),.I4(s_opa_i_23),.I5(v_count[4:4]),.O(s_fracta_52_o_0_e[31:31]));
defparam desc2628.INIT=64'h0000000000CC000A;
  LUT5 desc2629(.I0(N_1238),.I1(N_53),.I2(v_count[3:3]),.I3(s_opa_i_23),.I4(v_count[4:4]),.O(s_fracta_52_o_0_e[32:32]));
defparam desc2629.INIT=32'h00000A0C;
  LUT5 desc2630(.I0(N_1238),.I1(N_55),.I2(v_count[3:3]),.I3(s_opa_i_23),.I4(v_count[4:4]),.O(s_fracta_52_o_0_e[33:33]));
defparam desc2630.INIT=32'h00000C0A;
  LUT6 desc2631(.I0(N_1166),.I1(N_1174),.I2(N_1227),.I3(s_opa_i_4),.I4(s_opa_i_5),.I5(un2_s_snan_o_8),.O(pre_norm_div_dvdnd_0[49:49]));
defparam desc2631.INIT=64'hFFFFFFEFFFFFFFFF;
  LUT1 s_exp_tem_cry_7_outextlut(.I0(GND),.O(s_exp_tem_1[8:8]));
defparam s_exp_tem_cry_7_outextlut.INIT=2'h3;
  FD desc2632(.Q(pre_norm_sqrt_exp_o[2:2]),.D(s_exp_tem[3:3]),.C(clk_i));
  FD desc2633(.Q(pre_norm_sqrt_exp_o[3:3]),.D(s_exp_tem[4:4]),.C(clk_i));
  FD desc2634(.Q(pre_norm_sqrt_exp_o[6:6]),.D(s_exp_tem[7:7]),.C(clk_i));
  FD desc2635(.Q(pre_norm_sqrt_exp_o[7:7]),.D(s_exp_tem[8:8]),.C(clk_i));
  FDR desc2636(.Q(pre_norm_sqrt_exp_o[0:0]),.D(s_exp_tem[1:1]),.C(clk_i),.R(pre_norm_div_dvdnd_i[49:49]));
  FDR desc2637(.Q(pre_norm_sqrt_exp_o[1:1]),.D(s_exp_tem[2:2]),.C(clk_i),.R(pre_norm_div_dvdnd_i[49:49]));
  FDR desc2638(.Q(pre_norm_sqrt_exp_o[4:4]),.D(s_exp_tem[5:5]),.C(clk_i),.R(pre_norm_div_dvdnd_i[49:49]));
  FDR desc2639(.Q(pre_norm_sqrt_exp_o[5:5]),.D(s_exp_tem[6:6]),.C(clk_i),.R(pre_norm_div_dvdnd_i[49:49]));
  MUXCY s_exp_tem_cry_7_outext(.DI(GND),.CI(s_exp_tem_0[8:8]),.S(s_exp_tem_1[8:8]),.O(s_exp_tem[8:8]));
  LUT6 desc2640(.I0(s_opa_i_14),.I1(s_opa_i_12),.I2(s_opa_i_13),.I3(s_opa_i_15),.I4(un2_s_snan_o_20),.I5(N_208),.O(v_count_0_a2_1[2:2]));
defparam desc2640.INIT=64'h0001000100000001;
  LUT6_L s_exp_tem_axb_1_cZ(.I0(s_opa_i_21),.I1(s_opa_i_22),.I2(s_opa_i_20),.I3(s_opa_i_24),.I4(N_1077),.I5(v_count_1_0_0_a2_0[1:1]),.LO(s_exp_tem_axb_1));
defparam s_exp_tem_axb_1_cZ.INIT=64'h00FF00CC00FF00CD;
  LUT6 desc2641(.I0(s_opa_i_21),.I1(s_opa_i_22),.I2(s_opa_i_20),.I3(s_opa_i_24),.I4(N_1077),.I5(v_count_1_0_0_a2_0[1:1]),.O(v_count[1:1]));
defparam desc2641.INIT=64'h0000003300000032;
  LUT5 s_exp_tem_axb_0_cZ(.I0(s_opa_i_23),.I1(N_399),.I2(v_count_1_0_1),.I3(N_396),.I4(v_count_1_0_2),.O(s_exp_tem_axb_0));
defparam s_exp_tem_axb_0_cZ.INIT=32'hAAAAAAA9;
  LUT6 desc2642(.I0(N_1227),.I1(v_count[2:2]),.I2(N_44),.I3(N_1241),.I4(N_30_0),.I5(N_38_0),.O(N_92));
defparam desc2642.INIT=64'h1054327698DCBAFE;
  LUT6_L desc2643(.I0(s_opa_i_23),.I1(v_count[4:4]),.I2(v_count[2:2]),.I3(N_1620),.I4(N_92),.I5(pre_norm_div_dvdnd_18),.LO(pre_norm_sqrt_fracta_o_18));
defparam desc2643.INIT=64'h7F775D552A220800;
  LUT6_L desc2644(.I0(s_opa_i_23),.I1(v_count[4:4]),.I2(v_count[2:2]),.I3(N_1620),.I4(N_92),.I5(pre_norm_div_dvdnd_20),.LO(pre_norm_sqrt_fracta_o_19));
defparam desc2644.INIT=64'hBFBBAEAA15110400;
  LUT4_L desc2645(.I0(v_count[4:4]),.I1(v_count[2:2]),.I2(N_1620),.I3(N_92),.LO(pre_norm_div_dvdnd_19));
defparam desc2645.INIT=16'h7520;
  LUT5_L desc2646(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd[49:49]),.I2(v_count[4:4]),.I3(N_55),.I4(N_95),.LO(pre_norm_sqrt_fracta_o_22));
defparam desc2646.INIT=32'hDD8DD888;
  LUT1_L s_exp_tem_axb_7_cZ(.I0(s_opa_i_30),.LO(s_exp_tem_axb_7));
defparam s_exp_tem_axb_7_cZ.INIT=2'h2;
  LUT4_L desc2647(.I0(s_opa_i_14),.I1(s_opa_i_12),.I2(s_opa_i_13),.I3(s_opa_i_15),.LO(v_count_0_o3_i_o2_0[4:4]));
defparam desc2647.INIT=16'hFFFE;
  LUT5_L desc2648(.I0(s_opa_i_6),.I1(s_opa_i_7),.I2(s_opa_i_4),.I3(s_opa_i_5),.I4(N_1166),.LO(N_208));
defparam desc2648.INIT=32'h00010000;
  LUT6 desc2649(.I0(s_opa_i_21),.I1(s_opa_i_22),.I2(s_opa_i_20),.I3(un2_s_snan_o_22),.I4(v_count_0_a2_1[2:2]),.I5(result_i_o3_lut6_2_O6),.O(v_count[2:2]));
defparam desc2649.INIT=64'h0000000001010001;
  LUT2_L s_exp_tem_axb_4_cZ(.I0(s_opa_i_27),.I1(v_count[4:4]),.LO(s_exp_tem_axb_4));
defparam s_exp_tem_axb_4_cZ.INIT=4'h9;
  LUT2_L s_exp_tem_axb_2_cZ(.I0(s_opa_i_25),.I1(v_count[2:2]),.LO(s_exp_tem_axb_2));
defparam s_exp_tem_axb_2_cZ.INIT=4'h9;
  LUT6 desc2650(.I0(s_opa_i_4),.I1(s_opa_i_5),.I2(un2_s_snan_o_8),.I3(N_1166),.I4(N_1174),.I5(N_1227),.O(pre_norm_div_dvdnd[49:49]));
defparam desc2650.INIT=64'hFFFFFFEFFFFFFFFF;
  LUT6 desc2651(.I0(s_opa_i_4),.I1(s_opa_i_5),.I2(un2_s_snan_o_8),.I3(N_1166),.I4(N_1174),.I5(N_1227),.O(v_count[3:3]));
defparam desc2651.INIT=64'hFFFF001000000000;
  LUT2_L s_exp_tem_axb_3_cZ(.I0(s_opa_i_26),.I1(v_count[3:3]),.LO(s_exp_tem_axb_3));
defparam s_exp_tem_axb_3_cZ.INIT=4'h9;
  LUT6 desc2652(.I0(s_opa_i_4),.I1(s_opa_i_5),.I2(un2_s_snan_o_8),.I3(N_1166),.I4(N_1174),.I5(N_1227),.O(pre_norm_div_dvdnd_i[49:49]));
defparam desc2652.INIT=64'h0000001000000000;
  LUT5 desc2653(.I0(s_opa_i_0),.I1(v_count[1:1]),.I2(v_count[2:2]),.I3(v_count_i),.I4(N_1619),.O(N_53));
defparam desc2653.INIT=32'h2F0F2000;
  LUT6 desc2654(.I0(s_opa_i_0),.I1(v_count[1:1]),.I2(v_count[3:3]),.I3(v_count[2:2]),.I4(v_count_i),.I5(N_57),.O(pre_norm_div_dvdnd_8));
defparam desc2654.INIT=64'h0F2F0F0F00200000;
  LUT6 desc2655(.I0(v_count[3:3]),.I1(v_count[2:2]),.I2(N_1241),.I3(N_30_0),.I4(N_38_0),.I5(N_1620),.O(N_88));
defparam desc2655.INIT=64'h89CDABEF01452367;
  LUT6 desc2656(.I0(N_1174),.I1(N_1227),.I2(v_count[2:2]),.I3(N_30_0),.I4(N_38_0),.I5(N_1620),.O(pre_norm_div_dvdnd_11));
defparam desc2656.INIT=64'h080F787F00077077;
  LUT5_L desc2657(.I0(s_opa_i_23),.I1(v_count[3:3]),.I2(N_53),.I3(N_1242),.I4(pre_norm_div_dvdnd_11),.LO(pre_norm_sqrt_fracta_o_11));
defparam desc2657.INIT=32'hD5F780A2;
  LUT6_L desc2658(.I0(s_opa_i_23),.I1(v_count[3:3]),.I2(N_27_0),.I3(N_53),.I4(N_1242),.I5(N_1238),.LO(pre_norm_sqrt_fracta_o_12));
defparam desc2658.INIT=64'hCE8ADF9B46025713;
  LUT6_L desc2659(.I0(s_opa_i_23),.I1(v_count[3:3]),.I2(N_27_0),.I3(N_63),.I4(N_1238),.I5(N_55),.LO(pre_norm_sqrt_fracta_o_13));
defparam desc2659.INIT=64'hEFCDAB8967452301;
  LUT5 desc2660(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(N_69),.I3(N_53),.I4(N_1242),.O(pre_norm_div_dvdnd_20));
defparam desc2660.INIT=32'h54107632;
  LUT5 desc2661(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(N_73),.I3(N_1264),.I4(N_57),.O(pre_norm_div_dvdnd_16));
defparam desc2661.INIT=32'hE2F3C0D1;
  LUT5_L desc2662(.I0(s_opa_i_23),.I1(v_count[3:3]),.I2(N_63),.I3(N_55),.I4(N_88),.LO(pre_norm_sqrt_fracta_o_14));
defparam desc2662.INIT=32'hFEBA5410;
  LUT3_L desc2663(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd_21),.I2(pre_norm_div_dvdnd_20),.LO(pre_norm_sqrt_fracta_o_20));
defparam desc2663.INIT=8'hD8;
  XORCY s_exp_tem_s_7(.LI(s_exp_tem_axb_7),.CI(s_exp_tem_cry_6),.O(s_exp_tem[7:7]));
  MUXCY s_exp_tem_cry_7(.DI(GND),.CI(s_exp_tem_cry_6),.S(s_exp_tem_axb_7),.O(s_exp_tem_0[8:8]));
  XORCY s_exp_tem_s_6(.LI(s_opa_i_i[29:29]),.CI(s_exp_tem_cry_5),.O(s_exp_tem[6:6]));
  MUXCY_L s_exp_tem_cry_6_cZ(.DI(VCC),.CI(s_exp_tem_cry_5),.S(s_opa_i_i[29:29]),.LO(s_exp_tem_cry_6));
  XORCY s_exp_tem_s_5(.LI(s_opa_i_i[28:28]),.CI(s_exp_tem_cry_4),.O(s_exp_tem[5:5]));
  MUXCY_L s_exp_tem_cry_5_cZ(.DI(VCC),.CI(s_exp_tem_cry_4),.S(s_opa_i_i[28:28]),.LO(s_exp_tem_cry_5));
  XORCY s_exp_tem_s_4(.LI(s_exp_tem_axb_4),.CI(s_exp_tem_cry_3),.O(s_exp_tem[4:4]));
  MUXCY_L s_exp_tem_cry_4_cZ(.DI(s_opa_i_27),.CI(s_exp_tem_cry_3),.S(s_exp_tem_axb_4),.LO(s_exp_tem_cry_4));
  XORCY s_exp_tem_s_3(.LI(s_exp_tem_axb_3),.CI(s_exp_tem_cry_2),.O(s_exp_tem[3:3]));
  MUXCY_L s_exp_tem_cry_3_cZ(.DI(s_opa_i_26),.CI(s_exp_tem_cry_2),.S(s_exp_tem_axb_3),.LO(s_exp_tem_cry_3));
  XORCY s_exp_tem_s_2(.LI(s_exp_tem_axb_2),.CI(s_exp_tem_cry_1),.O(s_exp_tem[2:2]));
  MUXCY_L s_exp_tem_cry_2_cZ(.DI(s_opa_i_25),.CI(s_exp_tem_cry_1),.S(s_exp_tem_axb_2),.LO(s_exp_tem_cry_2));
  XORCY s_exp_tem_s_1(.LI(s_exp_tem_axb_1),.CI(s_exp_tem_cry_0),.O(s_exp_tem[1:1]));
  MUXCY_L s_exp_tem_cry_1_cZ(.DI(s_opa_i_24),.CI(s_exp_tem_cry_0),.S(s_exp_tem_axb_1),.LO(s_exp_tem_cry_1));
  MUXCY_L s_exp_tem_cry_0_cZ(.DI(s_opa_i_23),.CI(GND),.S(s_exp_tem_axb_0),.LO(s_exp_tem_cry_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT3 desc2664(.I0(N_53),.I1(v_count[3:3]),.I2(v_count[4:4]),.O(s_dvdnd_50_o_106_0_e));
defparam desc2664.INIT=8'h02;
  LUT3 desc2665(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(N_48_0),.O(m49_0_e));
defparam desc2665.INIT=8'h10;
  LUT3 desc2666(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd[26:26]),.I2(N_1245),.O(pre_norm_sqrt_fracta_o_0_d0));
defparam desc2666.INIT=8'hE4;
  LUT2 desc2667(.I0(pre_norm_div_dvdnd[49:49]),.I1(s_opa_i_23),.O(pre_norm_sqrt_fracta_o_0[51:51]));
defparam desc2667.INIT=4'h2;
  LUT5 desc2668(.I0(s_opa_i_23),.I1(v_count[4:4]),.I2(N_55),.I3(N_95),.I4(pre_norm_div_dvdnd_21),.O(pre_norm_sqrt_fracta_o_21));
defparam desc2668.INIT=32'hF7D5A280;
  LUT3 desc2669(.I0(v_count[4:4]),.I1(N_55),.I2(N_95),.O(pre_norm_div_dvdnd_22));
defparam desc2669.INIT=8'hD8;
  LUT2 desc2670(.I0(s_opa_i_6),.I1(s_opa_i_7),.O(un2_s_snan_o_8));
defparam desc2670.INIT=4'h1;
  LUT5 desc2671(.I0(s_opa_i_6),.I1(s_opa_i_7),.I2(s_opa_i_8),.I3(s_opa_i_9),.I4(s_opa_i_5),.O(v_count_56_0_2[4:4]));
defparam desc2671.INIT=32'h00000001;
  LUT5 desc2672(.I0(s_opa_i_8),.I1(s_opa_i_10),.I2(s_opa_i_11),.I3(s_opa_i_9),.I4(v_count_0_o3_i_o2_0[4:4]),.O(N_1174));
defparam desc2672.INIT=32'hFFFFFFFE;
  LUT3 desc2673(.I0(s_opa_i_10),.I1(s_opa_i_11),.I2(s_opa_i_9),.O(v_count_1_0_a2_7_i_0));
defparam desc2673.INIT=8'hDC;
  LUT4 desc2674(.I0(s_opa_i_2),.I1(s_opa_i_3),.I2(s_opa_i_1),.I3(s_opa_i_0),.O(N_1087));
defparam desc2674.INIT=16'hDCDD;
  LUT4 desc2675(.I0(s_opa_i_2),.I1(s_opa_i_3),.I2(s_opa_i_1),.I3(s_opa_i_0),.O(N_1166));
defparam desc2675.INIT=16'hFFFE;
  LUT3 desc2676(.I0(v_count[2:2]),.I1(N_1619),.I2(N_1624),.O(N_57));
defparam desc2676.INIT=8'hD8;
  LUT3 desc2677(.I0(v_count[2:2]),.I1(N_45),.I2(N_41),.O(N_69));
defparam desc2677.INIT=8'hE4;
  LUT5 desc2678(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(v_count[2:2]),.I3(N_38_0),.I4(N_1620),.O(pre_norm_div_dvdnd[33:33]));
defparam desc2678.INIT=32'h10110001;
  LUT4 desc2679(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(v_count[2:2]),.I3(N_1620),.O(s_dvdnd_50_o_105_0_e));
defparam desc2679.INIT=16'h0100;
  LUT3 desc2680(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd_9),.I2(pre_norm_div_dvdnd_8),.O(pre_norm_sqrt_fracta_o_8));
defparam desc2680.INIT=8'hD8;
  LUT3 desc2681(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd[33:33]),.I2(pre_norm_div_dvdnd_8),.O(pre_norm_sqrt_fracta_o_7));
defparam desc2681.INIT=8'hE4;
  LUT3 desc2682(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd_10),.I2(pre_norm_div_dvdnd_11),.O(pre_norm_sqrt_fracta_o_10));
defparam desc2682.INIT=8'hE4;
  LUT3 desc2683(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd_9),.I2(pre_norm_div_dvdnd_10),.O(pre_norm_sqrt_fracta_o_9));
defparam desc2683.INIT=8'hE4;
  LUT5 desc2684(.I0(s_opa_i_23),.I1(v_count[3:3]),.I2(v_count[4:4]),.I3(N_55),.I4(pre_norm_div_dvdnd[33:33]),.O(pre_norm_sqrt_fracta_o_6));
defparam desc2684.INIT=32'hABAA0100;
  LUT3 desc2685(.I0(v_count[3:3]),.I1(v_count[4:4]),.I2(N_55),.O(s_dvdnd_50_o_108_0_e));
defparam desc2685.INIT=8'h10;
  LUT3 desc2686(.I0(s_opa_i_23),.I1(N_88),.I2(pre_norm_div_dvdnd_16),.O(pre_norm_sqrt_fracta_o_15));
defparam desc2686.INIT=8'hE4;
  LUT3 desc2687(.I0(s_opa_i_23),.I1(pre_norm_div_dvdnd_17),.I2(pre_norm_div_dvdnd_16),.O(pre_norm_sqrt_fracta_o_16));
defparam desc2687.INIT=8'hD8;
endmodule
module sqrt_inj (s_state,s_fracta_52_o_0_e,sqrt_sqr_o,pre_norm_sqrt_fracta_o_0,pre_norm_sqrt_fracta_o_14,pre_norm_sqrt_fracta_o_15,pre_norm_sqrt_fracta_o_16,pre_norm_sqrt_fracta_o_17,pre_norm_sqrt_fracta_o_18,pre_norm_sqrt_fracta_o_19,pre_norm_sqrt_fracta_o_20,pre_norm_sqrt_fracta_o_21,pre_norm_sqrt_fracta_o_22,pre_norm_sqrt_fracta_o_23,pre_norm_sqrt_fracta_o_0_d0,pre_norm_sqrt_fracta_o_1,pre_norm_sqrt_fracta_o_7,pre_norm_sqrt_fracta_o_8,pre_norm_sqrt_fracta_o_9,pre_norm_sqrt_fracta_o_10,pre_norm_sqrt_fracta_o_11,pre_norm_sqrt_fracta_o_12,pre_norm_sqrt_fracta_o_13,s_start_i,un12_s_state_0_a2_lut6_2_O5,clk_i,s_start_i_0,sqrt_ine_o);
input s_state ;
input [33:29] s_fracta_52_o_0_e ;
output [24:0] sqrt_sqr_o ;
input [51:51] pre_norm_sqrt_fracta_o_0 ;
input pre_norm_sqrt_fracta_o_14 ;
input pre_norm_sqrt_fracta_o_15 ;
input pre_norm_sqrt_fracta_o_16 ;
input pre_norm_sqrt_fracta_o_17 ;
input pre_norm_sqrt_fracta_o_18 ;
input pre_norm_sqrt_fracta_o_19 ;
input pre_norm_sqrt_fracta_o_20 ;
input pre_norm_sqrt_fracta_o_21 ;
input pre_norm_sqrt_fracta_o_22 ;
input pre_norm_sqrt_fracta_o_23 ;
input pre_norm_sqrt_fracta_o_0_d0 ;
input pre_norm_sqrt_fracta_o_1 ;
input pre_norm_sqrt_fracta_o_7 ;
input pre_norm_sqrt_fracta_o_8 ;
input pre_norm_sqrt_fracta_o_9 ;
input pre_norm_sqrt_fracta_o_10 ;
input pre_norm_sqrt_fracta_o_11 ;
input pre_norm_sqrt_fracta_o_12 ;
input pre_norm_sqrt_fracta_o_13 ;
output s_start_i ;
output un12_s_state_0_a2_lut6_2_O5 ;
input clk_i ;
input s_start_i_0 ;
output sqrt_ine_o ;
wire pre_norm_sqrt_fracta_o_14 ;
wire pre_norm_sqrt_fracta_o_15 ;
wire pre_norm_sqrt_fracta_o_16 ;
wire pre_norm_sqrt_fracta_o_17 ;
wire pre_norm_sqrt_fracta_o_18 ;
wire pre_norm_sqrt_fracta_o_19 ;
wire pre_norm_sqrt_fracta_o_20 ;
wire pre_norm_sqrt_fracta_o_21 ;
wire pre_norm_sqrt_fracta_o_22 ;
wire pre_norm_sqrt_fracta_o_23 ;
wire pre_norm_sqrt_fracta_o_0_d0 ;
wire pre_norm_sqrt_fracta_o_1 ;
wire pre_norm_sqrt_fracta_o_7 ;
wire pre_norm_sqrt_fracta_o_8 ;
wire pre_norm_sqrt_fracta_o_9 ;
wire pre_norm_sqrt_fracta_o_10 ;
wire pre_norm_sqrt_fracta_o_11 ;
wire pre_norm_sqrt_fracta_o_12 ;
wire pre_norm_sqrt_fracta_o_13 ;
wire s_start_i ;
wire un12_s_state_0_a2_lut6_2_O5 ;
wire clk_i ;
wire s_start_i_0 ;
wire sqrt_ine_o ;
wire [51:0] r1_2 ;
wire [1:0] r1_2_i ;
wire [51:0] r0_2 ;
wire [51:27] s_rad_i ;
wire [4:0] c ;
wire [50:0] un14_s_state_cry ;
wire [25:0] r0 ;
wire [4:0] s_count ;
wire [25:0] r1 ;
wire [25:25] r1_RNIABVR_O5 ;
wire s_state_0 ;
wire [50:0] b_2 ;
wire [10:10] b_2_RNIMF314 ;
wire [22:22] r0_2_RNI9011F_O6 ;
wire [25:0] b ;
wire [51:0] v_r1_2_3 ;
wire [25:0] v_r1_3 ;
wire [24:0] s_sqr_o ;
wire [16:0] un31_s_count_0_data_tmp ;
wire [50:0] un27_s_count_cry ;
wire [11:11] r0_2_RNI351G4 ;
wire [22:22] b_2_RNI46VUE ;
wire [16:16] b_2_RNIRH7KV ;
wire [18:18] b_2_RNI5B6111 ;
wire [14:14] b_2_RNIT9A1G_0 ;
wire [23:23] r0_2_RNIM65S1 ;
wire [14:14] r0_2_RNIMOCU9 ;
wire b_2_fast ;
wire [1:0] r0_2_fast ;
wire c_i ;
wire [26:2] un33_s_count_a_5 ;
wire N_2876_i ;
wire m57_o5_inv ;
wire GND ;
wire VCC ;
wire un14_s_state_df2 ;
wire un14_s_state_lt2 ;
wire un14_s_state_df4 ;
wire un14_s_state_lt4 ;
wire un14_s_state_df6 ;
wire un14_s_state_lt6 ;
wire un14_s_state_df8 ;
wire un14_s_state_lt8 ;
wire un14_s_state_df10 ;
wire un14_s_state_lt10 ;
wire un14_s_state_df12 ;
wire un14_s_state_lt12 ;
wire un14_s_state_df14 ;
wire un14_s_state_lt14 ;
wire un14_s_state_df16 ;
wire un14_s_state_lt16 ;
wire un14_s_state_df18 ;
wire un14_s_state_lt18 ;
wire un14_s_state_df20 ;
wire un14_s_state_lt20 ;
wire un14_s_state_df22 ;
wire un14_s_state_lt22 ;
wire un14_s_state_df24 ;
wire un14_s_state_lt24 ;
wire un14_s_state_df26 ;
wire un14_s_state_lt26 ;
wire un14_s_state_df28 ;
wire un14_s_state_lt28 ;
wire un14_s_state_df30 ;
wire un14_s_state_lt30 ;
wire un14_s_state_df32 ;
wire un14_s_state_lt32 ;
wire un14_s_state_df34 ;
wire un14_s_state_lt34 ;
wire un14_s_state_df36 ;
wire un14_s_state_lt36 ;
wire un14_s_state_df38 ;
wire un14_s_state_lt38 ;
wire un14_s_state_df40 ;
wire un14_s_state_lt40 ;
wire un14_s_state_df42 ;
wire un14_s_state_lt42 ;
wire un14_s_state_df44 ;
wire un14_s_state_lt44 ;
wire un14_s_state_df46 ;
wire un14_s_state_lt46 ;
wire un14_s_state_df48 ;
wire un14_s_state_lt48 ;
wire un14_s_state_df50 ;
wire un14_s_state_lt50 ;
wire un27_s_count_df0 ;
wire un27_s_count_lt0 ;
wire un27_s_count_df2 ;
wire un27_s_count_lt2 ;
wire un27_s_count_df4 ;
wire un27_s_count_lt4 ;
wire un27_s_count_df6 ;
wire un27_s_count_lt6 ;
wire un27_s_count_df8 ;
wire un27_s_count_lt8 ;
wire un27_s_count_df10 ;
wire un27_s_count_lt10 ;
wire un27_s_count_df12 ;
wire un27_s_count_lt12 ;
wire un27_s_count_df14 ;
wire un27_s_count_lt14 ;
wire un27_s_count_df16 ;
wire un27_s_count_lt16 ;
wire un27_s_count_df18 ;
wire un27_s_count_lt18 ;
wire un27_s_count_df20 ;
wire un27_s_count_lt20 ;
wire un27_s_count_df22 ;
wire un27_s_count_lt22 ;
wire un27_s_count_df24 ;
wire un27_s_count_lt24 ;
wire un27_s_count_df26 ;
wire un27_s_count_lt26 ;
wire un27_s_count_df28 ;
wire un27_s_count_lt28 ;
wire un27_s_count_df30 ;
wire un27_s_count_lt30 ;
wire un27_s_count_df32 ;
wire un27_s_count_lt32 ;
wire un27_s_count_df34 ;
wire un27_s_count_lt34 ;
wire un27_s_count_df36 ;
wire un27_s_count_lt36 ;
wire un27_s_count_df38 ;
wire un27_s_count_lt38 ;
wire un27_s_count_df40 ;
wire un27_s_count_lt40 ;
wire un27_s_count_df42 ;
wire un27_s_count_lt42 ;
wire un27_s_count_df44 ;
wire un27_s_count_lt44 ;
wire un27_s_count_df46 ;
wire un27_s_count_lt46 ;
wire un27_s_count_df48 ;
wire un27_s_count_lt48 ;
wire un27_s_count_df50 ;
wire un27_s_count_lt50 ;
wire m143 ;
wire m159 ;
wire m121 ;
wire m180 ;
wire N_48_i ;
wire N_48_i_lut6_2_O5 ;
wire m47 ;
wire N_50_0 ;
wire m168_lut6_2_O6 ;
wire m168_lut6_2_O5 ;
wire m186 ;
wire m166 ;
wire m187_lut6_2_O6 ;
wire m187_lut6_2_O5 ;
wire m189 ;
wire m171 ;
wire m190_lut6_2_O6 ;
wire m190_lut6_2_O5 ;
wire m65 ;
wire m43 ;
wire m56 ;
wire m71_lut6_2_O6 ;
wire m73_lut6_2_O6 ;
wire m73_lut6_2_O5 ;
wire m136 ;
wire m139 ;
wire m141_lut6_2_O6 ;
wire m141_lut6_2_O5 ;
wire N_19_1 ;
wire N_84_0 ;
wire m84 ;
wire m25 ;
wire m26_lut6_2_O6 ;
wire N_86_0 ;
wire N_83_0 ;
wire N_2 ;
wire un3_s_count_0_a2_lut6_2_O6 ;
wire N_22_i_i ;
wire m127_lut6_2_O6 ;
wire m127_lut6_2_O5 ;
wire m154_lut6_2_O6 ;
wire m154_lut6_2_O5 ;
wire m138_lut6_2_O6 ;
wire m138_lut6_2_O5 ;
wire m24_lut6_2_O6 ;
wire m24_lut6_2_O5 ;
wire N_10_1 ;
wire m9_lut6_2_O5 ;
wire N_18_1 ;
wire m17_lut6_2_O5 ;
wire m55_lut6_2_O6 ;
wire m55_lut6_2_O5 ;
wire un33_s_count_a_5_0_axb_26 ;
wire un33_s_count_a_5_0_axb_2 ;
wire un33_s_count_a_5_0_axb_2_lut6_2_O5 ;
wire un12_s_state_0_a2_lut6_2_O6 ;
wire g4_0_2 ;
wire v_r1_2_3_31_0 ;
wire v_r1_2_3_42_0 ;
wire v_r1_2_3_44_lut6_2_O6 ;
wire v_r1_2_3_41_0 ;
wire v_r1_2_3_52_0 ;
wire g0_0_a4_0 ;
wire v_r1_2_3_59_0 ;
wire g0_i_1 ;
wire v_r1_2_3_73_0 ;
wire v_r1_2_3_73_0_lut6_2_O5 ;
wire v_r1_2_3_35_0 ;
wire v_r1_2_3_21_2_RNIMLGQ ;
wire g0_0_a4_0_2 ;
wire v_r1_2_3_35_0_RNI40J52_O5 ;
wire g1_0_0_2 ;
wire g0_0_a4_0_1 ;
wire g4_0_0 ;
wire g1_0_0_1 ;
wire g4_0_1 ;
wire g0_6_0 ;
wire m191 ;
wire m176 ;
wire g0_0_2 ;
wire g4_0_0_1 ;
wire v_r1_2_3_34_0 ;
wire g0_0_a3_0_2 ;
wire g1_1_1 ;
wire v_r1_2_3_21_2 ;
wire v_r1_2_3_27_0 ;
wire v_r1_2_3_21_2_RNIQ1CU_O5 ;
wire N_980_i ;
wire N_981_i ;
wire N_964_i ;
wire N_963_i ;
wire un31_s_count_0_N_116 ;
wire un31_s_count_0_N_109 ;
wire un31_s_count_0_N_102 ;
wire un31_s_count_0_N_95 ;
wire un31_s_count_0_N_88 ;
wire un31_s_count_0_N_81 ;
wire un31_s_count_0_N_74 ;
wire un31_s_count_0_N_67 ;
wire un31_s_count_0_N_60 ;
wire un14_s_state_df0 ;
wire N_2942_i ;
wire v_r1_2_3_73_0_lut6_2_RNIM5CP22 ;
wire v_r1_2_3_0_axb_24 ;
wire un33_s_count_a_5_0_axb_1 ;
wire un33_s_count_a_5_0_axb_3 ;
wire un33_s_count_a_5_0_axb_4 ;
wire un33_s_count_a_5_0_axb_5 ;
wire un33_s_count_a_5_0_axb_6 ;
wire un33_s_count_a_5_0_axb_7 ;
wire un33_s_count_a_5_0_axb_8 ;
wire un33_s_count_a_5_0_axb_9 ;
wire un33_s_count_a_5_0_axb_10 ;
wire un33_s_count_a_5_0_axb_11 ;
wire un33_s_count_a_5_0_axb_12 ;
wire un33_s_count_a_5_0_axb_13 ;
wire un33_s_count_a_5_0_axb_14 ;
wire un33_s_count_a_5_0_axb_15 ;
wire un33_s_count_a_5_0_axb_16 ;
wire un33_s_count_a_5_0_axb_17 ;
wire un33_s_count_a_5_0_axb_18 ;
wire un33_s_count_a_5_0_axb_19 ;
wire un33_s_count_a_5_0_axb_20 ;
wire un33_s_count_a_5_0_axb_21 ;
wire un33_s_count_a_5_0_axb_22 ;
wire un33_s_count_a_5_0_axb_23 ;
wire un33_s_count_a_5_0_axb_24 ;
wire un33_s_count_a_5_0_axb_25 ;
wire un33_s_count_a_5_0_axb_27 ;
wire un33_s_count_a_5_0_axb_28 ;
wire un33_s_count_a_5_0_axb_29 ;
wire un33_s_count_a_5_0_axb_30 ;
wire un33_s_count_a_5_0_axb_31 ;
wire un33_s_count_a_5_0_axb_32 ;
wire un33_s_count_a_5_0_axb_33 ;
wire un33_s_count_a_5_0_axb_34 ;
wire un33_s_count_a_5_0_axb_35 ;
wire un33_s_count_a_5_0_axb_36 ;
wire un33_s_count_a_5_0_axb_37 ;
wire un33_s_count_a_5_0_axb_38 ;
wire un33_s_count_a_5_0_axb_39 ;
wire un33_s_count_a_5_0_axb_40 ;
wire un33_s_count_a_5_0_axb_41 ;
wire un33_s_count_a_5_0_axb_42 ;
wire un33_s_count_a_5_0_axb_43 ;
wire un33_s_count_a_5_0_axb_44 ;
wire un33_s_count_a_5_0_axb_45 ;
wire un33_s_count_a_5_0_axb_46 ;
wire un33_s_count_a_5_0_axb_47 ;
wire un33_s_count_a_5_0_axb_48 ;
wire un33_s_count_a_5_0_axb_49 ;
wire un33_s_count_a_5_0_axb_50 ;
wire v_r1_3_axb_0 ;
wire v_r1_3_axb_1 ;
wire v_r1_3_axb_2 ;
wire v_r1_3_axb_3 ;
wire v_r1_3_axb_4 ;
wire v_r1_3_axb_5 ;
wire v_r1_3_axb_6 ;
wire v_r1_3_axb_7 ;
wire v_r1_3_axb_8 ;
wire v_r1_3_axb_9 ;
wire v_r1_3_axb_10 ;
wire v_r1_3_axb_11 ;
wire v_r1_3_axb_12 ;
wire v_r1_3_axb_13 ;
wire v_r1_3_axb_14 ;
wire v_r1_3_axb_15 ;
wire v_r1_3_axb_16 ;
wire v_r1_3_axb_17 ;
wire v_r1_3_axb_18 ;
wire v_r1_3_axb_19 ;
wire v_r1_3_axb_20 ;
wire v_r1_3_axb_21 ;
wire v_r1_3_axb_22 ;
wire v_r1_3_axb_23 ;
wire v_r1_3_axb_24 ;
wire v_r1_2_3_scalar ;
wire un31_s_count_0_N_3_i ;
wire s_ine_o ;
wire s_ine_o_0 ;
wire un31_s_count_0_I_139 ;
wire g0_5i0 ;
wire g0_5i1 ;
wire v_r1_2_3_56_0_tz ;
wire v_r1_2_3_35_0_RNIKOE74 ;
wire g3 ;
wire v_r1_2_3_63_2 ;
wire v_r1_2_3_72_0_N_2L1 ;
wire g2_0 ;
wire v_r1_2_3_49_0_tz ;
wire m45 ;
wire v_r1_2_3_28 ;
wire v_r1_2_3_65_c ;
wire v_r1_2_3_0_axb_22 ;
wire N_4 ;
wire g4_0 ;
wire g1_0 ;
wire v_r1_2_3_0_axb_21 ;
wire g0_0_0_0 ;
wire g4_0_0_0 ;
wire g4_1 ;
wire v_r1_2_3_31 ;
wire v_r1_2_3_0_cry_9_RNO ;
wire v_r1_2_3_22 ;
wire g5_0 ;
wire v_r1_2_3_65_0_0 ;
wire v_r1_2_3_77_0_tz ;
wire g0_0_a4_3 ;
wire v_r1_2_3_4 ;
wire v_r1_2_3_14_0 ;
wire N_5_0_0 ;
wire v_r1_2_3_28_0_tz ;
wire g0_i_0 ;
wire N_4_1 ;
wire v_r1_2_3_10 ;
wire g0_i_a3_0 ;
wire v_r1_2_3_48_0 ;
wire N_4_0 ;
wire g2_1_0 ;
wire N_6_1_0 ;
wire v_r1_2_3_14 ;
wire N_89_0 ;
wire N_12_1 ;
wire N_90_0 ;
wire m32 ;
wire m36 ;
wire m157 ;
wire m110 ;
wire m169 ;
wire m112 ;
wire m114 ;
wire m113 ;
wire m174 ;
wire v_r1_2_3_23 ;
wire m132 ;
wire v_r1_2_3_0_axb_8 ;
wire v_r1_2_3_0_cry_8_RNO ;
wire v_r1_2_3_63_2_0 ;
wire v_r1_2_3_25 ;
wire v_r1_2_3_0_axb_20 ;
wire v_r1_2_3_0_cry_20_RNO ;
wire m145 ;
wire m125 ;
wire v_r1_2_3_51 ;
wire v_r1_2_3_0_axb_16 ;
wire v_r1_2_3_9 ;
wire v_r1_2_3_0_axb_4 ;
wire v_r1_2_3_0_cry_4_RNO ;
wire m193 ;
wire v_r1_2_3_0_axb_1 ;
wire v_r1_2_3_0_cry_18_RNO ;
wire v_r1_2_3_0_axb_10 ;
wire m129 ;
wire v_r1_2_3_0_axb_12 ;
wire v_r1_2_3_16 ;
wire v_r1_2_3_0_axb_6 ;
wire m67 ;
wire v_r1_2_3_0_axb_14 ;
wire v_r1_2_3_2 ;
wire v_r1_2_3_0_axb_2 ;
wire v_r1_2_3_0_cry_1_RNO ;
wire v_r1_2_3_0_cry_2_RNO ;
wire v_r1_2_3_0_cry_3_RNO ;
wire m35 ;
wire m90 ;
wire N_95_0 ;
wire N_96_0 ;
wire m207 ;
wire N_3022_i ;
wire v_r1_2_3_0_cry_7_RNO ;
wire v_r1_2_3_0_cry_6_RNO ;
wire v_r1_2_3_0_cry_45_RNO ;
wire v_r1_2_3_0_cry_46_RNO ;
wire m100 ;
wire m108 ;
wire m182 ;
wire v_r1_2_3_0_cry_31_RNO ;
wire v_r1_2_3_0_cry_30_RNO ;
wire v_r1_2_3_0_cry_41_RNO ;
wire v_r1_2_3_0_cry_34_RNO ;
wire m203 ;
wire m200 ;
wire v_r1_2_3_0_cry_43_RNO ;
wire v_r1_2_3_0_cry_47_RNO ;
wire v_r1_2_3_0_cry_42_RNO ;
wire v_r1_2_3_0_cry_44_RNO ;
wire v_r1_2_3_0_cry_48_RNO ;
wire v_r1_2_3_0_cry_32_RNO ;
wire v_r1_2_3_0_cry_26_RNO ;
wire m211 ;
wire N_2891_i ;
wire v_r1_2_3_0_axb_27 ;
wire v_r1_2_3_175 ;
wire v_r1_2_3_0_cry_33_RNO ;
wire v_r1_2_3_0_cry_10_RNO ;
wire v_r1_2_3_0_cry_29_RNO ;
wire m210 ;
wire v_r1_2_3_0_cry_28_RNO ;
wire v_r1_2_3_0_cry_35_RNO ;
wire v_r1_2_3_0_cry_36_RNO ;
wire v_r1_2_3_0_cry_12_RNO ;
wire v_r1_2_3_0_cry_14_RNO ;
wire v_r1_2_3_0_cry_16_RNO ;
wire N_2895_i ;
wire v_r1_2_3_0_axb_18 ;
wire v_r1_2_3_49 ;
wire v_r1_2_3_0_cry_17_RNO ;
wire v_r1_2_3_0_cry_22_RNO ;
wire v_r1_2_3_0_cry_21_RNO ;
wire v_r1_2_3_0_axb_25 ;
wire v_r1_2_3_0_cry_0_cy ;
wire un1_r1_axb_24 ;
wire un1_r1_axb_23 ;
wire un1_r1_axb_22 ;
wire un1_r1_axb_21 ;
wire un1_r1_axb_20 ;
wire un1_r1_axb_19 ;
wire un1_r1_axb_18 ;
wire un1_r1_axb_17 ;
wire un1_r1_axb_16 ;
wire un1_r1_axb_15 ;
wire un1_r1_axb_14 ;
wire un1_r1_axb_13 ;
wire un1_r1_axb_12 ;
wire un1_r1_axb_11 ;
wire un1_r1_axb_10 ;
wire un1_r1_axb_9 ;
wire un1_r1_axb_8 ;
wire un1_r1_axb_7 ;
wire un1_r1_axb_6 ;
wire un1_r1_axb_5 ;
wire un1_r1_axb_4 ;
wire un1_r1_axb_3 ;
wire un1_r1_axb_2 ;
wire un1_r1_axb_1 ;
wire un1_r1_axb_0 ;
wire v_r1_2_3_0 ;
wire un33_s_count_NE_1_3 ;
wire un33_s_count_NE_0_3 ;
wire un33_s_count_a_5_0_o5_16 ;
wire un33_s_count_a_5_0_o5_21 ;
wire un33_s_count_a_5_0_o5_17 ;
wire un33_s_count_a_5_0_o5_4 ;
wire un33_s_count_a_5_0_o5_20 ;
wire un33_s_count_a_5_0_o5_18 ;
wire un33_s_count_a_5_0_o5_6 ;
wire un33_s_count_a_5_0_o5_3 ;
wire un33_s_count_a_5_0_o5_14 ;
wire un33_s_count_a_5_0_o5_23 ;
wire un33_s_count_a_5_0_o5_9 ;
wire un33_s_count_a_5_0_o5_10 ;
wire un33_s_count_a_5_0_o5_15 ;
wire un33_s_count_a_5_0_o5_19 ;
wire un33_s_count_a_5_0_o5_5 ;
wire un33_s_count_a_5_0_o5_8 ;
wire un33_s_count_a_5_0_o5_12 ;
wire un33_s_count_a_5_0_o5_24 ;
wire un33_s_count_a_5_0_o5_22 ;
wire un33_s_count_a_5_0_o5_13 ;
wire un33_s_count_a_5_0_o5_7 ;
wire un33_s_count_a_5_0_o5_11 ;
wire v_r1_3_axb_25 ;
wire un33_s_count_a_5_0_axb_51 ;
wire m109 ;
wire m106 ;
wire m105 ;
wire m42 ;
wire un33_s_count_29 ;
wire un33_s_count_30 ;
wire un33_s_count_31 ;
wire un33_s_count_32 ;
wire un33_s_count_33 ;
wire un33_s_count_34 ;
wire un33_s_count_NE_5 ;
wire un33_s_count_NE_3 ;
wire un33_s_count_NE_2 ;
wire un31_s_count_0_N_4 ;
wire un31_s_count_0_N_46 ;
wire un31_s_count_0_N_25 ;
wire un31_s_count_0_N_53 ;
wire un31_s_count_0_N_32 ;
wire un31_s_count_0_N_18 ;
wire un31_s_count_0_N_11 ;
wire un31_s_count_0_N_39 ;
wire v_r1_2_3_0_o5_26 ;
wire v_r1_2_3_0_o5_24 ;
wire m178 ;
wire m164 ;
wire m156 ;
wire m123 ;
wire m119 ;
wire m104 ;
wire un33_s_count_37 ;
wire un33_s_count_38 ;
wire un33_s_count_39 ;
wire un33_s_count_NE_6_3 ;
wire un33_s_count_1 ;
wire un33_s_count_27 ;
wire un33_s_count_28 ;
wire un33_s_count_NE_4_3 ;
wire v_r1_2_3_7 ;
wire m115 ;
wire un33_s_count_45 ;
wire un33_s_count_46 ;
wire un33_s_count_47 ;
wire un33_s_count_48 ;
wire un33_s_count_49 ;
wire un33_s_count_NE_8 ;
wire un33_s_count_40 ;
wire un33_s_count_41 ;
wire un33_s_count_42 ;
wire un33_s_count_43 ;
wire un33_s_count_44 ;
wire un33_s_count_NE_7 ;
wire un33_s_count_35 ;
wire un33_s_count_36 ;
wire un33_s_count_50 ;
wire un33_s_count_51 ;
wire un33_s_count_NE_1_4 ;
wire un33_s_count_NE_2_4 ;
wire m208 ;
wire m205 ;
wire m183 ;
wire m177 ;
wire m162 ;
wire m160 ;
wire m126 ;
wire m122 ;
wire m117 ;
wire m97 ;
wire N_93_0 ;
wire m87 ;
wire m59 ;
wire N_47_0 ;
wire N_29_0 ;
wire N_2951_i ;
wire v_r1_2_3_0_axb_0 ;
wire N_2939_i ;
wire N_2887_i ;
wire v_r1_2_3_0_axb_51 ;
wire v_r1_2_3_63_0_c ;
wire v_r1_2_3_56 ;
wire v_r1_2_3_63_0_d ;
wire v_r1_2_3_0_axb_3 ;
wire v_r1_2_3_0_axb_5 ;
wire v_r1_2_3_0_cry_5_RNO ;
wire v_r1_2_3_0_axb_7 ;
wire v_r1_2_3_0_axb_9 ;
wire v_r1_2_3_0_axb_11 ;
wire v_r1_2_3_0_cry_11_RNO ;
wire v_r1_2_3_0_axb_13 ;
wire v_r1_2_3_0_cry_13_RNO ;
wire v_r1_2_3_0_axb_15 ;
wire v_r1_2_3_0_cry_15_RNO ;
wire v_r1_2_3_0_axb_17 ;
wire v_r1_2_3_0_axb_19 ;
wire v_r1_2_3_0_cry_19_RNO ;
wire v_r1_2_3_0_axb_23 ;
wire v_r1_2_3_0_cry_23_RNO ;
wire v_r1_2_3_0_cry_24_RNO ;
wire v_r1_2_3_0_axb_26 ;
wire v_r1_2_3_0_axb_28 ;
wire v_r1_2_3_0_axb_29 ;
wire v_r1_2_3_0_axb_30 ;
wire v_r1_2_3_0_axb_31 ;
wire v_r1_2_3_0_axb_32 ;
wire v_r1_2_3_0_axb_33 ;
wire v_r1_2_3_0_axb_34 ;
wire v_r1_2_3_0_axb_35 ;
wire v_r1_2_3_0_axb_36 ;
wire v_r1_2_3_0_axb_37 ;
wire v_r1_2_3_0_cry_37_RNO ;
wire v_r1_2_3_0_axb_38 ;
wire v_r1_2_3_0_cry_38_RNO ;
wire v_r1_2_3_0_axb_39 ;
wire v_r1_2_3_0_cry_39_RNO ;
wire v_r1_2_3_0_axb_40 ;
wire v_r1_2_3_0_cry_40_RNO ;
wire v_r1_2_3_0_axb_41 ;
wire v_r1_2_3_0_axb_42 ;
wire v_r1_2_3_0_axb_43 ;
wire v_r1_2_3_0_axb_44 ;
wire v_r1_2_3_0_axb_45 ;
wire v_r1_2_3_0_axb_46 ;
wire v_r1_2_3_0_axb_47 ;
wire v_r1_2_3_0_axb_48 ;
wire v_r1_2_3_0_axb_49 ;
wire v_r1_2_3_0_cry_49_RNO ;
wire v_r1_2_3_0_axb_50 ;
wire v_r1_2_3_0_cry_50_RNO ;
wire un33_s_count_a_5_0_cry_26_RNO ;
wire un33_s_count_a_5_0_cry_28_RNO ;
wire un33_s_count_a_5_0_cry_29_RNO ;
wire un33_s_count_a_5_0_cry_30_RNO ;
wire un33_s_count_a_5_0_cry_31_RNO ;
wire un33_s_count_a_5_0_cry_32_RNO ;
wire un33_s_count_a_5_0_cry_33_RNO ;
wire un33_s_count_a_5_0_cry_34_RNO ;
wire un33_s_count_a_5_0_cry_35_RNO ;
wire un33_s_count_a_5_0_cry_36_RNO ;
wire un33_s_count_a_5_0_cry_37_RNO ;
wire un33_s_count_a_5_0_cry_38_RNO ;
wire un33_s_count_a_5_0_cry_39_RNO ;
wire un33_s_count_a_5_0_cry_40_RNO ;
wire un33_s_count_a_5_0_cry_41_RNO ;
wire un33_s_count_a_5_0_cry_42_RNO ;
wire un33_s_count_a_5_0_cry_43_RNO ;
wire un33_s_count_a_5_0_cry_44_RNO ;
wire un33_s_count_a_5_0_cry_45_RNO ;
wire un33_s_count_a_5_0_cry_46_RNO ;
wire un33_s_count_a_5_0_cry_47_RNO ;
wire un33_s_count_a_5_0_cry_48_RNO ;
wire un33_s_count_a_5_0_cry_49_RNO ;
wire un33_s_count_a_5_0_cry_50_RNO ;
wire un1_r1_cry_23 ;
wire un1_r1_s_24 ;
wire un1_r1_cry_22 ;
wire un1_r1_s_23 ;
wire un1_r1_cry_21 ;
wire un1_r1_s_22 ;
wire un1_r1_cry_20 ;
wire un1_r1_s_21 ;
wire un1_r1_cry_19 ;
wire un1_r1_s_20 ;
wire un1_r1_cry_18 ;
wire un1_r1_s_19 ;
wire un1_r1_cry_17 ;
wire un1_r1_s_18 ;
wire un1_r1_cry_16 ;
wire un1_r1_s_17 ;
wire un1_r1_cry_15 ;
wire un1_r1_s_16 ;
wire un1_r1_cry_14 ;
wire un1_r1_s_15 ;
wire un1_r1_cry_13 ;
wire un1_r1_s_14 ;
wire un1_r1_cry_12 ;
wire un1_r1_s_13 ;
wire un1_r1_cry_11 ;
wire un1_r1_s_12 ;
wire un1_r1_cry_10 ;
wire un1_r1_s_11 ;
wire un1_r1_cry_9 ;
wire un1_r1_s_10 ;
wire un1_r1_cry_8 ;
wire un1_r1_s_9 ;
wire un1_r1_cry_7 ;
wire un1_r1_s_8 ;
wire un1_r1_cry_6 ;
wire un1_r1_s_7 ;
wire un1_r1_cry_5 ;
wire un1_r1_s_6 ;
wire un1_r1_cry_4 ;
wire un1_r1_s_5 ;
wire un1_r1_cry_3 ;
wire un1_r1_s_4 ;
wire un1_r1_cry_2 ;
wire un1_r1_s_3 ;
wire un1_r1_cry_1 ;
wire un1_r1_s_2 ;
wire un1_r1_cry_0 ;
wire un1_r1_s_1 ;
wire v_r1_3_cry_24 ;
wire v_r1_3_cry_23 ;
wire v_r1_3_cry_22 ;
wire v_r1_3_cry_21 ;
wire v_r1_3_cry_20 ;
wire v_r1_3_cry_19 ;
wire v_r1_3_cry_18 ;
wire v_r1_3_cry_17 ;
wire v_r1_3_cry_16 ;
wire v_r1_3_cry_15 ;
wire v_r1_3_cry_14 ;
wire v_r1_3_cry_13 ;
wire v_r1_3_cry_12 ;
wire v_r1_3_cry_11 ;
wire v_r1_3_cry_10 ;
wire v_r1_3_cry_9 ;
wire v_r1_3_cry_8 ;
wire v_r1_3_cry_7 ;
wire v_r1_3_cry_6 ;
wire v_r1_3_cry_5 ;
wire v_r1_3_cry_4 ;
wire v_r1_3_cry_3 ;
wire v_r1_3_cry_2 ;
wire v_r1_3_cry_1 ;
wire v_r1_3_cry_0 ;
wire un33_s_count_a_5_0_cry_50 ;
wire un33_s_count_a_5_0_cry_49 ;
wire un33_s_count_a_5_0_cry_48 ;
wire un33_s_count_a_5_0_cry_47 ;
wire un33_s_count_a_5_0_cry_46 ;
wire un33_s_count_a_5_0_cry_45 ;
wire un33_s_count_a_5_0_cry_44 ;
wire un33_s_count_a_5_0_cry_43 ;
wire un33_s_count_a_5_0_cry_42 ;
wire un33_s_count_a_5_0_cry_41 ;
wire un33_s_count_a_5_0_cry_40 ;
wire un33_s_count_a_5_0_cry_39 ;
wire un33_s_count_a_5_0_cry_38 ;
wire un33_s_count_a_5_0_cry_37 ;
wire un33_s_count_a_5_0_cry_36 ;
wire un33_s_count_a_5_0_cry_35 ;
wire un33_s_count_a_5_0_cry_34 ;
wire un33_s_count_a_5_0_cry_33 ;
wire un33_s_count_a_5_0_cry_32 ;
wire un33_s_count_a_5_0_cry_31 ;
wire un33_s_count_a_5_0_cry_30 ;
wire un33_s_count_a_5_0_cry_29 ;
wire un33_s_count_a_5_0_cry_28 ;
wire un33_s_count_a_5_0_cry_27 ;
wire un33_s_count_a_5_0_cry_26 ;
wire un33_s_count_a_5_0_cry_25 ;
wire un33_s_count_a_5_0_cry_24 ;
wire un33_s_count_a_5_0_cry_23 ;
wire un33_s_count_a_5_0_cry_22 ;
wire un33_s_count_a_5_0_cry_21 ;
wire un33_s_count_a_5_0_cry_20 ;
wire un33_s_count_a_5_0_cry_19 ;
wire un33_s_count_a_5_0_cry_18 ;
wire un33_s_count_a_5_0_cry_17 ;
wire un33_s_count_a_5_0_cry_16 ;
wire un33_s_count_a_5_0_cry_15 ;
wire un33_s_count_a_5_0_cry_14 ;
wire un33_s_count_a_5_0_cry_13 ;
wire un33_s_count_a_5_0_cry_12 ;
wire un33_s_count_a_5_0_cry_11 ;
wire un33_s_count_a_5_0_cry_10 ;
wire un33_s_count_a_5_0_cry_9 ;
wire un33_s_count_a_5_0_cry_8 ;
wire un33_s_count_a_5_0_cry_7 ;
wire un33_s_count_a_5_0_cry_6 ;
wire un33_s_count_a_5_0_cry_5 ;
wire un33_s_count_a_5_0_cry_4 ;
wire un33_s_count_a_5_0_cry_3 ;
wire un33_s_count_a_5_0_cry_2 ;
wire un33_s_count_a_5_0_cry_1 ;
wire un33_s_count_a_5_0_cry_0 ;
wire v_r1_2_3_0_cry_50 ;
wire v_r1_2_3_0_cry_49 ;
wire v_r1_2_3_0_cry_48 ;
wire v_r1_2_3_0_cry_47 ;
wire v_r1_2_3_0_cry_46 ;
wire v_r1_2_3_0_cry_45 ;
wire v_r1_2_3_0_cry_44 ;
wire v_r1_2_3_0_cry_43 ;
wire v_r1_2_3_0_cry_42 ;
wire v_r1_2_3_0_cry_41 ;
wire v_r1_2_3_0_cry_40 ;
wire v_r1_2_3_0_cry_39 ;
wire v_r1_2_3_0_cry_38 ;
wire v_r1_2_3_0_cry_37 ;
wire v_r1_2_3_0_cry_36 ;
wire v_r1_2_3_0_cry_35 ;
wire v_r1_2_3_0_cry_34 ;
wire v_r1_2_3_0_cry_33 ;
wire v_r1_2_3_0_cry_32 ;
wire v_r1_2_3_0_cry_31 ;
wire v_r1_2_3_0_cry_30 ;
wire v_r1_2_3_0_cry_29 ;
wire v_r1_2_3_0_cry_28 ;
wire v_r1_2_3_0_cry_27 ;
wire v_r1_2_3_0_cry_26 ;
wire v_r1_2_3_0_cry_25 ;
wire v_r1_2_3_0_cry_24 ;
wire v_r1_2_3_0_cry_23 ;
wire v_r1_2_3_0_cry_22 ;
wire v_r1_2_3_0_cry_21 ;
wire v_r1_2_3_0_cry_20 ;
wire v_r1_2_3_0_cry_19 ;
wire v_r1_2_3_0_cry_18 ;
wire v_r1_2_3_0_cry_17 ;
wire v_r1_2_3_0_cry_16 ;
wire v_r1_2_3_0_cry_15 ;
wire v_r1_2_3_0_cry_14 ;
wire v_r1_2_3_0_cry_13 ;
wire v_r1_2_3_0_cry_12 ;
wire v_r1_2_3_0_cry_11 ;
wire v_r1_2_3_0_cry_10 ;
wire v_r1_2_3_0_cry_9 ;
wire v_r1_2_3_0_cry_8 ;
wire v_r1_2_3_0_cry_7 ;
wire v_r1_2_3_0_cry_6 ;
wire v_r1_2_3_0_cry_5 ;
wire v_r1_2_3_0_cry_4 ;
wire v_r1_2_3_0_cry_3 ;
wire v_r1_2_3_0_cry_2 ;
wire v_r1_2_3_0_cry_1 ;
wire v_r1_2_3_0_cry_0 ;
wire N_171 ;
wire N_170 ;
wire N_169 ;
wire N_168 ;
wire N_167 ;
wire N_166 ;
wire N_165 ;
wire N_164 ;
wire N_163 ;
wire N_162 ;
wire N_161 ;
wire N_160 ;
wire N_159 ;
wire N_158 ;
wire N_157 ;
wire N_156 ;
wire N_155 ;
wire N_154 ;
wire N_153 ;
wire N_152 ;
wire N_151 ;
wire N_150 ;
wire N_149 ;
wire N_148 ;
wire N_147 ;
wire N_146 ;
wire N_145 ;
wire N_144 ;
wire N_143 ;
wire N_142 ;
wire N_141 ;
wire N_140 ;
wire N_139 ;
wire N_138 ;
wire N_137 ;
wire N_136 ;
wire N_135 ;
wire N_134 ;
wire N_133 ;
wire N_132 ;
wire un14_s_state_lt0 ;
wire N_130 ;
wire N_129 ;
wire N_128 ;
wire N_127 ;
wire N_126 ;
wire N_125 ;
wire N_124 ;
wire N_123 ;
wire N_122 ;
wire N_121 ;
wire N_120 ;
wire N_119 ;
wire N_118 ;
wire N_117 ;
wire N_116 ;
wire N_115 ;
wire N_114 ;
wire N_113 ;
wire N_112 ;
wire N_111 ;
wire N_110 ;
wire N_109 ;
wire N_108 ;
wire N_107 ;
wire N_106 ;
wire N_105 ;
wire N_104 ;
wire N_103 ;
wire N_102 ;
wire N_2_0 ;
wire N_1 ;
// instances
  LUT1 un33_s_count_a_5_0_cry_1_RNO(.I0(r1_2[1:1]),.O(r1_2_i[1:1]));
defparam un33_s_count_a_5_0_cry_1_RNO.INIT=2'h1;
  INV desc2688(.I(N_2876_i),.O(m57_o5_inv));
  LUT6_2 desc2689(.I0(c[2:2]),.I1(un14_s_state_cry[50:50]),.I2(m65),.I3(m43),.I4(m56),.I5(c[3:3]),.O6(m71_lut6_2_O6),.O5(N_2876_i));
defparam desc2689.INIT=64'h727272720055AAFF;
  FD desc2690(.Q(s_rad_i[33:33]),.D(s_fracta_52_o_0_e[33:33]),.C(clk_i));
  FD desc2691(.Q(s_rad_i[32:32]),.D(s_fracta_52_o_0_e[32:32]),.C(clk_i));
  FD desc2692(.Q(s_rad_i[31:31]),.D(s_fracta_52_o_0_e[31:31]),.C(clk_i));
  FD desc2693(.Q(s_rad_i[30:30]),.D(s_fracta_52_o_0_e[30:30]),.C(clk_i));
  FD desc2694(.Q(s_rad_i[29:29]),.D(s_fracta_52_o_0_e[29:29]),.C(clk_i));
  FDSE desc2695(.Q(s_state_0),.D(GND),.C(clk_i),.S(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDSE desc2696(.Q(s_count[1:1]),.D(N_22_i_i),.C(clk_i),.S(s_start_i),.CE(s_state_0));
  FDSE desc2697(.Q(s_count[3:3]),.D(N_980_i),.C(clk_i),.S(s_start_i),.CE(s_state_0));
  FDRE desc2698(.Q(s_count[2:2]),.D(N_964_i),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDSE desc2699(.Q(s_count[4:4]),.D(N_981_i),.C(clk_i),.S(s_start_i),.CE(s_state_0));
  FDRE desc2700(.Q(s_count[0:0]),.D(N_963_i),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  LUT3 un31_s_count_0_I_10(.I0(r1_2[0:0]),.I1(r1_2[1:1]),.I2(r1_2[2:2]),.O(un31_s_count_0_N_116));
defparam un31_s_count_0_I_10.INIT=8'h01;
  LUT3 un31_s_count_0_I_18(.I0(r1_2[3:3]),.I1(r1_2[4:4]),.I2(r1_2[5:5]),.O(un31_s_count_0_N_109));
defparam un31_s_count_0_I_18.INIT=8'h01;
  LUT3 un31_s_count_0_I_26(.I0(r1_2[6:6]),.I1(r1_2[7:7]),.I2(r1_2[8:8]),.O(un31_s_count_0_N_102));
defparam un31_s_count_0_I_26.INIT=8'h01;
  LUT3 un31_s_count_0_I_34(.I0(r1_2[9:9]),.I1(r1_2[10:10]),.I2(r1_2[11:11]),.O(un31_s_count_0_N_95));
defparam un31_s_count_0_I_34.INIT=8'h01;
  LUT3 un31_s_count_0_I_42(.I0(r1_2[12:12]),.I1(r1_2[13:13]),.I2(r1_2[14:14]),.O(un31_s_count_0_N_88));
defparam un31_s_count_0_I_42.INIT=8'h01;
  LUT3 un31_s_count_0_I_50(.I0(r1_2[15:15]),.I1(r1_2[16:16]),.I2(r1_2[17:17]),.O(un31_s_count_0_N_81));
defparam un31_s_count_0_I_50.INIT=8'h01;
  LUT3 un31_s_count_0_I_58(.I0(r1_2[18:18]),.I1(r1_2[19:19]),.I2(r1_2[20:20]),.O(un31_s_count_0_N_74));
defparam un31_s_count_0_I_58.INIT=8'h01;
  LUT3 un31_s_count_0_I_66(.I0(r1_2[21:21]),.I1(r1_2[22:22]),.I2(r1_2[23:23]),.O(un31_s_count_0_N_67));
defparam un31_s_count_0_I_66.INIT=8'h01;
  LUT3 un31_s_count_0_I_74(.I0(r1_2[24:24]),.I1(r1_2[25:25]),.I2(r1_2[26:26]),.O(un31_s_count_0_N_60));
defparam un31_s_count_0_I_74.INIT=8'h01;
  LUT2 un14_s_state_df0_cZ(.I0(r0_2[0:0]),.I1(r0_2[1:1]),.O(un14_s_state_df0));
defparam un14_s_state_df0_cZ.INIT=4'h1;
  LUT4 desc2701(.I0(N_2942_i),.I1(v_r1_2_3_73_0_lut6_2_RNIM5CP22),.I2(b_2[24:24]),.I3(r0_2[24:24]),.O(v_r1_2_3_0_axb_24));
defparam desc2701.INIT=16'h6996;
  LUT1 un33_s_count_a_5_0_cry_0_RNO(.I0(r1_2[0:0]),.O(r1_2_i[0:0]));
defparam un33_s_count_a_5_0_cry_0_RNO.INIT=2'h1;
  LUT2 desc2702(.I0(r1[0:0]),.I1(r1_2[1:1]),.O(un33_s_count_a_5_0_axb_1));
defparam desc2702.INIT=4'h6;
  LUT4 un33_s_count_a_5_0_axb_3_cZ(.I0(r1[1:1]),.I1(r1[2:2]),.I2(r1_2[2:2]),.I3(r1_2[3:3]),.O(un33_s_count_a_5_0_axb_3));
defparam un33_s_count_a_5_0_axb_3_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_4_cZ(.I0(r1[2:2]),.I1(r1[3:3]),.I2(r1_2[3:3]),.I3(r1_2[4:4]),.O(un33_s_count_a_5_0_axb_4));
defparam un33_s_count_a_5_0_axb_4_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_5_cZ(.I0(r1[3:3]),.I1(r1[4:4]),.I2(r1_2[4:4]),.I3(r1_2[5:5]),.O(un33_s_count_a_5_0_axb_5));
defparam un33_s_count_a_5_0_axb_5_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_6_cZ(.I0(r1[4:4]),.I1(r1[5:5]),.I2(r1_2[5:5]),.I3(r1_2[6:6]),.O(un33_s_count_a_5_0_axb_6));
defparam un33_s_count_a_5_0_axb_6_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_7_cZ(.I0(r1[5:5]),.I1(r1[6:6]),.I2(r1_2[6:6]),.I3(r1_2[7:7]),.O(un33_s_count_a_5_0_axb_7));
defparam un33_s_count_a_5_0_axb_7_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_8_cZ(.I0(r1[6:6]),.I1(r1[7:7]),.I2(r1_2[7:7]),.I3(r1_2[8:8]),.O(un33_s_count_a_5_0_axb_8));
defparam un33_s_count_a_5_0_axb_8_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_9_cZ(.I0(r1[7:7]),.I1(r1[8:8]),.I2(r1_2[8:8]),.I3(r1_2[9:9]),.O(un33_s_count_a_5_0_axb_9));
defparam un33_s_count_a_5_0_axb_9_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_10_cZ(.I0(r1[8:8]),.I1(r1[9:9]),.I2(r1_2[9:9]),.I3(r1_2[10:10]),.O(un33_s_count_a_5_0_axb_10));
defparam un33_s_count_a_5_0_axb_10_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_11_cZ(.I0(r1[9:9]),.I1(r1[10:10]),.I2(r1_2[10:10]),.I3(r1_2[11:11]),.O(un33_s_count_a_5_0_axb_11));
defparam un33_s_count_a_5_0_axb_11_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_12_cZ(.I0(r1[10:10]),.I1(r1[11:11]),.I2(r1_2[11:11]),.I3(r1_2[12:12]),.O(un33_s_count_a_5_0_axb_12));
defparam un33_s_count_a_5_0_axb_12_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_13_cZ(.I0(r1[11:11]),.I1(r1[12:12]),.I2(r1_2[12:12]),.I3(r1_2[13:13]),.O(un33_s_count_a_5_0_axb_13));
defparam un33_s_count_a_5_0_axb_13_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_14_cZ(.I0(r1[12:12]),.I1(r1[13:13]),.I2(r1_2[13:13]),.I3(r1_2[14:14]),.O(un33_s_count_a_5_0_axb_14));
defparam un33_s_count_a_5_0_axb_14_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_15_cZ(.I0(r1[13:13]),.I1(r1[14:14]),.I2(r1_2[14:14]),.I3(r1_2[15:15]),.O(un33_s_count_a_5_0_axb_15));
defparam un33_s_count_a_5_0_axb_15_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_16_cZ(.I0(r1[14:14]),.I1(r1[15:15]),.I2(r1_2[15:15]),.I3(r1_2[16:16]),.O(un33_s_count_a_5_0_axb_16));
defparam un33_s_count_a_5_0_axb_16_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_17_cZ(.I0(r1[15:15]),.I1(r1[16:16]),.I2(r1_2[16:16]),.I3(r1_2[17:17]),.O(un33_s_count_a_5_0_axb_17));
defparam un33_s_count_a_5_0_axb_17_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_18_cZ(.I0(r1[16:16]),.I1(r1[17:17]),.I2(r1_2[17:17]),.I3(r1_2[18:18]),.O(un33_s_count_a_5_0_axb_18));
defparam un33_s_count_a_5_0_axb_18_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_19_cZ(.I0(r1[17:17]),.I1(r1[18:18]),.I2(r1_2[18:18]),.I3(r1_2[19:19]),.O(un33_s_count_a_5_0_axb_19));
defparam un33_s_count_a_5_0_axb_19_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_20_cZ(.I0(r1[18:18]),.I1(r1[19:19]),.I2(r1_2[19:19]),.I3(r1_2[20:20]),.O(un33_s_count_a_5_0_axb_20));
defparam un33_s_count_a_5_0_axb_20_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_21_cZ(.I0(r1[19:19]),.I1(r1[20:20]),.I2(r1_2[20:20]),.I3(r1_2[21:21]),.O(un33_s_count_a_5_0_axb_21));
defparam un33_s_count_a_5_0_axb_21_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_22_cZ(.I0(r1[20:20]),.I1(r1[21:21]),.I2(r1_2[21:21]),.I3(r1_2[22:22]),.O(un33_s_count_a_5_0_axb_22));
defparam un33_s_count_a_5_0_axb_22_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_23_cZ(.I0(r1[21:21]),.I1(r1[22:22]),.I2(r1_2[22:22]),.I3(r1_2[23:23]),.O(un33_s_count_a_5_0_axb_23));
defparam un33_s_count_a_5_0_axb_23_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_24_cZ(.I0(r1[22:22]),.I1(r1[23:23]),.I2(r1_2[23:23]),.I3(r1_2[24:24]),.O(un33_s_count_a_5_0_axb_24));
defparam un33_s_count_a_5_0_axb_24_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_25_cZ(.I0(r1[23:23]),.I1(r1[24:24]),.I2(r1_2[24:24]),.I3(r1_2[25:25]),.O(un33_s_count_a_5_0_axb_25));
defparam un33_s_count_a_5_0_axb_25_cZ.INIT=16'hC639;
  LUT4 un33_s_count_a_5_0_axb_27_cZ(.I0(r1[25:25]),.I1(r1_2[26:26]),.I2(r1_2[27:27]),.I3(s_rad_i[27:27]),.O(un33_s_count_a_5_0_axb_27));
defparam un33_s_count_a_5_0_axb_27_cZ.INIT=16'h2DD2;
  LUT4 desc2703(.I0(r1_2[27:27]),.I1(r1_2[28:28]),.I2(s_rad_i[27:27]),.I3(s_rad_i[28:28]),.O(un33_s_count_a_5_0_axb_28));
defparam desc2703.INIT=16'hC639;
  LUT4 desc2704(.I0(r1_2[28:28]),.I1(r1_2[29:29]),.I2(s_rad_i[28:28]),.I3(s_rad_i[29:29]),.O(un33_s_count_a_5_0_axb_29));
defparam desc2704.INIT=16'hC639;
  LUT4 desc2705(.I0(r1_2[29:29]),.I1(r1_2[30:30]),.I2(s_rad_i[29:29]),.I3(s_rad_i[30:30]),.O(un33_s_count_a_5_0_axb_30));
defparam desc2705.INIT=16'hC639;
  LUT4 desc2706(.I0(r1_2[30:30]),.I1(r1_2[31:31]),.I2(s_rad_i[30:30]),.I3(s_rad_i[31:31]),.O(un33_s_count_a_5_0_axb_31));
defparam desc2706.INIT=16'hC639;
  LUT4 desc2707(.I0(r1_2[31:31]),.I1(r1_2[32:32]),.I2(s_rad_i[31:31]),.I3(s_rad_i[32:32]),.O(un33_s_count_a_5_0_axb_32));
defparam desc2707.INIT=16'hC639;
  LUT4 desc2708(.I0(r1_2[32:32]),.I1(r1_2[33:33]),.I2(s_rad_i[32:32]),.I3(s_rad_i[33:33]),.O(un33_s_count_a_5_0_axb_33));
defparam desc2708.INIT=16'hC639;
  LUT4 desc2709(.I0(r1_2[33:33]),.I1(r1_2[34:34]),.I2(s_rad_i[33:33]),.I3(s_rad_i[34:34]),.O(un33_s_count_a_5_0_axb_34));
defparam desc2709.INIT=16'hC639;
  LUT4 desc2710(.I0(r1_2[34:34]),.I1(r1_2[35:35]),.I2(s_rad_i[34:34]),.I3(s_rad_i[35:35]),.O(un33_s_count_a_5_0_axb_35));
defparam desc2710.INIT=16'hC639;
  LUT4 desc2711(.I0(r1_2[35:35]),.I1(r1_2[36:36]),.I2(s_rad_i[35:35]),.I3(s_rad_i[36:36]),.O(un33_s_count_a_5_0_axb_36));
defparam desc2711.INIT=16'hC639;
  LUT4 desc2712(.I0(r1_2[36:36]),.I1(r1_2[37:37]),.I2(s_rad_i[36:36]),.I3(s_rad_i[37:37]),.O(un33_s_count_a_5_0_axb_37));
defparam desc2712.INIT=16'hC639;
  LUT4 desc2713(.I0(r1_2[37:37]),.I1(r1_2[38:38]),.I2(s_rad_i[37:37]),.I3(s_rad_i[38:38]),.O(un33_s_count_a_5_0_axb_38));
defparam desc2713.INIT=16'hC639;
  LUT4 desc2714(.I0(r1_2[38:38]),.I1(r1_2[39:39]),.I2(s_rad_i[38:38]),.I3(s_rad_i[39:39]),.O(un33_s_count_a_5_0_axb_39));
defparam desc2714.INIT=16'hC639;
  LUT4 desc2715(.I0(r1_2[39:39]),.I1(r1_2[40:40]),.I2(s_rad_i[39:39]),.I3(s_rad_i[40:40]),.O(un33_s_count_a_5_0_axb_40));
defparam desc2715.INIT=16'hC639;
  LUT4 desc2716(.I0(r1_2[40:40]),.I1(r1_2[41:41]),.I2(s_rad_i[40:40]),.I3(s_rad_i[41:41]),.O(un33_s_count_a_5_0_axb_41));
defparam desc2716.INIT=16'hC639;
  LUT4 desc2717(.I0(r1_2[41:41]),.I1(r1_2[42:42]),.I2(s_rad_i[41:41]),.I3(s_rad_i[42:42]),.O(un33_s_count_a_5_0_axb_42));
defparam desc2717.INIT=16'hC639;
  LUT4 desc2718(.I0(r1_2[42:42]),.I1(r1_2[43:43]),.I2(s_rad_i[42:42]),.I3(s_rad_i[43:43]),.O(un33_s_count_a_5_0_axb_43));
defparam desc2718.INIT=16'hC639;
  LUT4 desc2719(.I0(r1_2[43:43]),.I1(r1_2[44:44]),.I2(s_rad_i[43:43]),.I3(s_rad_i[44:44]),.O(un33_s_count_a_5_0_axb_44));
defparam desc2719.INIT=16'hC639;
  LUT4 desc2720(.I0(r1_2[44:44]),.I1(r1_2[45:45]),.I2(s_rad_i[44:44]),.I3(s_rad_i[45:45]),.O(un33_s_count_a_5_0_axb_45));
defparam desc2720.INIT=16'hC639;
  LUT4 desc2721(.I0(r1_2[45:45]),.I1(r1_2[46:46]),.I2(s_rad_i[45:45]),.I3(s_rad_i[46:46]),.O(un33_s_count_a_5_0_axb_46));
defparam desc2721.INIT=16'hC639;
  LUT4 desc2722(.I0(r1_2[46:46]),.I1(r1_2[47:47]),.I2(s_rad_i[46:46]),.I3(s_rad_i[47:47]),.O(un33_s_count_a_5_0_axb_47));
defparam desc2722.INIT=16'hC639;
  LUT4 desc2723(.I0(r1_2[47:47]),.I1(r1_2[48:48]),.I2(s_rad_i[47:47]),.I3(s_rad_i[48:48]),.O(un33_s_count_a_5_0_axb_48));
defparam desc2723.INIT=16'hC639;
  LUT4 desc2724(.I0(r1_2[48:48]),.I1(r1_2[49:49]),.I2(s_rad_i[48:48]),.I3(s_rad_i[49:49]),.O(un33_s_count_a_5_0_axb_49));
defparam desc2724.INIT=16'hC639;
  LUT4 desc2725(.I0(r1_2[49:49]),.I1(r1_2[50:50]),.I2(s_rad_i[49:49]),.I3(s_rad_i[50:50]),.O(un33_s_count_a_5_0_axb_50));
defparam desc2725.INIT=16'hC639;
  LUT3 v_r1_3_axb_0_cZ(.I0(b[0:0]),.I1(r0[0:0]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_0));
defparam v_r1_3_axb_0_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_1_cZ(.I0(b[1:1]),.I1(r0[1:1]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_1));
defparam v_r1_3_axb_1_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_2_cZ(.I0(b[2:2]),.I1(r0[2:2]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_2));
defparam v_r1_3_axb_2_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_3_cZ(.I0(b[3:3]),.I1(r0[3:3]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_3));
defparam v_r1_3_axb_3_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_4_cZ(.I0(b[4:4]),.I1(r0[4:4]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_4));
defparam v_r1_3_axb_4_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_5_cZ(.I0(b[5:5]),.I1(r0[5:5]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_5));
defparam v_r1_3_axb_5_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_6_cZ(.I0(b[6:6]),.I1(r0[6:6]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_6));
defparam v_r1_3_axb_6_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_7_cZ(.I0(b[7:7]),.I1(r0[7:7]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_7));
defparam v_r1_3_axb_7_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_8_cZ(.I0(b[8:8]),.I1(r0[8:8]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_8));
defparam v_r1_3_axb_8_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_9_cZ(.I0(b[9:9]),.I1(r0[9:9]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_9));
defparam v_r1_3_axb_9_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_10_cZ(.I0(b[10:10]),.I1(r0[10:10]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_10));
defparam v_r1_3_axb_10_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_11_cZ(.I0(b[11:11]),.I1(r0[11:11]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_11));
defparam v_r1_3_axb_11_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_12_cZ(.I0(b[12:12]),.I1(r0[12:12]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_12));
defparam v_r1_3_axb_12_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_13_cZ(.I0(b[13:13]),.I1(r0[13:13]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_13));
defparam v_r1_3_axb_13_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_14_cZ(.I0(b[14:14]),.I1(r0[14:14]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_14));
defparam v_r1_3_axb_14_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_15_cZ(.I0(b[15:15]),.I1(r0[15:15]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_15));
defparam v_r1_3_axb_15_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_16_cZ(.I0(b[16:16]),.I1(r0[16:16]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_16));
defparam v_r1_3_axb_16_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_17_cZ(.I0(b[17:17]),.I1(r0[17:17]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_17));
defparam v_r1_3_axb_17_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_18_cZ(.I0(b[18:18]),.I1(r0[18:18]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_18));
defparam v_r1_3_axb_18_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_19_cZ(.I0(b[19:19]),.I1(r0[19:19]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_19));
defparam v_r1_3_axb_19_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_20_cZ(.I0(b[20:20]),.I1(r0[20:20]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_20));
defparam v_r1_3_axb_20_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_21_cZ(.I0(b[21:21]),.I1(r0[21:21]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_21));
defparam v_r1_3_axb_21_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_22_cZ(.I0(b[22:22]),.I1(r0[22:22]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_22));
defparam v_r1_3_axb_22_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_23_cZ(.I0(b[23:23]),.I1(r0[23:23]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_23));
defparam v_r1_3_axb_23_cZ.INIT=8'h96;
  LUT3 v_r1_3_axb_24_cZ(.I0(b[24:24]),.I1(r0[24:24]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_24));
defparam v_r1_3_axb_24_cZ.INIT=8'h96;
  LUT2 v_r1_2_3_cZ(.I0(b_2[0:0]),.I1(r0_2[0:0]),.O(v_r1_2_3_scalar));
defparam v_r1_2_3_cZ.INIT=4'h6;
  LUT2 un31_s_count_0_N_3_i_cZ(.I0(r1_2[51:51]),.I1(s_rad_i[51:51]),.O(un31_s_count_0_N_3_i));
defparam un31_s_count_0_N_3_i_cZ.INIT=4'h9;
  FD s_ine_o_Z(.Q(s_ine_o),.D(s_ine_o_0),.C(clk_i));
  FDE desc2726(.Q(r1_2[0:0]),.D(v_r1_2_3[0:0]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2727(.Q(r1_2[1:1]),.D(v_r1_2_3[1:1]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2728(.Q(r1_2[2:2]),.D(v_r1_2_3[2:2]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2729(.Q(r1_2[3:3]),.D(v_r1_2_3[3:3]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2730(.Q(r1_2[4:4]),.D(v_r1_2_3[4:4]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2731(.Q(r1_2[5:5]),.D(v_r1_2_3[5:5]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2732(.Q(r1_2[6:6]),.D(v_r1_2_3[6:6]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2733(.Q(r1_2[7:7]),.D(v_r1_2_3[7:7]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2734(.Q(r1_2[8:8]),.D(v_r1_2_3[8:8]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2735(.Q(r1_2[9:9]),.D(v_r1_2_3[9:9]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2736(.Q(r1_2[10:10]),.D(v_r1_2_3[10:10]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2737(.Q(r1_2[11:11]),.D(v_r1_2_3[11:11]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2738(.Q(r1_2[12:12]),.D(v_r1_2_3[12:12]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2739(.Q(r1_2[13:13]),.D(v_r1_2_3[13:13]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2740(.Q(r1_2[14:14]),.D(v_r1_2_3[14:14]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2741(.Q(r1_2[15:15]),.D(v_r1_2_3[15:15]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2742(.Q(r1_2[16:16]),.D(v_r1_2_3[16:16]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2743(.Q(r1_2[17:17]),.D(v_r1_2_3[17:17]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2744(.Q(r1_2[18:18]),.D(v_r1_2_3[18:18]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2745(.Q(r1_2[19:19]),.D(v_r1_2_3[19:19]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2746(.Q(r1_2[20:20]),.D(v_r1_2_3[20:20]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2747(.Q(r1_2[21:21]),.D(v_r1_2_3[21:21]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2748(.Q(r1_2[22:22]),.D(v_r1_2_3[22:22]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2749(.Q(r1_2[23:23]),.D(v_r1_2_3[23:23]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2750(.Q(r1_2[24:24]),.D(v_r1_2_3[24:24]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2751(.Q(r1_2[25:25]),.D(v_r1_2_3[25:25]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2752(.Q(r1_2[26:26]),.D(v_r1_2_3[26:26]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2753(.Q(r1_2[27:27]),.D(v_r1_2_3[27:27]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2754(.Q(r1_2[28:28]),.D(v_r1_2_3[28:28]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2755(.Q(r1_2[29:29]),.D(v_r1_2_3[29:29]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2756(.Q(r1_2[30:30]),.D(v_r1_2_3[30:30]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2757(.Q(r1_2[31:31]),.D(v_r1_2_3[31:31]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2758(.Q(r1_2[32:32]),.D(v_r1_2_3[32:32]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2759(.Q(r1_2[33:33]),.D(v_r1_2_3[33:33]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2760(.Q(r1_2[34:34]),.D(v_r1_2_3[34:34]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2761(.Q(r1_2[35:35]),.D(v_r1_2_3[35:35]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2762(.Q(r1_2[36:36]),.D(v_r1_2_3[36:36]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2763(.Q(r1_2[37:37]),.D(v_r1_2_3[37:37]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2764(.Q(r1_2[38:38]),.D(v_r1_2_3[38:38]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2765(.Q(r1_2[39:39]),.D(v_r1_2_3[39:39]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2766(.Q(r1_2[40:40]),.D(v_r1_2_3[40:40]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2767(.Q(r1_2[41:41]),.D(v_r1_2_3[41:41]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2768(.Q(r1_2[42:42]),.D(v_r1_2_3[42:42]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2769(.Q(r1_2[43:43]),.D(v_r1_2_3[43:43]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2770(.Q(r1_2[44:44]),.D(v_r1_2_3[44:44]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2771(.Q(r1_2[45:45]),.D(v_r1_2_3[45:45]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2772(.Q(r1_2[46:46]),.D(v_r1_2_3[46:46]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2773(.Q(r1_2[47:47]),.D(v_r1_2_3[47:47]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2774(.Q(r1_2[48:48]),.D(v_r1_2_3[48:48]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2775(.Q(r1_2[49:49]),.D(v_r1_2_3[49:49]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2776(.Q(r1_2[50:50]),.D(v_r1_2_3[50:50]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2777(.Q(r1_2[51:51]),.D(v_r1_2_3[51:51]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2778(.Q(r1[0:0]),.D(v_r1_3[0:0]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2779(.Q(r1[1:1]),.D(v_r1_3[1:1]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2780(.Q(r1[2:2]),.D(v_r1_3[2:2]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2781(.Q(r1[3:3]),.D(v_r1_3[3:3]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2782(.Q(r1[4:4]),.D(v_r1_3[4:4]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2783(.Q(r1[5:5]),.D(v_r1_3[5:5]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2784(.Q(r1[6:6]),.D(v_r1_3[6:6]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2785(.Q(r1[7:7]),.D(v_r1_3[7:7]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2786(.Q(r1[8:8]),.D(v_r1_3[8:8]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2787(.Q(r1[9:9]),.D(v_r1_3[9:9]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2788(.Q(r1[10:10]),.D(v_r1_3[10:10]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2789(.Q(r1[11:11]),.D(v_r1_3[11:11]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2790(.Q(r1[12:12]),.D(v_r1_3[12:12]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2791(.Q(r1[13:13]),.D(v_r1_3[13:13]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2792(.Q(r1[14:14]),.D(v_r1_3[14:14]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2793(.Q(r1[15:15]),.D(v_r1_3[15:15]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2794(.Q(r1[16:16]),.D(v_r1_3[16:16]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2795(.Q(r1[17:17]),.D(v_r1_3[17:17]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2796(.Q(r1[18:18]),.D(v_r1_3[18:18]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2797(.Q(r1[19:19]),.D(v_r1_3[19:19]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2798(.Q(r1[20:20]),.D(v_r1_3[20:20]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2799(.Q(r1[21:21]),.D(v_r1_3[21:21]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2800(.Q(r1[22:22]),.D(v_r1_3[22:22]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2801(.Q(r1[23:23]),.D(v_r1_3[23:23]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2802(.Q(r1[24:24]),.D(v_r1_3[24:24]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FDE desc2803(.Q(r1[25:25]),.D(v_r1_3[25:25]),.C(clk_i),.CE(un12_s_state_0_a2_lut6_2_O6));
  FD desc2804(.Q(sqrt_sqr_o[12:12]),.D(s_sqr_o[12:12]),.C(clk_i));
  FD desc2805(.Q(sqrt_sqr_o[13:13]),.D(s_sqr_o[13:13]),.C(clk_i));
  FD desc2806(.Q(sqrt_sqr_o[14:14]),.D(s_sqr_o[14:14]),.C(clk_i));
  FD desc2807(.Q(sqrt_sqr_o[15:15]),.D(s_sqr_o[15:15]),.C(clk_i));
  FD desc2808(.Q(sqrt_sqr_o[16:16]),.D(s_sqr_o[16:16]),.C(clk_i));
  FD desc2809(.Q(sqrt_sqr_o[17:17]),.D(s_sqr_o[17:17]),.C(clk_i));
  FD desc2810(.Q(sqrt_sqr_o[18:18]),.D(s_sqr_o[18:18]),.C(clk_i));
  FD desc2811(.Q(sqrt_sqr_o[19:19]),.D(s_sqr_o[19:19]),.C(clk_i));
  FD desc2812(.Q(sqrt_sqr_o[20:20]),.D(s_sqr_o[20:20]),.C(clk_i));
  FD desc2813(.Q(sqrt_sqr_o[21:21]),.D(s_sqr_o[21:21]),.C(clk_i));
  FD desc2814(.Q(sqrt_sqr_o[22:22]),.D(s_sqr_o[22:22]),.C(clk_i));
  FD desc2815(.Q(sqrt_sqr_o[23:23]),.D(s_sqr_o[23:23]),.C(clk_i));
  FD desc2816(.Q(sqrt_sqr_o[24:24]),.D(s_sqr_o[24:24]),.C(clk_i));
  FD desc2817(.Q(sqrt_sqr_o[0:0]),.D(s_sqr_o[0:0]),.C(clk_i));
  FD desc2818(.Q(sqrt_sqr_o[1:1]),.D(s_sqr_o[1:1]),.C(clk_i));
  FD desc2819(.Q(sqrt_sqr_o[2:2]),.D(s_sqr_o[2:2]),.C(clk_i));
  FD desc2820(.Q(sqrt_sqr_o[3:3]),.D(s_sqr_o[3:3]),.C(clk_i));
  FD desc2821(.Q(sqrt_sqr_o[4:4]),.D(s_sqr_o[4:4]),.C(clk_i));
  FD desc2822(.Q(sqrt_sqr_o[5:5]),.D(s_sqr_o[5:5]),.C(clk_i));
  FD desc2823(.Q(sqrt_sqr_o[6:6]),.D(s_sqr_o[6:6]),.C(clk_i));
  FD desc2824(.Q(sqrt_sqr_o[7:7]),.D(s_sqr_o[7:7]),.C(clk_i));
  FD desc2825(.Q(sqrt_sqr_o[8:8]),.D(s_sqr_o[8:8]),.C(clk_i));
  FD desc2826(.Q(sqrt_sqr_o[9:9]),.D(s_sqr_o[9:9]),.C(clk_i));
  FD desc2827(.Q(sqrt_sqr_o[10:10]),.D(s_sqr_o[10:10]),.C(clk_i));
  FD desc2828(.Q(sqrt_sqr_o[11:11]),.D(s_sqr_o[11:11]),.C(clk_i));
  FD desc2829(.Q(s_rad_i[41:41]),.D(pre_norm_sqrt_fracta_o_14),.C(clk_i));
  FD desc2830(.Q(s_rad_i[42:42]),.D(pre_norm_sqrt_fracta_o_15),.C(clk_i));
  FD desc2831(.Q(s_rad_i[43:43]),.D(pre_norm_sqrt_fracta_o_16),.C(clk_i));
  FD desc2832(.Q(s_rad_i[44:44]),.D(pre_norm_sqrt_fracta_o_17),.C(clk_i));
  FD desc2833(.Q(s_rad_i[45:45]),.D(pre_norm_sqrt_fracta_o_18),.C(clk_i));
  FD desc2834(.Q(s_rad_i[46:46]),.D(pre_norm_sqrt_fracta_o_19),.C(clk_i));
  FD desc2835(.Q(s_rad_i[47:47]),.D(pre_norm_sqrt_fracta_o_20),.C(clk_i));
  FD desc2836(.Q(s_rad_i[48:48]),.D(pre_norm_sqrt_fracta_o_21),.C(clk_i));
  FD desc2837(.Q(s_rad_i[49:49]),.D(pre_norm_sqrt_fracta_o_22),.C(clk_i));
  FD desc2838(.Q(s_rad_i[50:50]),.D(pre_norm_sqrt_fracta_o_23),.C(clk_i));
  FD desc2839(.Q(s_rad_i[51:51]),.D(pre_norm_sqrt_fracta_o_0[51:51]),.C(clk_i));
  FD desc2840(.Q(s_rad_i[27:27]),.D(pre_norm_sqrt_fracta_o_0_d0),.C(clk_i));
  FD desc2841(.Q(s_rad_i[28:28]),.D(pre_norm_sqrt_fracta_o_1),.C(clk_i));
  FD desc2842(.Q(s_rad_i[34:34]),.D(pre_norm_sqrt_fracta_o_7),.C(clk_i));
  FD desc2843(.Q(s_rad_i[35:35]),.D(pre_norm_sqrt_fracta_o_8),.C(clk_i));
  FD desc2844(.Q(s_rad_i[36:36]),.D(pre_norm_sqrt_fracta_o_9),.C(clk_i));
  FD desc2845(.Q(s_rad_i[37:37]),.D(pre_norm_sqrt_fracta_o_10),.C(clk_i));
  FD desc2846(.Q(s_rad_i[38:38]),.D(pre_norm_sqrt_fracta_o_11),.C(clk_i));
  FD desc2847(.Q(s_rad_i[39:39]),.D(pre_norm_sqrt_fracta_o_12),.C(clk_i));
  FD desc2848(.Q(s_rad_i[40:40]),.D(pre_norm_sqrt_fracta_o_13),.C(clk_i));
  FD s_start_i_Z(.Q(s_start_i),.D(s_start_i_0),.C(clk_i));
  FD desc2849(.Q(b_2[50:50]),.D(s_start_i),.C(clk_i));
  FD ine_o_Z(.Q(sqrt_ine_o),.D(s_ine_o),.C(clk_i));
  MUXCY un31_s_count_0_I_139_cZ(.DI(GND),.CI(un31_s_count_0_data_tmp[16:16]),.S(un31_s_count_0_N_3_i),.O(un31_s_count_0_I_139));
  MUXCY desc2850(.DI(un14_s_state_lt50),.CI(un14_s_state_cry[48:48]),.S(un14_s_state_df50),.O(un14_s_state_cry[50:50]));
  MUXCY desc2851(.DI(un27_s_count_lt50),.CI(un27_s_count_cry[48:48]),.S(un27_s_count_df50),.O(un27_s_count_cry[50:50]));
  MUXF7 desc2852(.I0(g0_5i0),.I1(g0_5i1),.S(r0_2[14:14]),.O(v_r1_2_3_56_0_tz));
  LUT5 desc2853(.I0(b_2[14:14]),.I1(r0_2[13:13]),.I2(r0_2[16:16]),.I3(r0_2[15:15]),.I4(v_r1_2_3_35_0_RNIKOE74),.O(g0_5i1));
defparam desc2853.INIT=32'hFEF0FAF0;
  LUT6 desc2854(.I0(b_2[14:14]),.I1(r0_2[13:13]),.I2(r0_2[16:16]),.I3(r0_2[15:15]),.I4(g3),.I5(v_r1_2_3_42_0),.O(g0_5i0));
defparam desc2854.INIT=64'hF8F0F8F0F8F0F0F0;
  LUT3_L v_r1_2_3_72_0_N_2L1_cZ(.I0(r0_2[20:20]),.I1(r0_2[19:19]),.I2(v_r1_2_3_63_2),.LO(v_r1_2_3_72_0_N_2L1));
defparam v_r1_2_3_72_0_N_2L1_cZ.INIT=8'h7F;
  LUT2_L desc2855(.I0(r0_2[11:11]),.I1(b_2_RNIMF314[10:10]),.LO(r0_2_RNI351G4[11:11]));
defparam desc2855.INIT=4'h7;
  LUT6 desc2856(.I0(b_2[12:12]),.I1(r0_2[12:12]),.I2(r0_2[14:14]),.I3(r0_2[13:13]),.I4(g2_0),.I5(r0_2_RNI351G4[11:11]),.O(v_r1_2_3_49_0_tz));
defparam desc2856.INIT=64'hFAF0F8F0FEF0FCF0;
  LUT5 desc2857(.I0(b_2[22:22]),.I1(r0_2[22:22]),.I2(c[4:4]),.I3(m73_lut6_2_O6),.I4(m45),.O(b_2_RNI46VUE[22:22]));
defparam desc2857.INIT=32'h96669969;
  LUT5_L desc2858(.I0(b_2[18:18]),.I1(r0_2[20:20]),.I2(r0_2[19:19]),.I3(r0_2[18:18]),.I4(b_2_RNIRH7KV[16:16]),.LO(b_2_RNI5B6111[18:18]));
defparam desc2858.INIT=32'h13331313;
  LUT6 desc2859(.I0(b_2[20:20]),.I1(r0_2[21:21]),.I2(b_2_RNI46VUE[22:22]),.I3(v_r1_2_3_28),.I4(v_r1_2_3_65_c),.I5(b_2_RNI5B6111[18:18]),.O(v_r1_2_3_0_axb_22));
defparam desc2859.INIT=64'hC387C30FC387C387;
  LUT5 desc2860(.I0(b_2[14:14]),.I1(r0_2[16:16]),.I2(r0_2[15:15]),.I3(v_r1_2_3_49_0_tz),.I4(N_4),.O(b_2_RNIT9A1G_0[14:14]));
defparam desc2860.INIT=32'h00007FFF;
  LUT4_L desc2861(.I0(b_2[16:16]),.I1(r0_2[17:17]),.I2(b_2_RNIT9A1G_0[14:14]),.I3(v_r1_2_3_56_0_tz),.LO(b_2_RNIRH7KV[16:16]));
defparam desc2861.INIT=16'h73F3;
  LUT4 v_r1_2_3_73_0_lut6_2_RNIM5CP22_cZ(.I0(v_r1_2_3_73_0_lut6_2_O5),.I1(r0_2_RNIM65S1[23:23]),.I2(g4_0),.I3(v_r1_2_3_65_c),.O(v_r1_2_3_73_0_lut6_2_RNIM5CP22));
defparam v_r1_2_3_73_0_lut6_2_RNIM5CP22_cZ.INIT=16'hBBB8;
  LUT6 desc2862(.I0(r0_2[23:23]),.I1(b_2[22:22]),.I2(r0_2[22:22]),.I3(b_2[20:20]),.I4(r0_2[21:21]),.I5(r0_2[20:20]),.O(r0_2_RNIM65S1[23:23]));
defparam desc2862.INIT=64'hFFD7FFFFD7FFFFFF;
  LUT5 desc2863(.I0(b_2[20:20]),.I1(r0_2[20:20]),.I2(r0_2_RNI9011F_O6[22:22]),.I3(g1_0),.I4(v_r1_2_3_65_c),.O(v_r1_2_3_0_axb_21));
defparam desc2863.INIT=32'hE1E1E187;
  LUT4_L desc2864(.I0(b_2[16:16]),.I1(r0_2_RNIMOCU9[14:14]),.I2(g0_0_0_0),.I3(N_4),.LO(g4_0_0_0));
defparam desc2864.INIT=16'hFFA8;
  LUT5 desc2865(.I0(r0_2[14:14]),.I1(r0_2[13:13]),.I2(g1_0_0_2),.I3(g3),.I4(v_r1_2_3_42_0),.O(r0_2_RNIMOCU9[14:14]));
defparam desc2865.INIT=32'hE0E0E0A0;
  LUT4 v_r1_2_3_21_2_RNIMLGQ_cZ(.I0(b_2[8:8]),.I1(r0_2[8:8]),.I2(r0_2[7:7]),.I3(v_r1_2_3_21_2),.O(v_r1_2_3_21_2_RNIMLGQ));
defparam v_r1_2_3_21_2_RNIMLGQ_cZ.INIT=16'hE888;
  LUT5 desc2866(.I0(b_2[20:20]),.I1(r0_2[20:20]),.I2(g0_0_2),.I3(g4_1),.I4(v_r1_2_3_65_c),.O(v_r1_2_3_31));
defparam desc2866.INIT=32'hE0E0E080;
  LUT5 v_r1_2_3_0_cry_9_RNO_cZ(.I0(b_2[8:8]),.I1(r0_2[8:8]),.I2(r0_2[7:7]),.I3(r0_2[9:9]),.I4(v_r1_2_3_21_2),.O(v_r1_2_3_0_cry_9_RNO));
defparam v_r1_2_3_0_cry_9_RNO_cZ.INIT=32'h17E87788;
  FDR desc2867(.Q(b_2_fast),.D(b_2[2:2]),.C(clk_i),.R(s_start_i));
  FDRE desc2868(.Q(r0_2_fast[1:1]),.D(v_r1_2_3[1:1]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc2869(.Q(r0_2_fast[0:0]),.D(v_r1_2_3[0:0]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  LUT6 desc2870(.I0(r0_2[19:19]),.I1(r0_2[18:18]),.I2(b_2[16:16]),.I3(r0_2[17:17]),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_65_c));
defparam desc2870.INIT=64'h8800800088000000;
  LUT5 desc2871(.I0(r0_2[14:14]),.I1(r0_2[13:13]),.I2(r0_2[16:16]),.I3(r0_2[15:15]),.I4(v_r1_2_3_35_0_RNIKOE74),.O(N_4));
defparam desc2871.INIT=32'h80000000;
  LUT6 desc2872(.I0(r0_2[20:20]),.I1(b_2[16:16]),.I2(r0_2[17:17]),.I3(g0_6_0),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.O(g5_0));
defparam desc2872.INIT=64'hFAAAEAAAFAAAAAAA;
  LUT6 desc2873(.I0(r0_2[18:18]),.I1(r0_2[17:17]),.I2(g1_0_0_1),.I3(g1_1_1),.I4(v_r1_2_3_49_0_tz),.I5(g4_0_0_0),.O(g1_0));
defparam desc2873.INIT=64'hE0E0E0E0E0A0A0A0;
  LUT2 desc2874(.I0(r0_2[20:20]),.I1(g1_0),.O(v_r1_2_3_65_0_0));
defparam desc2874.INIT=4'hE;
  LUT6 v_r1_2_3_72_0_N_2L1_RNIMAAJ42(.I0(r0_2[22:22]),.I1(b_2[20:20]),.I2(r0_2[21:21]),.I3(g5_0),.I4(g1_0),.I5(v_r1_2_3_72_0_N_2L1),.O(v_r1_2_3_77_0_tz));
defparam v_r1_2_3_72_0_N_2L1_RNIMAAJ42.INIT=64'hEAEAEAAAFAFAFAFA;
  LUT6 v_r1_2_3_13_RNIHH162(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(g0_0_a4_3),.I4(v_r1_2_3_4),.I5(v_r1_2_3_14_0),.O(N_5_0_0));
defparam v_r1_2_3_13_RNIHH162.INIT=64'hF800F800F8008800;
  LUT6 desc2875(.I0(b_2[10:10]),.I1(b_2[8:8]),.I2(r0_2[10:10]),.I3(r0_2[9:9]),.I4(N_5_0_0),.I5(v_r1_2_3_28_0_tz),.O(b_2_RNIMF314[10:10]));
defparam desc2875.INIT=64'hFFFFE8A0FFFFA0A0;
  LUT3 desc2876(.I0(r0_2[12:12]),.I1(r0_2[11:11]),.I2(b_2_RNIMF314[10:10]),.O(g3));
defparam desc2876.INIT=8'h80;
  LUT6 v_r1_2_3_35_0_RNI0PKK2(.I0(b_2[12:12]),.I1(r0_2[12:12]),.I2(r0_2[11:11]),.I3(g4_0_0_1),.I4(v_r1_2_3_35_0),.I5(v_r1_2_3_21_2_RNIMLGQ),.O(v_r1_2_3_42_0));
defparam v_r1_2_3_35_0_RNI0PKK2.INIT=64'hA8A8A888A8A88888;
  LUT2 v_r1_2_3_35_RNO_0(.I0(r0_2[8:8]),.I1(r0_2[7:7]),.O(g0_i_0));
defparam v_r1_2_3_35_RNO_0.INIT=4'h8;
  LUT2_L desc2877(.I0(b_2[10:10]),.I1(r0_2[10:10]),.LO(N_4_1));
defparam desc2877.INIT=4'hE;
  LUT6 desc2878(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[8:8]),.I3(r0_2[7:7]),.I4(r0_2[9:9]),.I5(N_4_1),.O(g0_0_a4_3));
defparam desc2878.INIT=64'hE000000000000000;
  LUT6 v_r1_2_3_35_0_RNO(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(g0_i_0),.I4(v_r1_2_3_4),.I5(v_r1_2_3_14_0),.O(v_r1_2_3_10));
defparam v_r1_2_3_35_0_RNO.INIT=64'hE800E800E8008800;
  LUT6 desc2879(.I0(b_2[18:18]),.I1(b_2[14:14]),.I2(r0_2[18:18]),.I3(r0_2[16:16]),.I4(r0_2[15:15]),.I5(v_r1_2_3_49_0_tz),.O(g0_i_a3_0));
defparam desc2879.INIT=64'hECA0A0A0A0A0A0A0;
  LUT6 v_r1_2_3_35_0_RNIKOE74_cZ(.I0(b_2[12:12]),.I1(r0_2[12:12]),.I2(r0_2[11:11]),.I3(g0_0_a4_0_2),.I4(v_r1_2_3_35_0),.I5(v_r1_2_3_21_2_RNIMLGQ),.O(v_r1_2_3_35_0_RNIKOE74));
defparam v_r1_2_3_35_0_RNIKOE74_cZ.INIT=64'hE8E8E888E8E88888;
  LUT6 desc2880(.I0(b_2[14:14]),.I1(r0_2[16:16]),.I2(r0_2[15:15]),.I3(g0_0_a3_0_2),.I4(v_r1_2_3_35_0_RNIKOE74),.I5(v_r1_2_3_49_0_tz),.O(v_r1_2_3_22));
defparam desc2880.INIT=64'hFF808080FF000000;
  LUT6 v_r1_2_3_59_0_lut6_2_RNII8ONV(.I0(b_2[16:16]),.I1(g0_i_1),.I2(g0_0_a3_0_2),.I3(v_r1_2_3_35_0_RNIKOE74),.I4(g0_i_a3_0),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_28));
defparam v_r1_2_3_59_0_lut6_2_RNII8ONV.INIT=64'hCCCCC888CCCCC000;
  LUT2 v_r1_2_3_0_cry_16_RNO_0(.I0(r0_2[14:14]),.I1(r0_2[13:13]),.O(v_r1_2_3_48_0));
defparam v_r1_2_3_0_cry_16_RNO_0.INIT=4'h8;
  LUT3 v_r1_2_3_21_2_RNIJUQF(.I0(r0_2[8:8]),.I1(r0_2[7:7]),.I2(v_r1_2_3_21_2),.O(N_4_0));
defparam v_r1_2_3_21_2_RNIJUQF.INIT=8'h80;
  LUT6 v_r1_2_3_35_0_RNIM6633(.I0(b_2[8:8]),.I1(r0_2[11:11]),.I2(g4_0_2),.I3(v_r1_2_3_28_0_tz),.I4(N_4_0),.I5(v_r1_2_3_35_0),.O(g2_0));
defparam v_r1_2_3_35_0_RNIM6633.INIT=64'hCCCCCCCCC0C08000;
  LUT5 desc2881(.I0(r0_2[14:14]),.I1(r0_2[13:13]),.I2(r0_2[16:16]),.I3(r0_2[15:15]),.I4(v_r1_2_3_35_0_RNIKOE74),.O(g0_0_0_0));
defparam desc2881.INIT=32'hF8F0F0F0;
  LUT5 desc2882(.I0(b_2[14:14]),.I1(r0_2[16:16]),.I2(r0_2[15:15]),.I3(v_r1_2_3_49_0_tz),.I4(N_4),.O(g2_1_0));
defparam desc2882.INIT=32'hFFFF8000;
  LUT6 desc2883(.I0(r0_2[18:18]),.I1(b_2[16:16]),.I2(r0_2[17:17]),.I3(g4_0_1),.I4(g2_1_0),.I5(v_r1_2_3_56_0_tz),.O(g4_1));
defparam desc2883.INIT=64'hFA00EA00FA00AA00;
  LUT5 desc2884(.I0(r0_2[14:14]),.I1(b_2[14:14]),.I2(r0_2[13:13]),.I3(v_r1_2_3_35_0_RNIKOE74),.I4(v_r1_2_3_49_0_tz),.O(N_6_1_0));
defparam desc2884.INIT=32'hECCCA000;
  LUT6 v_r1_2_3_52_0_lut6_2_RNIU7M301(.I0(r0_2[18:18]),.I1(g4_0_0),.I2(g0_0_a4_0),.I3(g0_0_a4_0_1),.I4(N_6_1_0),.I5(v_r1_2_3_56_0_tz),.O(g4_0));
defparam v_r1_2_3_52_0_lut6_2_RNIU7M301.INIT=64'hCCC8C8C8CC888888;
  LUT6 v_r1_2_3_14_RNI66FT(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(r0_2[8:8]),.I4(r0_2[7:7]),.I5(v_r1_2_3_14),.O(v_r1_2_3_28_0_tz));
defparam v_r1_2_3_14_RNI66FT.INIT=64'hFFE8FF00FF88FF00;
  LUT6 desc2885(.I0(r0[25:25]),.I1(c[1:1]),.I2(c[2:2]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(N_84_0),.O(N_89_0));
defparam desc2885.INIT=64'hF7FFF8F0070F0800;
  LUT6 desc2886(.I0(r0[25:25]),.I1(c[1:1]),.I2(c[2:2]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(N_10_1),.O(N_12_1));
defparam desc2886.INIT=64'hDFFFE0C01F3F2000;
  LUT6 desc2887(.I0(r0[13:13]),.I1(r0[14:14]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m24_lut6_2_O6),.O(N_90_0));
defparam desc2887.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2888(.I0(r0[12:12]),.I1(r0[11:11]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m32),.O(m36));
defparam desc2888.INIT=64'h3F5FCFAF3050C0A0;
  LUT6 desc2889(.I0(r0[19:19]),.I1(r0[18:18]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m17_lut6_2_O5),.O(m157));
defparam desc2889.INIT=64'h3F5FCFAF3050C0A0;
  LUT6 desc2890(.I0(r0[10:10]),.I1(r0[11:11]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m110),.O(m169));
defparam desc2890.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2891(.I0(r0[8:8]),.I1(r0[9:9]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m112),.O(m114));
defparam desc2891.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2892(.I0(r0[7:7]),.I1(r0[6:6]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m113),.O(m174));
defparam desc2892.INIT=64'h3F5FCFAF3050C0A0;
  LUT6 desc2893(.I0(r0[7:7]),.I1(r0[6:6]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m55_lut6_2_O5),.O(m136));
defparam desc2893.INIT=64'hF3F5FCFA03050C0A;
  LUT6 v_r1_2_3_23_RNI0E9E7(.I0(b_2[8:8]),.I1(r0_2[8:8]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(v_r1_2_3_23),.I5(m132),.O(v_r1_2_3_0_axb_8));
defparam v_r1_2_3_23_RNI0E9E7.INIT=64'h6999966666969969;
  LUT3 v_r1_2_3_0_cry_8_RNO_cZ(.I0(b_2[8:8]),.I1(r0_2[8:8]),.I2(v_r1_2_3_23),.O(v_r1_2_3_0_cry_8_RNO));
defparam v_r1_2_3_0_cry_8_RNO_cZ.INIT=8'h96;
  LUT6 v_r1_2_3_63_2_0_RNI05SSU(.I0(b_2[20:20]),.I1(r0_2[20:20]),.I2(r0_2[19:19]),.I3(N_48_i),.I4(v_r1_2_3_63_2_0),.I5(v_r1_2_3_25),.O(v_r1_2_3_0_axb_20));
defparam v_r1_2_3_63_2_0_RNI05SSU.INIT=64'h6996699669969966;
  LUT5 v_r1_2_3_0_cry_20_RNO_cZ(.I0(b_2[20:20]),.I1(r0_2[20:20]),.I2(r0_2[19:19]),.I3(v_r1_2_3_63_2_0),.I4(v_r1_2_3_25),.O(v_r1_2_3_0_cry_20_RNO));
defparam v_r1_2_3_0_cry_20_RNO_cZ.INIT=32'h96969666;
  LUT6 v_r1_2_3_51_RNIV701C(.I0(b_2[16:16]),.I1(r0_2[16:16]),.I2(c[4:4]),.I3(m145),.I4(m125),.I5(v_r1_2_3_51),.O(v_r1_2_3_0_axb_16));
defparam v_r1_2_3_51_RNIV701C.INIT=64'h9666996969996696;
  LUT6 v_r1_2_3_9_RNI0RGH5(.I0(b_2[4:4]),.I1(r0_2[4:4]),.I2(c[4:4]),.I3(v_r1_2_3_9),.I4(un14_s_state_cry[50:50]),.I5(m143),.O(v_r1_2_3_0_axb_4));
defparam v_r1_2_3_9_RNI0RGH5.INIT=64'h6996996666999669;
  LUT3 v_r1_2_3_0_cry_4_RNO_cZ(.I0(b_2[4:4]),.I1(r0_2[4:4]),.I2(v_r1_2_3_9),.O(v_r1_2_3_0_cry_4_RNO));
defparam v_r1_2_3_0_cry_4_RNO_cZ.INIT=8'h96;
  LUT6 desc2894(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[0:0]),.I3(c[4:4]),.I4(un14_s_state_cry[50:50]),.I5(m193),.O(v_r1_2_3_0_axb_1));
defparam desc2894.INIT=64'h936C6C6C93936C93;
  LUT6 v_r1_2_3_0_cry_18_RNO_cZ(.I0(b_2[18:18]),.I1(r0_2[18:18]),.I2(b_2[16:16]),.I3(r0_2[17:17]),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_0_cry_18_RNO));
defparam v_r1_2_3_0_cry_18_RNO_cZ.INIT=64'h9966966699666666;
  LUT6_L v_r1_2_3_51_cZ(.I0(r0_2[14:14]),.I1(b_2[14:14]),.I2(r0_2[13:13]),.I3(r0_2[15:15]),.I4(v_r1_2_3_35_0_RNIKOE74),.I5(v_r1_2_3_49_0_tz),.LO(v_r1_2_3_51));
defparam v_r1_2_3_51_cZ.INIT=64'hEC00CC00A0000000;
  LUT6 desc2895(.I0(b_2[10:10]),.I1(r0_2[10:10]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(v_r1_2_3_21_2_RNIQ1CU_O5),.I5(m71_lut6_2_O6),.O(v_r1_2_3_0_axb_10));
defparam desc2895.INIT=64'h6999966666969969;
  LUT6 desc2896(.I0(b_2[12:12]),.I1(r0_2[12:12]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(v_r1_2_3_35_0_RNI40J52_O5),.I5(m129),.O(v_r1_2_3_0_axb_12));
defparam desc2896.INIT=64'h6999966666969969;
  LUT6 v_r1_2_3_16_RNI4ECC5(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(c[4:4]),.I3(v_r1_2_3_16),.I4(un14_s_state_cry[50:50]),.I5(m73_lut6_2_O6),.O(v_r1_2_3_0_axb_6));
defparam v_r1_2_3_16_RNI4ECC5.INIT=64'h6996996666999669;
  LUT6 v_r1_2_3_44_lut6_2_RNIL0LI9(.I0(r0_2[14:14]),.I1(b_2[14:14]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(v_r1_2_3_44_lut6_2_O6),.I5(m67),.O(v_r1_2_3_0_axb_14));
defparam v_r1_2_3_44_lut6_2_RNIL0LI9.INIT=64'h6999966666969969;
  LUT6 v_r1_2_3_2_RNI7PDE5(.I0(b_2[2:2]),.I1(r0_2[2:2]),.I2(c[4:4]),.I3(v_r1_2_3_2),.I4(un14_s_state_cry[50:50]),.I5(m73_lut6_2_O5),.O(v_r1_2_3_0_axb_2));
defparam v_r1_2_3_2_RNI7PDE5.INIT=64'h6996996666999669;
  LUT3 v_r1_2_3_0_cry_1_RNO_cZ(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[0:0]),.O(v_r1_2_3_0_cry_1_RNO));
defparam v_r1_2_3_0_cry_1_RNO_cZ.INIT=8'h6C;
  LUT5 v_r1_2_3_0_cry_2_RNO_cZ(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[0:0]),.I3(b_2[2:2]),.I4(r0_2[2:2]),.O(v_r1_2_3_0_cry_2_RNO));
defparam v_r1_2_3_0_cry_2_RNO_cZ.INIT=32'h807F7F80;
  LUT6 v_r1_2_3_0_cry_3_RNO_cZ(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[3:3]),.I3(r0_2[0:0]),.I4(b_2[2:2]),.I5(r0_2[2:2]),.O(v_r1_2_3_0_cry_3_RNO));
defparam v_r1_2_3_0_cry_3_RNO_cZ.INIT=64'h0F0F78F078F0F0F0;
  LUT5 desc2897(.I0(c[1:1]),.I1(c[2:2]),.I2(m35),.I3(m32),.I4(m25),.O(N_50_0));
defparam desc2897.INIT=32'hF7B3C480;
  LUT5 desc2898(.I0(c[1:1]),.I1(c[2:2]),.I2(m24_lut6_2_O6),.I3(m32),.I4(m84),.O(m90));
defparam desc2898.INIT=32'hFB73C840;
  LUT5 desc2899(.I0(c[1:1]),.I1(c[2:2]),.I2(m24_lut6_2_O6),.I3(m32),.I4(N_95_0),.O(N_96_0));
defparam desc2899.INIT=32'hFEDC3210;
  LUT6 desc2900(.I0(c[2:2]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m139),.I5(m207),.O(N_3022_i));
defparam desc2900.INIT=64'hFF1FEF0FF010E000;
  LUT6 v_r1_2_3_0_cry_7_RNO_cZ(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(r0_2[7:7]),.I4(v_r1_2_3_4),.I5(v_r1_2_3_14_0),.O(v_r1_2_3_0_cry_7_RNO));
defparam v_r1_2_3_0_cry_7_RNO_cZ.INIT=64'h17E817E817E87788;
  LUT5 v_r1_2_3_0_cry_6_RNO_cZ(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(v_r1_2_3_4),.I4(v_r1_2_3_14_0),.O(v_r1_2_3_0_cry_6_RNO));
defparam v_r1_2_3_0_cry_6_RNO_cZ.INIT=32'h96969666;
  LUT4 v_r1_2_3_0_cry_45_RNO_cZ(.I0(r0_2[45:45]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m166),.O(v_r1_2_3_0_cry_45_RNO));
defparam v_r1_2_3_0_cry_45_RNO_cZ.INIT=16'h569A;
  LUT4 v_r1_2_3_0_cry_46_RNO_cZ(.I0(r0_2[45:45]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m166),.O(v_r1_2_3_0_cry_46_RNO));
defparam v_r1_2_3_0_cry_46_RNO_cZ.INIT=16'hA820;
  LUT6 v_r1_2_3_0_cry_31_RNO_cZ(.I0(r0_2[31:31]),.I1(c[3:3]),.I2(c[4:4]),.I3(m100),.I4(m108),.I5(m182),.O(v_r1_2_3_0_cry_31_RNO));
defparam v_r1_2_3_0_cry_31_RNO_cZ.INIT=64'h595A5556A9AAA5A6;
  LUT4 v_r1_2_3_0_cry_30_RNO_cZ(.I0(r0_2[29:29]),.I1(c[4:4]),.I2(m186),.I3(m166),.O(v_r1_2_3_0_cry_30_RNO));
defparam v_r1_2_3_0_cry_30_RNO_cZ.INIT=16'h2A08;
  LUT4 v_r1_2_3_0_cry_41_RNO_cZ(.I0(r0_2[41:41]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m171),.O(v_r1_2_3_0_cry_41_RNO));
defparam v_r1_2_3_0_cry_41_RNO_cZ.INIT=16'h569A;
  LUT4 v_r1_2_3_0_cry_34_RNO_cZ(.I0(r0_2[33:33]),.I1(c[4:4]),.I2(m159),.I3(m180),.O(v_r1_2_3_0_cry_34_RNO));
defparam v_r1_2_3_0_cry_34_RNO_cZ.INIT=16'hA820;
  LUT6 v_r1_2_3_0_cry_43_RNO_cZ(.I0(r0_2[43:43]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m203),.I5(m200),.O(v_r1_2_3_0_cry_43_RNO));
defparam v_r1_2_3_0_cry_43_RNO_cZ.INIT=64'h555A959A656AA5AA;
  LUT6 v_r1_2_3_0_cry_47_RNO_cZ(.I0(r0_2[47:47]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m100),.I5(m108),.O(v_r1_2_3_0_cry_47_RNO));
defparam v_r1_2_3_0_cry_47_RNO_cZ.INIT=64'h959AA5AA555A656A;
  LUT4 v_r1_2_3_0_cry_42_RNO_cZ(.I0(r0_2[41:41]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m171),.O(v_r1_2_3_0_cry_42_RNO));
defparam v_r1_2_3_0_cry_42_RNO_cZ.INIT=16'hA820;
  LUT6 v_r1_2_3_0_cry_44_RNO_cZ(.I0(r0_2[43:43]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m203),.I5(m200),.O(v_r1_2_3_0_cry_44_RNO));
defparam v_r1_2_3_0_cry_44_RNO_cZ.INIT=64'hAAA02A208A800A00;
  LUT6 v_r1_2_3_0_cry_48_RNO_cZ(.I0(r0_2[47:47]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m100),.I5(m108),.O(v_r1_2_3_0_cry_48_RNO));
defparam v_r1_2_3_0_cry_48_RNO_cZ.INIT=64'h2A200A00AAA08A80;
  LUT6 v_r1_2_3_0_cry_32_RNO_cZ(.I0(r0_2[31:31]),.I1(c[3:3]),.I2(c[4:4]),.I3(m100),.I4(m108),.I5(m182),.O(v_r1_2_3_0_cry_32_RNO));
defparam v_r1_2_3_0_cry_32_RNO_cZ.INIT=64'hA2A0AAA802000A08;
  LUT4 v_r1_2_3_0_cry_26_RNO_cZ(.I0(r0_2[25:25]),.I1(c[4:4]),.I2(m189),.I3(m171),.O(v_r1_2_3_0_cry_26_RNO));
defparam v_r1_2_3_0_cry_26_RNO_cZ.INIT=16'h2A08;
  LUT5 v_r1_2_3_0_axb_27_cZ(.I0(b_2[26:26]),.I1(r0_2[26:26]),.I2(r0_2[27:27]),.I3(m211),.I4(N_2891_i),.O(v_r1_2_3_0_axb_27));
defparam v_r1_2_3_0_axb_27_cZ.INIT=32'h1EE17887;
  LUT6_L v_r1_2_3_175_cZ(.I0(b_2[50:50]),.I1(r0_2[50:50]),.I2(c[3:3]),.I3(c[4:4]),.I4(un14_s_state_cry[50:50]),.I5(m47),.LO(v_r1_2_3_175));
defparam v_r1_2_3_175_cZ.INIT=64'hEEEEE8888EEE8888;
  LUT4 v_r1_2_3_0_cry_33_RNO_cZ(.I0(r0_2[33:33]),.I1(c[4:4]),.I2(m159),.I3(m180),.O(v_r1_2_3_0_cry_33_RNO));
defparam v_r1_2_3_0_cry_33_RNO_cZ.INIT=16'h569A;
  LUT6 v_r1_2_3_0_cry_10_RNO_cZ(.I0(b_2[8:8]),.I1(r0_2[9:9]),.I2(v_r1_2_3_31_0),.I3(v_r1_2_3_27_0),.I4(v_r1_2_3_28_0_tz),.I5(v_r1_2_3_21_2),.O(v_r1_2_3_0_cry_10_RNO));
defparam v_r1_2_3_0_cry_10_RNO_cZ.INIT=64'h3C783CF07878F0F0;
  LUT4 v_r1_2_3_0_cry_29_RNO_cZ(.I0(r0_2[29:29]),.I1(c[4:4]),.I2(m186),.I3(m166),.O(v_r1_2_3_0_cry_29_RNO));
defparam v_r1_2_3_0_cry_29_RNO_cZ.INIT=16'h95A6;
  LUT6 v_r1_2_3_0_cry_28_RNO_cZ(.I0(r0_2[27:27]),.I1(c[3:3]),.I2(c[4:4]),.I3(m203),.I4(m200),.I5(m210),.O(v_r1_2_3_0_cry_28_RNO));
defparam v_r1_2_3_0_cry_28_RNO_cZ.INIT=64'h0A020800AAA2A8A0;
  LUT6 v_r1_2_3_0_cry_35_RNO_cZ(.I0(r0_2[35:35]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m200),.I5(m207),.O(v_r1_2_3_0_cry_35_RNO));
defparam v_r1_2_3_0_cry_35_RNO_cZ.INIT=64'h5556595AA5A6A9AA;
  LUT6 v_r1_2_3_0_cry_36_RNO_cZ(.I0(r0_2[35:35]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m200),.I5(m207),.O(v_r1_2_3_0_cry_36_RNO));
defparam v_r1_2_3_0_cry_36_RNO_cZ.INIT=64'hAAA8A2A00A080200;
  LUT6 v_r1_2_3_0_cry_12_RNO_cZ(.I0(b_2[12:12]),.I1(r0_2[12:12]),.I2(r0_2[11:11]),.I3(v_r1_2_3_34_0),.I4(v_r1_2_3_35_0),.I5(v_r1_2_3_21_2_RNIMLGQ),.O(v_r1_2_3_0_cry_12_RNO));
defparam v_r1_2_3_0_cry_12_RNO_cZ.INIT=64'h9696966696966666;
  LUT6 v_r1_2_3_0_cry_14_RNO_cZ(.I0(r0_2[14:14]),.I1(b_2[14:14]),.I2(r0_2[13:13]),.I3(v_r1_2_3_41_0),.I4(b_2_RNIMF314[10:10]),.I5(v_r1_2_3_42_0),.O(v_r1_2_3_0_cry_14_RNO));
defparam v_r1_2_3_0_cry_14_RNO_cZ.INIT=64'h9696969696666666;
  LUT6 v_r1_2_3_0_cry_16_RNO_cZ(.I0(b_2[14:14]),.I1(r0_2[15:15]),.I2(v_r1_2_3_48_0),.I3(v_r1_2_3_52_0),.I4(v_r1_2_3_35_0_RNIKOE74),.I5(v_r1_2_3_49_0_tz),.O(v_r1_2_3_0_cry_16_RNO));
defparam v_r1_2_3_0_cry_16_RNO_cZ.INIT=64'h37C877883FC0FF00;
  LUT6 v_r1_2_3_59_0_lut6_2_RNIF122G1(.I0(b_2[16:16]),.I1(r0_2[17:17]),.I2(v_r1_2_3_59_0),.I3(N_2895_i),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_0_axb_18));
defparam v_r1_2_3_59_0_lut6_2_RNIF122G1.INIT=64'hC33C8778C33C0FF0;
  LUT6 v_r1_2_3_0_cry_17_RNO_cZ(.I0(b_2[16:16]),.I1(r0_2[16:16]),.I2(r0_2[17:17]),.I3(r0_2[15:15]),.I4(v_r1_2_3_49),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_0_cry_17_RNO));
defparam v_r1_2_3_0_cry_17_RNO_cZ.INIT=64'h1E5A5A5A3CF0F0F0;
  LUT6 v_r1_2_3_0_cry_22_RNO_cZ(.I0(b_2[20:20]),.I1(r0_2[21:21]),.I2(v_r1_2_3_73_0),.I3(v_r1_2_3_28),.I4(v_r1_2_3_65_c),.I5(v_r1_2_3_65_0_0),.O(v_r1_2_3_0_cry_22_RNO));
defparam v_r1_2_3_0_cry_22_RNO_cZ.INIT=64'h3C783C783C783CF0;
  LUT5 v_r1_2_3_0_cry_21_RNO_cZ(.I0(b_2[20:20]),.I1(r0_2[21:21]),.I2(v_r1_2_3_28),.I3(v_r1_2_3_65_c),.I4(v_r1_2_3_65_0_0),.O(v_r1_2_3_0_cry_21_RNO));
defparam v_r1_2_3_0_cry_21_RNO_cZ.INIT=32'h3636363C;
  LUT5 v_r1_2_3_0_axb_25_cZ(.I0(b_2[24:24]),.I1(r0_2[25:25]),.I2(r0_2[24:24]),.I3(m190_lut6_2_O6),.I4(v_r1_2_3_73_0_lut6_2_RNIM5CP22),.O(v_r1_2_3_0_axb_25));
defparam v_r1_2_3_0_axb_25_cZ.INIT=32'h36C96C93;
  MUXCY_L v_r1_2_3_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(v_r1_2_3_scalar),.LO(v_r1_2_3_0_cry_0_cy));
  LUT2_L un1_r1_axb_24_cZ(.I0(r1[24:24]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_24));
defparam un1_r1_axb_24_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_23_cZ(.I0(r1[23:23]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_23));
defparam un1_r1_axb_23_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_22_cZ(.I0(r1[22:22]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_22));
defparam un1_r1_axb_22_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_21_cZ(.I0(r1[21:21]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_21));
defparam un1_r1_axb_21_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_20_cZ(.I0(r1[20:20]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_20));
defparam un1_r1_axb_20_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_19_cZ(.I0(r1[19:19]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_19));
defparam un1_r1_axb_19_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_18_cZ(.I0(r1[18:18]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_18));
defparam un1_r1_axb_18_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_17_cZ(.I0(r1[17:17]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_17));
defparam un1_r1_axb_17_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_16_cZ(.I0(r1[16:16]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_16));
defparam un1_r1_axb_16_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_15_cZ(.I0(r1[15:15]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_15));
defparam un1_r1_axb_15_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_14_cZ(.I0(r1[14:14]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_14));
defparam un1_r1_axb_14_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_13_cZ(.I0(r1[13:13]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_13));
defparam un1_r1_axb_13_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_12_cZ(.I0(r1[12:12]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_12));
defparam un1_r1_axb_12_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_11_cZ(.I0(r1[11:11]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_11));
defparam un1_r1_axb_11_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_10_cZ(.I0(r1[10:10]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_10));
defparam un1_r1_axb_10_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_9_cZ(.I0(r1[9:9]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_9));
defparam un1_r1_axb_9_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_8_cZ(.I0(r1[8:8]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_8));
defparam un1_r1_axb_8_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_7_cZ(.I0(r1[7:7]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_7));
defparam un1_r1_axb_7_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_6_cZ(.I0(r1[6:6]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_6));
defparam un1_r1_axb_6_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_5_cZ(.I0(r1[5:5]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_5));
defparam un1_r1_axb_5_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_4_cZ(.I0(r1[4:4]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_4));
defparam un1_r1_axb_4_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_3_cZ(.I0(r1[3:3]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_3));
defparam un1_r1_axb_3_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_2_cZ(.I0(r1[2:2]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_2));
defparam un1_r1_axb_2_cZ.INIT=4'h6;
  LUT2_L un1_r1_axb_1_cZ(.I0(r1[1:1]),.I1(un27_s_count_cry[50:50]),.LO(un1_r1_axb_1));
defparam un1_r1_axb_1_cZ.INIT=4'h6;
  LUT2 un1_r1_axb_0_cZ(.I0(r1[0:0]),.I1(un27_s_count_cry[50:50]),.O(un1_r1_axb_0));
defparam un1_r1_axb_0_cZ.INIT=4'h6;
  LUT2_L v_r1_2_3_0_cZ(.I0(b_2_fast),.I1(r0_2_fast[0:0]),.LO(v_r1_2_3_0));
defparam v_r1_2_3_0_cZ.INIT=4'h8;
  LUT1_L desc2901(.I0(c[0:0]),.LO(c_i));
defparam desc2901.INIT=2'h1;
  LUT4 s_ine_o_e_RNO_8(.I0(un33_s_count_a_5[8:8]),.I1(un33_s_count_a_5[9:9]),.I2(un33_s_count_a_5[10:10]),.I3(un33_s_count_a_5[11:11]),.O(un33_s_count_NE_1_3));
defparam s_ine_o_e_RNO_8.INIT=16'h7FFF;
  LUT4_L s_ine_o_e_RNO_7(.I0(un33_s_count_a_5[2:2]),.I1(un33_s_count_a_5[3:3]),.I2(un33_s_count_a_5[4:4]),.I3(un33_s_count_a_5[5:5]),.LO(un33_s_count_NE_0_3));
defparam s_ine_o_e_RNO_7.INIT=16'h7FFF;
  LUT2 un33_s_count_a_5_0_o5_16_cZ(.I0(r1[15:15]),.I1(r1_2[16:16]),.O(un33_s_count_a_5_0_o5_16));
defparam un33_s_count_a_5_0_o5_16_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_21_cZ(.I0(r1[20:20]),.I1(r1_2[21:21]),.O(un33_s_count_a_5_0_o5_21));
defparam un33_s_count_a_5_0_o5_21_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_17_cZ(.I0(r1[16:16]),.I1(r1_2[17:17]),.O(un33_s_count_a_5_0_o5_17));
defparam un33_s_count_a_5_0_o5_17_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_4_cZ(.I0(r1[3:3]),.I1(r1_2[4:4]),.O(un33_s_count_a_5_0_o5_4));
defparam un33_s_count_a_5_0_o5_4_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_20_cZ(.I0(r1[19:19]),.I1(r1_2[20:20]),.O(un33_s_count_a_5_0_o5_20));
defparam un33_s_count_a_5_0_o5_20_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_18_cZ(.I0(r1[17:17]),.I1(r1_2[18:18]),.O(un33_s_count_a_5_0_o5_18));
defparam un33_s_count_a_5_0_o5_18_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_6_cZ(.I0(r1[5:5]),.I1(r1_2[6:6]),.O(un33_s_count_a_5_0_o5_6));
defparam un33_s_count_a_5_0_o5_6_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_3_cZ(.I0(r1[2:2]),.I1(r1_2[3:3]),.O(un33_s_count_a_5_0_o5_3));
defparam un33_s_count_a_5_0_o5_3_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_14_cZ(.I0(r1[13:13]),.I1(r1_2[14:14]),.O(un33_s_count_a_5_0_o5_14));
defparam un33_s_count_a_5_0_o5_14_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_23_cZ(.I0(r1[22:22]),.I1(r1_2[23:23]),.O(un33_s_count_a_5_0_o5_23));
defparam un33_s_count_a_5_0_o5_23_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_9_cZ(.I0(r1[8:8]),.I1(r1_2[9:9]),.O(un33_s_count_a_5_0_o5_9));
defparam un33_s_count_a_5_0_o5_9_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_10_cZ(.I0(r1[9:9]),.I1(r1_2[10:10]),.O(un33_s_count_a_5_0_o5_10));
defparam un33_s_count_a_5_0_o5_10_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_15_cZ(.I0(r1[14:14]),.I1(r1_2[15:15]),.O(un33_s_count_a_5_0_o5_15));
defparam un33_s_count_a_5_0_o5_15_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_19_cZ(.I0(r1[18:18]),.I1(r1_2[19:19]),.O(un33_s_count_a_5_0_o5_19));
defparam un33_s_count_a_5_0_o5_19_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_5_cZ(.I0(r1[4:4]),.I1(r1_2[5:5]),.O(un33_s_count_a_5_0_o5_5));
defparam un33_s_count_a_5_0_o5_5_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_8_cZ(.I0(r1[7:7]),.I1(r1_2[8:8]),.O(un33_s_count_a_5_0_o5_8));
defparam un33_s_count_a_5_0_o5_8_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_12_cZ(.I0(r1[11:11]),.I1(r1_2[12:12]),.O(un33_s_count_a_5_0_o5_12));
defparam un33_s_count_a_5_0_o5_12_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_24_cZ(.I0(r1[23:23]),.I1(r1_2[24:24]),.O(un33_s_count_a_5_0_o5_24));
defparam un33_s_count_a_5_0_o5_24_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_22_cZ(.I0(r1[21:21]),.I1(r1_2[22:22]),.O(un33_s_count_a_5_0_o5_22));
defparam un33_s_count_a_5_0_o5_22_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_13_cZ(.I0(r1[12:12]),.I1(r1_2[13:13]),.O(un33_s_count_a_5_0_o5_13));
defparam un33_s_count_a_5_0_o5_13_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_7_cZ(.I0(r1[6:6]),.I1(r1_2[7:7]),.O(un33_s_count_a_5_0_o5_7));
defparam un33_s_count_a_5_0_o5_7_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_o5_11_cZ(.I0(r1[10:10]),.I1(r1_2[11:11]),.O(un33_s_count_a_5_0_o5_11));
defparam un33_s_count_a_5_0_o5_11_cZ.INIT=4'hD;
  LUT3 v_r1_3_axb_25_cZ(.I0(b[25:25]),.I1(r0[25:25]),.I2(un14_s_state_cry[50:50]),.O(v_r1_3_axb_25));
defparam v_r1_3_axb_25_cZ.INIT=8'h96;
  LUT4 un33_s_count_a_5_0_axb_51_cZ(.I0(r1_2[51:51]),.I1(r1_2[50:50]),.I2(s_rad_i[51:51]),.I3(s_rad_i[50:50]),.O(un33_s_count_a_5_0_axb_51));
defparam un33_s_count_a_5_0_axb_51_cZ.INIT=16'hA569;
  LUT3 v_r1_2_3_2_cZ(.I0(b_2_fast),.I1(r0_2_fast[0:0]),.I2(r0_2_fast[1:1]),.O(v_r1_2_3_2));
defparam v_r1_2_3_2_cZ.INIT=8'h80;
  LUT4 desc2902(.I0(r0[8:8]),.I1(r0[9:9]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m113));
defparam desc2902.INIT=16'h53AC;
  LUT4 desc2903(.I0(r0[10:10]),.I1(r0[11:11]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m112));
defparam desc2903.INIT=16'h53AC;
  LUT4 desc2904(.I0(r0[12:12]),.I1(r0[13:13]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m110));
defparam desc2904.INIT=16'h53AC;
  LUT4 desc2905(.I0(r0[15:15]),.I1(r0[14:14]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m109));
defparam desc2905.INIT=16'h35CA;
  LUT4 desc2906(.I0(r0[16:16]),.I1(r0[17:17]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m106));
defparam desc2906.INIT=16'hAC53;
  LUT4 desc2907(.I0(r0[19:19]),.I1(r0[18:18]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m105));
defparam desc2907.INIT=16'h35CA;
  LUT4 desc2908(.I0(r0[7:7]),.I1(r0[8:8]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m42));
defparam desc2908.INIT=16'h53AC;
  LUT4 desc2909(.I0(r0[12:12]),.I1(r0[11:11]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m35));
defparam desc2909.INIT=16'h35CA;
  LUT4 desc2910(.I0(r0[13:13]),.I1(r0[14:14]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m32));
defparam desc2910.INIT=16'h53AC;
  LUT6 s_ine_o_e_RNO_3(.I0(un33_s_count_29),.I1(un33_s_count_30),.I2(un33_s_count_31),.I3(un33_s_count_32),.I4(un33_s_count_33),.I5(un33_s_count_34),.O(un33_s_count_NE_5));
defparam s_ine_o_e_RNO_3.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L s_ine_o_e_RNO_6(.I0(un33_s_count_a_5[18:18]),.I1(un33_s_count_a_5[19:19]),.I2(un33_s_count_a_5[20:20]),.I3(un33_s_count_a_5[21:21]),.I4(un33_s_count_a_5[22:22]),.I5(un33_s_count_a_5[23:23]),.LO(un33_s_count_NE_3));
defparam s_ine_o_e_RNO_6.INIT=64'h7FFFFFFFFFFFFFFF;
  LUT6_L s_ine_o_e_RNO_9(.I0(un33_s_count_a_5[12:12]),.I1(un33_s_count_a_5[13:13]),.I2(un33_s_count_a_5[14:14]),.I3(un33_s_count_a_5[15:15]),.I4(un33_s_count_a_5[16:16]),.I5(un33_s_count_a_5[17:17]),.LO(un33_s_count_NE_2));
defparam s_ine_o_e_RNO_9.INIT=64'h7FFFFFFFFFFFFFFF;
  LUT6 un31_s_count_0_I_138(.I0(r1_2[50:50]),.I1(r1_2[48:48]),.I2(r1_2[49:49]),.I3(s_rad_i[50:50]),.I4(s_rad_i[48:48]),.I5(s_rad_i[49:49]),.O(un31_s_count_0_N_4));
defparam un31_s_count_0_I_138.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_90(.I0(r1_2[30:30]),.I1(r1_2[31:31]),.I2(r1_2[32:32]),.I3(s_rad_i[30:30]),.I4(s_rad_i[31:31]),.I5(s_rad_i[32:32]),.O(un31_s_count_0_N_46));
defparam un31_s_count_0_I_90.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_114(.I0(r1_2[39:39]),.I1(r1_2[40:40]),.I2(r1_2[41:41]),.I3(s_rad_i[39:39]),.I4(s_rad_i[40:40]),.I5(s_rad_i[41:41]),.O(un31_s_count_0_N_25));
defparam un31_s_count_0_I_114.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_82(.I0(r1_2[27:27]),.I1(r1_2[28:28]),.I2(r1_2[29:29]),.I3(s_rad_i[27:27]),.I4(s_rad_i[28:28]),.I5(s_rad_i[29:29]),.O(un31_s_count_0_N_53));
defparam un31_s_count_0_I_82.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_106(.I0(r1_2[36:36]),.I1(r1_2[37:37]),.I2(r1_2[38:38]),.I3(s_rad_i[36:36]),.I4(s_rad_i[37:37]),.I5(s_rad_i[38:38]),.O(un31_s_count_0_N_32));
defparam un31_s_count_0_I_106.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_122(.I0(r1_2[42:42]),.I1(r1_2[43:43]),.I2(r1_2[44:44]),.I3(s_rad_i[42:42]),.I4(s_rad_i[43:43]),.I5(s_rad_i[44:44]),.O(un31_s_count_0_N_18));
defparam un31_s_count_0_I_122.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_130(.I0(r1_2[45:45]),.I1(r1_2[46:46]),.I2(r1_2[47:47]),.I3(s_rad_i[45:45]),.I4(s_rad_i[46:46]),.I5(s_rad_i[47:47]),.O(un31_s_count_0_N_11));
defparam un31_s_count_0_I_130.INIT=64'h8040201008040201;
  LUT6 un31_s_count_0_I_98(.I0(r1_2[33:33]),.I1(r1_2[34:34]),.I2(r1_2[35:35]),.I3(s_rad_i[33:33]),.I4(s_rad_i[34:34]),.I5(s_rad_i[35:35]),.O(un31_s_count_0_N_39));
defparam un31_s_count_0_I_98.INIT=64'h8040201008040201;
  LUT3 v_r1_2_3_0_o5_26_cZ(.I0(b_2[26:26]),.I1(r0_2[26:26]),.I2(N_2891_i),.O(v_r1_2_3_0_o5_26));
defparam v_r1_2_3_0_o5_26_cZ.INIT=8'hE8;
  LUT3 v_r1_2_3_0_o5_24_cZ(.I0(b_2[24:24]),.I1(r0_2[24:24]),.I2(v_r1_2_3_73_0_lut6_2_RNIM5CP22),.O(v_r1_2_3_0_o5_24));
defparam v_r1_2_3_0_o5_24_cZ.INIT=8'hE8;
  LUT6 desc2911(.I0(r0[3:3]),.I1(r0[2:2]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m55_lut6_2_O5),.O(m178));
defparam desc2911.INIT=64'h3F5FCFAF3050C0A0;
  LUT6 desc2912(.I0(r0[15:15]),.I1(r0[14:14]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m106),.O(m164));
defparam desc2912.INIT=64'h3050C0A03F5FCFAF;
  LUT6 desc2913(.I0(r0[23:23]),.I1(r0[22:22]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m9_lut6_2_O5),.O(m156));
defparam desc2913.INIT=64'h3F5FCFAF3050C0A0;
  LUT6 desc2914(.I0(r0[3:3]),.I1(r0[2:2]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m138_lut6_2_O6),.O(m139));
defparam desc2914.INIT=64'hF3F5FCFA03050C0A;
  LUT6 desc2915(.I0(r0[1:1]),.I1(r0[2:2]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m55_lut6_2_O6),.O(m123));
defparam desc2915.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2916(.I0(r0[5:5]),.I1(r0[6:6]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m42),.O(m119));
defparam desc2916.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2917(.I0(r0[23:23]),.I1(r0[22:22]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m17_lut6_2_O5),.O(m104));
defparam desc2917.INIT=64'hF3F5FCFA03050C0A;
  LUT6 desc2918(.I0(r0[9:9]),.I1(r0[10:10]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m35),.O(N_95_0));
defparam desc2918.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2919(.I0(r0[17:17]),.I1(r0[18:18]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(N_18_1),.O(m84));
defparam desc2919.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2920(.I0(r0[21:21]),.I1(r0[22:22]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(N_10_1),.O(N_84_0));
defparam desc2920.INIT=64'h5F3FAFCF5030A0C0;
  LUT6 desc2921(.I0(r0[1:1]),.I1(r0[2:2]),.I2(r0[0:0]),.I3(c[1:1]),.I4(c[0:0]),.I5(un14_s_state_cry[50:50]),.O(m65));
defparam desc2921.INIT=64'h00AAF0CCFF550F33;
  LUT6 desc2922(.I0(r0[5:5]),.I1(r0[6:6]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m55_lut6_2_O6),.O(m56));
defparam desc2922.INIT=64'hF5F3FAFC05030A0C;
  LUT6 desc2923(.I0(r0[9:9]),.I1(r0[10:10]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m42),.O(m43));
defparam desc2923.INIT=64'hF5F3FAFC05030A0C;
  LUT6 desc2924(.I0(r0[17:17]),.I1(r0[18:18]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(m24_lut6_2_O6),.O(m25));
defparam desc2924.INIT=64'hF5F3FAFC05030A0C;
  LUT6 desc2925(.I0(r0[21:21]),.I1(r0[22:22]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.I5(N_18_1),.O(N_19_1));
defparam desc2925.INIT=64'hF5F3FAFC05030A0C;
  LUT6_L s_ine_o_e_RNO_4(.I0(un33_s_count_a_5[6:6]),.I1(un33_s_count_a_5[7:7]),.I2(un33_s_count_NE_1_3),.I3(un33_s_count_37),.I4(un33_s_count_38),.I5(un33_s_count_39),.LO(un33_s_count_NE_6_3));
defparam s_ine_o_e_RNO_4.INIT=64'hFFFFFFFFFFFFFFF7;
  LUT6 s_ine_o_e_RNO_2(.I0(r1_2[0:0]),.I1(un33_s_count_1),.I2(un33_s_count_a_5[26:26]),.I3(un33_s_count_27),.I4(un33_s_count_28),.I5(un33_s_count_NE_0_3),.O(un33_s_count_NE_4_3));
defparam s_ine_o_e_RNO_2.INIT=64'hFFFFFFFFFFFFFFDF;
  LUT5 v_r1_2_3_7_cZ(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[0:0]),.I3(b_2[2:2]),.I4(r0_2[2:2]),.O(v_r1_2_3_7));
defparam v_r1_2_3_7_cZ.INIT=32'hFF808000;
  LUT6 desc2926(.I0(c[1:1]),.I1(c[2:2]),.I2(m105),.I3(m109),.I4(m106),.I5(m110),.O(m203));
defparam desc2926.INIT=64'hDC98FEBA54107632;
  LUT5 desc2927(.I0(c[1:1]),.I1(c[2:2]),.I2(un14_s_state_cry[50:50]),.I3(m9_lut6_2_O5),.I4(m104),.O(m200));
defparam desc2927.INIT=32'hFEDC3210;
  LUT6 desc2928(.I0(c[1:1]),.I1(c[2:2]),.I2(m109),.I3(m112),.I4(m113),.I5(m110),.O(m115));
defparam desc2928.INIT=64'hFEBA7632DC985410;
  LUT5 desc2929(.I0(c[1:1]),.I1(c[2:2]),.I2(m105),.I3(m106),.I4(m104),.O(m108));
defparam desc2929.INIT=32'h8C04BF37;
  LUT6 desc2930(.I0(r0[24:24]),.I1(r0[25:25]),.I2(c[1:1]),.I3(c[2:2]),.I4(c[0:0]),.I5(un14_s_state_cry[50:50]),.O(m100));
defparam desc2930.INIT=64'h5FFF3FFFA000C000;
  LUT5 desc2931(.I0(c[1:1]),.I1(c[2:2]),.I2(m24_lut6_2_O5),.I3(N_10_1),.I4(N_19_1),.O(m47));
defparam desc2931.INIT=32'hFEDC3210;
  LUT6 s_ine_o_e_RNO_0(.I0(un33_s_count_45),.I1(un33_s_count_46),.I2(un33_s_count_47),.I3(un33_s_count_48),.I4(un33_s_count_49),.I5(un33_s_count_NE_3),.O(un33_s_count_NE_8));
defparam s_ine_o_e_RNO_0.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6_L s_ine_o_e_RNO_5(.I0(un33_s_count_40),.I1(un33_s_count_41),.I2(un33_s_count_42),.I3(un33_s_count_43),.I4(un33_s_count_44),.I5(un33_s_count_NE_2),.LO(un33_s_count_NE_7));
defparam s_ine_o_e_RNO_5.INIT=64'hFFFFFFFFFFFFFFFE;
  LUT6 v_r1_2_3_13(.I0(r0_2_fast[1:1]),.I1(r0_2[4:4]),.I2(r0_2[3:3]),.I3(b_2[2:2]),.I4(r0_2[2:2]),.I5(v_r1_2_3_0),.O(v_r1_2_3_4));
defparam v_r1_2_3_13.INIT=64'hC0808000C0000000;
  LUT6 v_r1_2_3_9_cZ(.I0(b_2[0:0]),.I1(r0_2[1:1]),.I2(r0_2[3:3]),.I3(r0_2[0:0]),.I4(b_2[2:2]),.I5(r0_2[2:2]),.O(v_r1_2_3_9));
defparam v_r1_2_3_9_cZ.INIT=64'hF0F0800080000000;
  LUT5 s_ine_o_e_RNO(.I0(un33_s_count_35),.I1(un33_s_count_36),.I2(un33_s_count_50),.I3(un33_s_count_51),.I4(un33_s_count_NE_6_3),.O(un33_s_count_NE_1_4));
defparam s_ine_o_e_RNO.INIT=32'hFFFFFFFE;
  LUT6 v_r1_2_3_14_0_cZ(.I0(b_2[4:4]),.I1(r0_2[4:4]),.I2(r0_2[3:3]),.I3(b_2[2:2]),.I4(r0_2[2:2]),.I5(v_r1_2_3_2),.O(v_r1_2_3_14_0));
defparam v_r1_2_3_14_0_cZ.INIT=64'hA8A8A888A8888888;
  LUT6 desc2932(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m114),.I4(m136),.I5(m139),.O(m210));
defparam desc2932.INIT=64'h08192A3B4C5D6E7F;
  LUT5 desc2933(.I0(c[2:2]),.I1(c[3:3]),.I2(m114),.I3(m136),.I4(m203),.O(m207));
defparam desc2933.INIT=32'hFB73C840;
  LUT5 desc2934(.I0(c[1:1]),.I1(c[2:2]),.I2(c[3:3]),.I3(un14_s_state_cry[50:50]),.I4(m138_lut6_2_O6),.O(m193));
defparam desc2934.INIT=32'h00FE01FF;
  LUT5 desc2935(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m138_lut6_2_O5),.I4(m178),.O(m191));
defparam desc2935.INIT=32'h2E0C3F1D;
  LUT6 desc2936(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m138_lut6_2_O5),.I4(m174),.I5(m178),.O(m189));
defparam desc2936.INIT=64'h4C085D196E2A7F3B;
  LUT6 desc2937(.I0(c[2:2]),.I1(c[3:3]),.I2(m138_lut6_2_O5),.I3(m174),.I4(m178),.I5(m169),.O(m186));
defparam desc2937.INIT=64'h80A2C4E691B3D5F7;
  LUT5 desc2938(.I0(c[2:2]),.I1(c[3:3]),.I2(m136),.I3(m139),.I4(m115),.O(m182));
defparam desc2938.INIT=32'hFB73C840;
  LUT6 desc2939(.I0(c[2:2]),.I1(c[3:3]),.I2(m174),.I3(m178),.I4(m164),.I5(m169),.O(m180));
defparam desc2939.INIT=64'hFB73EA62D951C840;
  LUT6 desc2940(.I0(c[2:2]),.I1(c[3:3]),.I2(m174),.I3(m157),.I4(m164),.I5(m169),.O(m176));
defparam desc2940.INIT=64'hF7E6D5C4B3A29180;
  LUT6 desc2941(.I0(c[2:2]),.I1(c[3:3]),.I2(m156),.I3(m157),.I4(m164),.I5(m169),.O(m171));
defparam desc2941.INIT=64'hFEDCBA9876543210;
  LUT6 desc2942(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m156),.I4(m157),.I5(m164),.O(m166));
defparam desc2942.INIT=64'hFEDCBA9876543210;
  LUT5 desc2943(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m156),.I4(m157),.O(m159));
defparam desc2943.INIT=32'hFCB87430;
  LUT6 desc2944(.I0(r0[0:0]),.I1(c[1:1]),.I2(c[2:2]),.I3(c[0:0]),.I4(c[3:3]),.I5(un14_s_state_cry[50:50]),.O(m145));
defparam desc2944.INIT=64'h00000002FFFFFFFD;
  LUT5 desc2945(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m127_lut6_2_O6),.I4(m123),.O(m143));
defparam desc2945.INIT=32'h2E0C3F1D;
  LUT6 desc2946(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m127_lut6_2_O6),.I4(m119),.I5(m123),.O(m132));
defparam desc2946.INIT=64'h4C085D196E2A7F3B;
  LUT6 desc2947(.I0(c[2:2]),.I1(c[3:3]),.I2(m127_lut6_2_O6),.I3(N_95_0),.I4(m119),.I5(m123),.O(m129));
defparam desc2947.INIT=64'h8091A2B3C4D5E6F7;
  LUT6 desc2948(.I0(c[2:2]),.I1(c[3:3]),.I2(N_90_0),.I3(N_95_0),.I4(m119),.I5(m123),.O(m125));
defparam desc2948.INIT=64'hFEDCBA9876543210;
  LUT6 desc2949(.I0(c[2:2]),.I1(c[3:3]),.I2(m84),.I3(N_90_0),.I4(N_95_0),.I5(m119),.O(m121));
defparam desc2949.INIT=64'hFEDCBA9876543210;
  LUT6 desc2950(.I0(c[2:2]),.I1(c[3:3]),.I2(m65),.I3(m36),.I4(m43),.I5(m56),.O(m67));
defparam desc2950.INIT=64'h8091A2B3C4D5E6F7;
  LUT6 desc2951(.I0(c[2:2]),.I1(c[3:3]),.I2(N_19_1),.I3(m36),.I4(m43),.I5(m25),.O(m45));
defparam desc2951.INIT=64'hFEBA7632DC985410;
  LUT5_L s_ine_o_e_RNO_1(.I0(un33_s_count_a_5[24:24]),.I1(un33_s_count_a_5[25:25]),.I2(un33_s_count_NE_4_3),.I3(un33_s_count_NE_5),.I4(un33_s_count_NE_7),.LO(un33_s_count_NE_2_4));
defparam s_ine_o_e_RNO_1.INIT=32'hFFFFFFF7;
  LUT6 v_r1_2_3_14_cZ(.I0(b_2[4:4]),.I1(r0_2[4:4]),.I2(r0_2[3:3]),.I3(b_2[2:2]),.I4(r0_2[2:2]),.I5(v_r1_2_3_2),.O(v_r1_2_3_14));
defparam v_r1_2_3_14_cZ.INIT=64'hE8E8E888E8888888;
  LUT5 desc2952(.I0(c[3:3]),.I1(c[4:4]),.I2(m203),.I3(m200),.I4(m210),.O(m211));
defparam desc2952.INIT=32'hCEDF0213;
  LUT5 desc2953(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m200),.I4(m207),.O(m208));
defparam desc2953.INIT=32'hFEDC3210;
  LUT5 desc2954(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m203),.I4(m200),.O(m205));
defparam desc2954.INIT=32'hFC74B830;
  LUT5 desc2955(.I0(c[3:3]),.I1(c[4:4]),.I2(m100),.I3(m108),.I4(m182),.O(m183));
defparam desc2955.INIT=32'hDCFE1032;
  LUT6 desc2956(.I0(c[2:2]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m156),.I5(m176),.O(m177));
defparam desc2956.INIT=64'hFFF8F7F00F080700;
  LUT5 desc2957(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m100),.I4(m108),.O(m162));
defparam desc2957.INIT=32'h8BCF0347;
  LUT6 desc2958(.I0(c[2:2]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m156),.I5(m157),.O(m160));
defparam desc2958.INIT=64'hFFC0BF807F403F00;
  LUT5 desc2959(.I0(c[3:3]),.I1(c[4:4]),.I2(N_83_0),.I3(N_86_0),.I4(m125),.O(m126));
defparam desc2959.INIT=32'hFEDC3210;
  LUT5 desc2960(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(N_89_0),.I4(m121),.O(m122));
defparam desc2960.INIT=32'hFEDC3210;
  LUT6 desc2961(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m100),.I4(m115),.I5(m108),.O(m117));
defparam desc2961.INIT=64'hBA983210FEDC7654;
  LUT6 desc2962(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(N_83_0),.I4(N_96_0),.I5(N_86_0),.O(m97));
defparam desc2962.INIT=64'hFEDC7654BA983210;
  LUT5 desc2963(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m90),.I4(N_89_0),.O(N_93_0));
defparam desc2963.INIT=32'hFC74B830;
  LUT5 desc2964(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(N_83_0),.I4(N_86_0),.O(m87));
defparam desc2964.INIT=32'hFCB87430;
  LUT6 desc2965(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m47),.I4(m57_o5_inv),.I5(N_50_0),.O(m59));
defparam desc2965.INIT=64'hFEDC7654BA983210;
  LUT5 desc2966(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(N_12_1),.I4(m45),.O(N_47_0));
defparam desc2966.INIT=32'hFEDC3210;
  LUT5 desc2967(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(N_12_1),.I4(m26_lut6_2_O6),.O(N_29_0));
defparam desc2967.INIT=32'hFCB87430;
  LUT3 v_r1_2_3_16_cZ(.I0(r0_2[5:5]),.I1(v_r1_2_3_4),.I2(v_r1_2_3_14_0),.O(v_r1_2_3_16));
defparam v_r1_2_3_16_cZ.INIT=8'hA8;
  LUT5 desc2968(.I0(c[3:3]),.I1(c[4:4]),.I2(N_96_0),.I3(m132),.I4(N_86_0),.O(N_2942_i));
defparam desc2968.INIT=32'h31FD20EC;
  LUT5 desc2969(.I0(c[3:3]),.I1(c[4:4]),.I2(m115),.I3(m108),.I4(m141_lut6_2_O6),.O(N_2951_i));
defparam desc2969.INIT=32'h2031ECFD;
  LUT5 desc2970(.I0(c[3:3]),.I1(c[4:4]),.I2(m73_lut6_2_O5),.I3(m57_o5_inv),.I4(N_50_0),.O(N_2895_i));
defparam desc2970.INIT=32'h3F1D2E0C;
  LUT5 v_r1_2_3_0_axb_0_cZ(.I0(c[2:2]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m127_lut6_2_O6),.O(v_r1_2_3_0_axb_0));
defparam v_r1_2_3_0_axb_0_cZ.INIT=32'h01000001;
  LUT5 desc2971(.I0(c[3:3]),.I1(c[4:4]),.I2(m47),.I3(m71_lut6_2_O6),.I4(N_50_0),.O(N_2891_i));
defparam desc2971.INIT=32'h32FE10DC;
  LUT5 desc2972(.I0(c[3:3]),.I1(c[4:4]),.I2(m90),.I3(N_89_0),.I4(m129),.O(N_2939_i));
defparam desc2972.INIT=32'h3120FDEC;
  LUT5 desc2973(.I0(c[3:3]),.I1(c[4:4]),.I2(N_12_1),.I3(m26_lut6_2_O6),.I4(m67),.O(N_2887_i));
defparam desc2973.INIT=32'h3210FEDC;
  LUT6 v_r1_2_3_0_axb_51_cZ(.I0(r0_2[51:51]),.I1(c[3:3]),.I2(c[4:4]),.I3(un14_s_state_cry[50:50]),.I4(m200),.I5(v_r1_2_3_175),.O(v_r1_2_3_0_axb_51));
defparam v_r1_2_3_0_axb_51_cZ.INIT=64'hAA956A55556A95AA;
  LUT5 v_r1_2_3_21_2_cZ(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(v_r1_2_3_4),.I4(v_r1_2_3_14_0),.O(v_r1_2_3_21_2));
defparam v_r1_2_3_21_2_cZ.INIT=32'hE8E8E888;
  LUT6_L s_ine_o_e(.I0(s_ine_o),.I1(un3_s_count_0_a2_lut6_2_O6),.I2(un31_s_count_0_I_139),.I3(un33_s_count_NE_1_4),.I4(un33_s_count_NE_8),.I5(un33_s_count_NE_2_4),.LO(s_ine_o_0));
defparam s_ine_o_e.INIT=64'h2E2E2E2E2E2E2E22;
  LUT6 v_r1_2_3_23_cZ(.I0(b_2[6:6]),.I1(r0_2[6:6]),.I2(r0_2[5:5]),.I3(r0_2[7:7]),.I4(v_r1_2_3_4),.I5(v_r1_2_3_14_0),.O(v_r1_2_3_23));
defparam v_r1_2_3_23_cZ.INIT=64'hE800E800E8008800;
  LUT6 v_r1_2_3_35_0_cZ(.I0(b_2[10:10]),.I1(b_2[8:8]),.I2(r0_2[10:10]),.I3(r0_2[9:9]),.I4(v_r1_2_3_10),.I5(v_r1_2_3_28_0_tz),.O(v_r1_2_3_35_0));
defparam v_r1_2_3_35_0_cZ.INIT=64'hAAA0A8A0AAA0A0A0;
  LUT6 v_r1_2_3_49_cZ(.I0(r0_2[14:14]),.I1(b_2[14:14]),.I2(r0_2[13:13]),.I3(v_r1_2_3_41_0),.I4(b_2_RNIMF314[10:10]),.I5(v_r1_2_3_42_0),.O(v_r1_2_3_49));
defparam v_r1_2_3_49_cZ.INIT=64'hE8E8E8E8E8888888;
  LUT5 v_r1_2_3_63_0_c_cZ(.I0(b_2[18:18]),.I1(r0_2[16:16]),.I2(r0_2[17:17]),.I3(r0_2[15:15]),.I4(v_r1_2_3_49),.O(v_r1_2_3_63_0_c));
defparam v_r1_2_3_63_0_c_cZ.INIT=32'h80000000;
  LUT5_L v_r1_2_3_56_cZ(.I0(b_2[16:16]),.I1(r0_2[16:16]),.I2(r0_2[15:15]),.I3(v_r1_2_3_49),.I4(v_r1_2_3_56_0_tz),.LO(v_r1_2_3_56));
defparam v_r1_2_3_56_cZ.INIT=32'hEAAAC000;
  LUT5 v_r1_2_3_63_tz_0_0(.I0(b_2[18:18]),.I1(r0_2[18:18]),.I2(b_2[16:16]),.I3(r0_2[17:17]),.I4(v_r1_2_3_56_0_tz),.O(v_r1_2_3_63_0_d));
defparam v_r1_2_3_63_tz_0_0.INIT=32'hA8888888;
  LUT5 v_r1_2_3_62(.I0(r0_2[18:18]),.I1(b_2[16:16]),.I2(r0_2[17:17]),.I3(v_r1_2_3_22),.I4(v_r1_2_3_56_0_tz),.O(v_r1_2_3_25));
defparam v_r1_2_3_62.INIT=32'hA080A000;
  LUT6 v_r1_2_3_63_2_0_cZ(.I0(b_2[18:18]),.I1(r0_2[18:18]),.I2(b_2[16:16]),.I3(r0_2[17:17]),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.O(v_r1_2_3_63_2_0));
defparam v_r1_2_3_63_2_0_cZ.INIT=64'hAA88A888AA888888;
  LUT6_L v_r1_2_3_63_2_cZ(.I0(b_2[18:18]),.I1(r0_2[18:18]),.I2(b_2[16:16]),.I3(r0_2[17:17]),.I4(v_r1_2_3_22),.I5(v_r1_2_3_56_0_tz),.LO(v_r1_2_3_63_2));
defparam v_r1_2_3_63_2_cZ.INIT=64'hEE88E888EE888888;
  LUT5 v_r1_2_3_7_RNIQJM46(.I0(r0_2[3:3]),.I1(c[4:4]),.I2(v_r1_2_3_7),.I3(un14_s_state_cry[50:50]),.I4(m141_lut6_2_O5),.O(v_r1_2_3_0_axb_3));
defparam v_r1_2_3_7_RNIQJM46.INIT=32'h965AA569;
  LUT5 v_r1_2_3_14_RNIE7KT4(.I0(r0_2[5:5]),.I1(c[4:4]),.I2(v_r1_2_3_14),.I3(un14_s_state_cry[50:50]),.I4(m191),.O(v_r1_2_3_0_axb_5));
defparam v_r1_2_3_14_RNIE7KT4.INIT=32'h965AA569;
  LUT2 v_r1_2_3_0_cry_5_RNO_cZ(.I0(r0_2[5:5]),.I1(v_r1_2_3_14),.O(v_r1_2_3_0_cry_5_RNO));
defparam v_r1_2_3_0_cry_5_RNO_cZ.INIT=4'h6;
  LUT5 v_r1_2_3_21_2_RNIR2D76(.I0(r0_2[7:7]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(v_r1_2_3_21_2),.I4(m141_lut6_2_O6),.O(v_r1_2_3_0_axb_7));
defparam v_r1_2_3_21_2_RNIR2D76.INIT=32'h956AA659;
  LUT5 desc2974(.I0(r0_2[9:9]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(v_r1_2_3_21_2_RNIMLGQ),.I4(m189),.O(v_r1_2_3_0_axb_9));
defparam desc2974.INIT=32'h956AA659;
  LUT5 desc2975(.I0(r0_2[11:11]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(b_2_RNIMF314[10:10]),.I4(m210),.O(v_r1_2_3_0_axb_11));
defparam desc2975.INIT=32'h956AA659;
  LUT2 v_r1_2_3_0_cry_11_RNO_cZ(.I0(r0_2[11:11]),.I1(b_2_RNIMF314[10:10]),.O(v_r1_2_3_0_cry_11_RNO));
defparam v_r1_2_3_0_cry_11_RNO_cZ.INIT=4'h6;
  LUT5 desc2976(.I0(r0_2[13:13]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(v_r1_2_3_35_0_RNIKOE74),.I4(m186),.O(v_r1_2_3_0_axb_13));
defparam desc2976.INIT=32'h956AA659;
  LUT2 v_r1_2_3_0_cry_13_RNO_cZ(.I0(r0_2[13:13]),.I1(v_r1_2_3_35_0_RNIKOE74),.O(v_r1_2_3_0_cry_13_RNO));
defparam v_r1_2_3_0_cry_13_RNO_cZ.INIT=4'h6;
  LUT5 v_r1_2_3_49_RNIAKEIA(.I0(r0_2[15:15]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m182),.I4(v_r1_2_3_49),.O(v_r1_2_3_0_axb_15));
defparam v_r1_2_3_49_RNIAKEIA.INIT=32'hA695596A;
  LUT2 v_r1_2_3_0_cry_15_RNO_cZ(.I0(r0_2[15:15]),.I1(v_r1_2_3_49),.O(v_r1_2_3_0_cry_15_RNO));
defparam v_r1_2_3_0_cry_15_RNO_cZ.INIT=4'h6;
  LUT5 v_r1_2_3_56_RNI26FIC(.I0(r0_2[17:17]),.I1(c[4:4]),.I2(m193),.I3(m180),.I4(v_r1_2_3_56),.O(v_r1_2_3_0_axb_17));
defparam v_r1_2_3_56_RNI26FIC.INIT=32'h6A5995A6;
  LUT5 v_r1_2_3_63_tz_0_0_RNIQEK1E(.I0(r0_2[19:19]),.I1(N_3022_i),.I2(v_r1_2_3_63_0_c),.I3(v_r1_2_3_63_0_d),.I4(v_r1_2_3_25),.O(v_r1_2_3_0_axb_19));
defparam v_r1_2_3_63_tz_0_0_RNIQEK1E.INIT=32'h99999996;
  LUT4 v_r1_2_3_0_cry_19_RNO_cZ(.I0(r0_2[19:19]),.I1(v_r1_2_3_63_0_c),.I2(v_r1_2_3_63_0_d),.I3(v_r1_2_3_25),.O(v_r1_2_3_0_cry_19_RNO));
defparam v_r1_2_3_0_cry_19_RNO_cZ.INIT=16'h5556;
  LUT5 desc2977(.I0(r0_2[23:23]),.I1(b_2[22:22]),.I2(N_2951_i),.I3(v_r1_2_3_31),.I4(v_r1_2_3_77_0_tz),.O(v_r1_2_3_0_axb_23));
defparam desc2977.INIT=32'hA596A55A;
  LUT4 v_r1_2_3_0_cry_23_RNO_cZ(.I0(r0_2[23:23]),.I1(b_2[22:22]),.I2(v_r1_2_3_31),.I3(v_r1_2_3_77_0_tz),.O(v_r1_2_3_0_cry_23_RNO));
defparam v_r1_2_3_0_cry_23_RNO_cZ.INIT=16'h565A;
  LUT3 v_r1_2_3_0_cry_24_RNO_cZ(.I0(b_2[24:24]),.I1(r0_2[24:24]),.I2(v_r1_2_3_73_0_lut6_2_RNIM5CP22),.O(v_r1_2_3_0_cry_24_RNO));
defparam v_r1_2_3_0_cry_24_RNO_cZ.INIT=8'h96;
  LUT5 desc2978(.I0(b_2[26:26]),.I1(r0_2[25:25]),.I2(r0_2[26:26]),.I3(N_2891_i),.I4(m190_lut6_2_O6),.O(v_r1_2_3_0_axb_26));
defparam desc2978.INIT=32'hA55A6996;
  LUT5 desc2979(.I0(b_2[28:28]),.I1(r0_2[28:28]),.I2(r0_2[27:27]),.I3(m211),.I4(N_2939_i),.O(v_r1_2_3_0_axb_28));
defparam desc2979.INIT=32'h99696696;
  LUT5 desc2980(.I0(b_2[28:28]),.I1(r0_2[28:28]),.I2(r0_2[29:29]),.I3(N_2939_i),.I4(m187_lut6_2_O6),.O(v_r1_2_3_0_axb_29));
defparam desc2980.INIT=32'h1E78E187;
  LUT5 desc2981(.I0(b_2[30:30]),.I1(r0_2[30:30]),.I2(r0_2[29:29]),.I3(N_2887_i),.I4(m187_lut6_2_O6),.O(v_r1_2_3_0_axb_30));
defparam desc2981.INIT=32'h99666996;
  LUT5 desc2982(.I0(b_2[30:30]),.I1(r0_2[30:30]),.I2(r0_2[31:31]),.I3(N_2887_i),.I4(m183),.O(v_r1_2_3_0_axb_31));
defparam desc2982.INIT=32'hE1871E78;
  LUT5 desc2983(.I0(b_2[32:32]),.I1(r0_2[32:32]),.I2(r0_2[31:31]),.I3(m126),.I4(m183),.O(v_r1_2_3_0_axb_32));
defparam desc2983.INIT=32'h69969966;
  LUT5 desc2984(.I0(b_2[32:32]),.I1(r0_2[32:32]),.I2(r0_2[33:33]),.I3(m126),.I4(N_48_i_lut6_2_O5),.O(v_r1_2_3_0_axb_33));
defparam desc2984.INIT=32'hE1871E78;
  LUT5 desc2985(.I0(b_2[34:34]),.I1(r0_2[34:34]),.I2(r0_2[33:33]),.I3(m59),.I4(N_48_i_lut6_2_O5),.O(v_r1_2_3_0_axb_34));
defparam desc2985.INIT=32'h69969966;
  LUT5 desc2986(.I0(b_2[34:34]),.I1(r0_2[34:34]),.I2(r0_2[35:35]),.I3(m59),.I4(m208),.O(v_r1_2_3_0_axb_35));
defparam desc2986.INIT=32'hE1871E78;
  LUT5 desc2987(.I0(b_2[36:36]),.I1(r0_2[36:36]),.I2(r0_2[35:35]),.I3(m122),.I4(m208),.O(v_r1_2_3_0_axb_36));
defparam desc2987.INIT=32'h69969966;
  LUT5 desc2988(.I0(b_2[36:36]),.I1(r0_2[36:36]),.I2(r0_2[37:37]),.I3(m122),.I4(m177),.O(v_r1_2_3_0_axb_37));
defparam desc2988.INIT=32'hE1871E78;
  LUT2 v_r1_2_3_0_cry_37_RNO_cZ(.I0(r0_2[37:37]),.I1(m177),.O(v_r1_2_3_0_cry_37_RNO));
defparam v_r1_2_3_0_cry_37_RNO_cZ.INIT=4'h6;
  LUT5 desc2989(.I0(b_2[38:38]),.I1(r0_2[38:38]),.I2(r0_2[37:37]),.I3(N_47_0),.I4(m177),.O(v_r1_2_3_0_axb_38));
defparam desc2989.INIT=32'h69969966;
  LUT2 v_r1_2_3_0_cry_38_RNO_cZ(.I0(r0_2[37:37]),.I1(m177),.O(v_r1_2_3_0_cry_38_RNO));
defparam v_r1_2_3_0_cry_38_RNO_cZ.INIT=4'h8;
  LUT5 desc2990(.I0(b_2[38:38]),.I1(r0_2[38:38]),.I2(r0_2[39:39]),.I3(m117),.I4(N_47_0),.O(v_r1_2_3_0_axb_39));
defparam desc2990.INIT=32'hE11E8778;
  LUT2 v_r1_2_3_0_cry_39_RNO_cZ(.I0(r0_2[39:39]),.I1(m117),.O(v_r1_2_3_0_cry_39_RNO));
defparam v_r1_2_3_0_cry_39_RNO_cZ.INIT=4'h6;
  LUT5 desc2991(.I0(b_2[40:40]),.I1(r0_2[40:40]),.I2(r0_2[39:39]),.I3(m97),.I4(m117),.O(v_r1_2_3_0_axb_40));
defparam desc2991.INIT=32'h69969966;
  LUT2 v_r1_2_3_0_cry_40_RNO_cZ(.I0(r0_2[39:39]),.I1(m117),.O(v_r1_2_3_0_cry_40_RNO));
defparam v_r1_2_3_0_cry_40_RNO_cZ.INIT=4'h8;
  LUT5 desc2992(.I0(b_2[40:40]),.I1(r0_2[40:40]),.I2(r0_2[41:41]),.I3(m97),.I4(m190_lut6_2_O5),.O(v_r1_2_3_0_axb_41));
defparam desc2992.INIT=32'hE1871E78;
  LUT5 desc2993(.I0(b_2[42:42]),.I1(r0_2[42:42]),.I2(r0_2[41:41]),.I3(m168_lut6_2_O6),.I4(m190_lut6_2_O5),.O(v_r1_2_3_0_axb_42));
defparam desc2993.INIT=32'h69969966;
  LUT5 desc2994(.I0(b_2[42:42]),.I1(r0_2[42:42]),.I2(r0_2[43:43]),.I3(m205),.I4(m168_lut6_2_O6),.O(v_r1_2_3_0_axb_43));
defparam desc2994.INIT=32'hE11E8778;
  LUT5 desc2995(.I0(b_2[44:44]),.I1(r0_2[44:44]),.I2(r0_2[43:43]),.I3(N_93_0),.I4(m205),.O(v_r1_2_3_0_axb_44));
defparam desc2995.INIT=32'h69969966;
  LUT5 desc2996(.I0(b_2[44:44]),.I1(r0_2[44:44]),.I2(r0_2[45:45]),.I3(N_93_0),.I4(m187_lut6_2_O5),.O(v_r1_2_3_0_axb_45));
defparam desc2996.INIT=32'hE1871E78;
  LUT5 desc2997(.I0(b_2[46:46]),.I1(r0_2[46:46]),.I2(r0_2[45:45]),.I3(N_29_0),.I4(m187_lut6_2_O5),.O(v_r1_2_3_0_axb_46));
defparam desc2997.INIT=32'h69969966;
  LUT5 desc2998(.I0(b_2[46:46]),.I1(r0_2[46:46]),.I2(r0_2[47:47]),.I3(m162),.I4(N_29_0),.O(v_r1_2_3_0_axb_47));
defparam desc2998.INIT=32'h1EE17887;
  LUT5 desc2999(.I0(b_2[48:48]),.I1(r0_2[48:48]),.I2(r0_2[47:47]),.I3(m162),.I4(m87),.O(v_r1_2_3_0_axb_48));
defparam desc2999.INIT=32'h99696696;
  LUT5 desc3000(.I0(b_2[48:48]),.I1(r0_2[48:48]),.I2(r0_2[49:49]),.I3(m160),.I4(m87),.O(v_r1_2_3_0_axb_49));
defparam desc3000.INIT=32'hE11E8778;
  LUT2 v_r1_2_3_0_cry_49_RNO_cZ(.I0(r0_2[49:49]),.I1(m160),.O(v_r1_2_3_0_cry_49_RNO));
defparam v_r1_2_3_0_cry_49_RNO_cZ.INIT=4'h6;
  LUT5 desc3001(.I0(b_2[50:50]),.I1(r0_2[50:50]),.I2(r0_2[49:49]),.I3(m160),.I4(m168_lut6_2_O5),.O(v_r1_2_3_0_axb_50));
defparam desc3001.INIT=32'h69999666;
  LUT2 v_r1_2_3_0_cry_50_RNO_cZ(.I0(r0_2[49:49]),.I1(m160),.O(v_r1_2_3_0_cry_50_RNO));
defparam v_r1_2_3_0_cry_50_RNO_cZ.INIT=4'h8;
  LUT2 un33_s_count_a_5_0_cry_26_RNO_cZ(.I0(r1[24:24]),.I1(r1_2[25:25]),.O(un33_s_count_a_5_0_cry_26_RNO));
defparam un33_s_count_a_5_0_cry_26_RNO_cZ.INIT=4'hD;
  LUT2 un33_s_count_a_5_0_cry_28_RNO_cZ(.I0(r1_2[27:27]),.I1(s_rad_i[27:27]),.O(un33_s_count_a_5_0_cry_28_RNO));
defparam un33_s_count_a_5_0_cry_28_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_29_RNO_cZ(.I0(r1_2[28:28]),.I1(s_rad_i[28:28]),.O(un33_s_count_a_5_0_cry_29_RNO));
defparam un33_s_count_a_5_0_cry_29_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_30_RNO_cZ(.I0(r1_2[29:29]),.I1(s_rad_i[29:29]),.O(un33_s_count_a_5_0_cry_30_RNO));
defparam un33_s_count_a_5_0_cry_30_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_31_RNO_cZ(.I0(r1_2[30:30]),.I1(s_rad_i[30:30]),.O(un33_s_count_a_5_0_cry_31_RNO));
defparam un33_s_count_a_5_0_cry_31_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_32_RNO_cZ(.I0(r1_2[31:31]),.I1(s_rad_i[31:31]),.O(un33_s_count_a_5_0_cry_32_RNO));
defparam un33_s_count_a_5_0_cry_32_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_33_RNO_cZ(.I0(r1_2[32:32]),.I1(s_rad_i[32:32]),.O(un33_s_count_a_5_0_cry_33_RNO));
defparam un33_s_count_a_5_0_cry_33_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_34_RNO_cZ(.I0(r1_2[33:33]),.I1(s_rad_i[33:33]),.O(un33_s_count_a_5_0_cry_34_RNO));
defparam un33_s_count_a_5_0_cry_34_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_35_RNO_cZ(.I0(r1_2[34:34]),.I1(s_rad_i[34:34]),.O(un33_s_count_a_5_0_cry_35_RNO));
defparam un33_s_count_a_5_0_cry_35_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_36_RNO_cZ(.I0(r1_2[35:35]),.I1(s_rad_i[35:35]),.O(un33_s_count_a_5_0_cry_36_RNO));
defparam un33_s_count_a_5_0_cry_36_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_37_RNO_cZ(.I0(r1_2[36:36]),.I1(s_rad_i[36:36]),.O(un33_s_count_a_5_0_cry_37_RNO));
defparam un33_s_count_a_5_0_cry_37_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_38_RNO_cZ(.I0(r1_2[37:37]),.I1(s_rad_i[37:37]),.O(un33_s_count_a_5_0_cry_38_RNO));
defparam un33_s_count_a_5_0_cry_38_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_39_RNO_cZ(.I0(r1_2[38:38]),.I1(s_rad_i[38:38]),.O(un33_s_count_a_5_0_cry_39_RNO));
defparam un33_s_count_a_5_0_cry_39_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_40_RNO_cZ(.I0(r1_2[39:39]),.I1(s_rad_i[39:39]),.O(un33_s_count_a_5_0_cry_40_RNO));
defparam un33_s_count_a_5_0_cry_40_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_41_RNO_cZ(.I0(r1_2[40:40]),.I1(s_rad_i[40:40]),.O(un33_s_count_a_5_0_cry_41_RNO));
defparam un33_s_count_a_5_0_cry_41_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_42_RNO_cZ(.I0(r1_2[41:41]),.I1(s_rad_i[41:41]),.O(un33_s_count_a_5_0_cry_42_RNO));
defparam un33_s_count_a_5_0_cry_42_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_43_RNO_cZ(.I0(r1_2[42:42]),.I1(s_rad_i[42:42]),.O(un33_s_count_a_5_0_cry_43_RNO));
defparam un33_s_count_a_5_0_cry_43_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_44_RNO_cZ(.I0(r1_2[43:43]),.I1(s_rad_i[43:43]),.O(un33_s_count_a_5_0_cry_44_RNO));
defparam un33_s_count_a_5_0_cry_44_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_45_RNO_cZ(.I0(r1_2[44:44]),.I1(s_rad_i[44:44]),.O(un33_s_count_a_5_0_cry_45_RNO));
defparam un33_s_count_a_5_0_cry_45_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_46_RNO_cZ(.I0(r1_2[45:45]),.I1(s_rad_i[45:45]),.O(un33_s_count_a_5_0_cry_46_RNO));
defparam un33_s_count_a_5_0_cry_46_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_47_RNO_cZ(.I0(r1_2[46:46]),.I1(s_rad_i[46:46]),.O(un33_s_count_a_5_0_cry_47_RNO));
defparam un33_s_count_a_5_0_cry_47_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_48_RNO_cZ(.I0(r1_2[47:47]),.I1(s_rad_i[47:47]),.O(un33_s_count_a_5_0_cry_48_RNO));
defparam un33_s_count_a_5_0_cry_48_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_49_RNO_cZ(.I0(r1_2[48:48]),.I1(s_rad_i[48:48]),.O(un33_s_count_a_5_0_cry_49_RNO));
defparam un33_s_count_a_5_0_cry_49_RNO_cZ.INIT=4'h2;
  LUT2 un33_s_count_a_5_0_cry_50_RNO_cZ(.I0(r1_2[49:49]),.I1(s_rad_i[49:49]),.O(un33_s_count_a_5_0_cry_50_RNO));
defparam un33_s_count_a_5_0_cry_50_RNO_cZ.INIT=4'h2;
  XORCY un1_r1_s_24_cZ(.LI(un1_r1_axb_24),.CI(un1_r1_cry_23),.O(un1_r1_s_24));
  XORCY un1_r1_s_23_cZ(.LI(un1_r1_axb_23),.CI(un1_r1_cry_22),.O(un1_r1_s_23));
  MUXCY_L un1_r1_cry_23_cZ(.DI(r1[23:23]),.CI(un1_r1_cry_22),.S(un1_r1_axb_23),.LO(un1_r1_cry_23));
  XORCY un1_r1_s_22_cZ(.LI(un1_r1_axb_22),.CI(un1_r1_cry_21),.O(un1_r1_s_22));
  MUXCY_L un1_r1_cry_22_cZ(.DI(r1[22:22]),.CI(un1_r1_cry_21),.S(un1_r1_axb_22),.LO(un1_r1_cry_22));
  XORCY un1_r1_s_21_cZ(.LI(un1_r1_axb_21),.CI(un1_r1_cry_20),.O(un1_r1_s_21));
  MUXCY_L un1_r1_cry_21_cZ(.DI(r1[21:21]),.CI(un1_r1_cry_20),.S(un1_r1_axb_21),.LO(un1_r1_cry_21));
  XORCY un1_r1_s_20_cZ(.LI(un1_r1_axb_20),.CI(un1_r1_cry_19),.O(un1_r1_s_20));
  MUXCY_L un1_r1_cry_20_cZ(.DI(r1[20:20]),.CI(un1_r1_cry_19),.S(un1_r1_axb_20),.LO(un1_r1_cry_20));
  XORCY un1_r1_s_19_cZ(.LI(un1_r1_axb_19),.CI(un1_r1_cry_18),.O(un1_r1_s_19));
  MUXCY_L un1_r1_cry_19_cZ(.DI(r1[19:19]),.CI(un1_r1_cry_18),.S(un1_r1_axb_19),.LO(un1_r1_cry_19));
  XORCY un1_r1_s_18_cZ(.LI(un1_r1_axb_18),.CI(un1_r1_cry_17),.O(un1_r1_s_18));
  MUXCY_L un1_r1_cry_18_cZ(.DI(r1[18:18]),.CI(un1_r1_cry_17),.S(un1_r1_axb_18),.LO(un1_r1_cry_18));
  XORCY un1_r1_s_17_cZ(.LI(un1_r1_axb_17),.CI(un1_r1_cry_16),.O(un1_r1_s_17));
  MUXCY_L un1_r1_cry_17_cZ(.DI(r1[17:17]),.CI(un1_r1_cry_16),.S(un1_r1_axb_17),.LO(un1_r1_cry_17));
  XORCY un1_r1_s_16_cZ(.LI(un1_r1_axb_16),.CI(un1_r1_cry_15),.O(un1_r1_s_16));
  MUXCY_L un1_r1_cry_16_cZ(.DI(r1[16:16]),.CI(un1_r1_cry_15),.S(un1_r1_axb_16),.LO(un1_r1_cry_16));
  XORCY un1_r1_s_15_cZ(.LI(un1_r1_axb_15),.CI(un1_r1_cry_14),.O(un1_r1_s_15));
  MUXCY_L un1_r1_cry_15_cZ(.DI(r1[15:15]),.CI(un1_r1_cry_14),.S(un1_r1_axb_15),.LO(un1_r1_cry_15));
  XORCY un1_r1_s_14_cZ(.LI(un1_r1_axb_14),.CI(un1_r1_cry_13),.O(un1_r1_s_14));
  MUXCY_L un1_r1_cry_14_cZ(.DI(r1[14:14]),.CI(un1_r1_cry_13),.S(un1_r1_axb_14),.LO(un1_r1_cry_14));
  XORCY un1_r1_s_13_cZ(.LI(un1_r1_axb_13),.CI(un1_r1_cry_12),.O(un1_r1_s_13));
  MUXCY_L un1_r1_cry_13_cZ(.DI(r1[13:13]),.CI(un1_r1_cry_12),.S(un1_r1_axb_13),.LO(un1_r1_cry_13));
  XORCY un1_r1_s_12_cZ(.LI(un1_r1_axb_12),.CI(un1_r1_cry_11),.O(un1_r1_s_12));
  MUXCY_L un1_r1_cry_12_cZ(.DI(r1[12:12]),.CI(un1_r1_cry_11),.S(un1_r1_axb_12),.LO(un1_r1_cry_12));
  XORCY un1_r1_s_11_cZ(.LI(un1_r1_axb_11),.CI(un1_r1_cry_10),.O(un1_r1_s_11));
  MUXCY_L un1_r1_cry_11_cZ(.DI(r1[11:11]),.CI(un1_r1_cry_10),.S(un1_r1_axb_11),.LO(un1_r1_cry_11));
  XORCY un1_r1_s_10_cZ(.LI(un1_r1_axb_10),.CI(un1_r1_cry_9),.O(un1_r1_s_10));
  MUXCY_L un1_r1_cry_10_cZ(.DI(r1[10:10]),.CI(un1_r1_cry_9),.S(un1_r1_axb_10),.LO(un1_r1_cry_10));
  XORCY un1_r1_s_9_cZ(.LI(un1_r1_axb_9),.CI(un1_r1_cry_8),.O(un1_r1_s_9));
  MUXCY_L un1_r1_cry_9_cZ(.DI(r1[9:9]),.CI(un1_r1_cry_8),.S(un1_r1_axb_9),.LO(un1_r1_cry_9));
  XORCY un1_r1_s_8_cZ(.LI(un1_r1_axb_8),.CI(un1_r1_cry_7),.O(un1_r1_s_8));
  MUXCY_L un1_r1_cry_8_cZ(.DI(r1[8:8]),.CI(un1_r1_cry_7),.S(un1_r1_axb_8),.LO(un1_r1_cry_8));
  XORCY un1_r1_s_7_cZ(.LI(un1_r1_axb_7),.CI(un1_r1_cry_6),.O(un1_r1_s_7));
  MUXCY_L un1_r1_cry_7_cZ(.DI(r1[7:7]),.CI(un1_r1_cry_6),.S(un1_r1_axb_7),.LO(un1_r1_cry_7));
  XORCY un1_r1_s_6_cZ(.LI(un1_r1_axb_6),.CI(un1_r1_cry_5),.O(un1_r1_s_6));
  MUXCY_L un1_r1_cry_6_cZ(.DI(r1[6:6]),.CI(un1_r1_cry_5),.S(un1_r1_axb_6),.LO(un1_r1_cry_6));
  XORCY un1_r1_s_5_cZ(.LI(un1_r1_axb_5),.CI(un1_r1_cry_4),.O(un1_r1_s_5));
  MUXCY_L un1_r1_cry_5_cZ(.DI(r1[5:5]),.CI(un1_r1_cry_4),.S(un1_r1_axb_5),.LO(un1_r1_cry_5));
  XORCY un1_r1_s_4_cZ(.LI(un1_r1_axb_4),.CI(un1_r1_cry_3),.O(un1_r1_s_4));
  MUXCY_L un1_r1_cry_4_cZ(.DI(r1[4:4]),.CI(un1_r1_cry_3),.S(un1_r1_axb_4),.LO(un1_r1_cry_4));
  XORCY un1_r1_s_3_cZ(.LI(un1_r1_axb_3),.CI(un1_r1_cry_2),.O(un1_r1_s_3));
  MUXCY_L un1_r1_cry_3_cZ(.DI(r1[3:3]),.CI(un1_r1_cry_2),.S(un1_r1_axb_3),.LO(un1_r1_cry_3));
  XORCY un1_r1_s_2_cZ(.LI(un1_r1_axb_2),.CI(un1_r1_cry_1),.O(un1_r1_s_2));
  MUXCY_L un1_r1_cry_2_cZ(.DI(r1[2:2]),.CI(un1_r1_cry_1),.S(un1_r1_axb_2),.LO(un1_r1_cry_2));
  XORCY un1_r1_s_1_cZ(.LI(un1_r1_axb_1),.CI(un1_r1_cry_0),.O(un1_r1_s_1));
  MUXCY_L un1_r1_cry_1_cZ(.DI(r1[1:1]),.CI(un1_r1_cry_0),.S(un1_r1_axb_1),.LO(un1_r1_cry_1));
  MUXCY_L un1_r1_cry_0_cZ(.DI(r1[0:0]),.CI(GND),.S(un1_r1_axb_0),.LO(un1_r1_cry_0));
  XORCY v_r1_3_s_25(.LI(v_r1_3_axb_25),.CI(v_r1_3_cry_24),.O(v_r1_3[25:25]));
  XORCY v_r1_3_s_24(.LI(v_r1_3_axb_24),.CI(v_r1_3_cry_23),.O(v_r1_3[24:24]));
  MUXCY_L v_r1_3_cry_24_cZ(.DI(r0[24:24]),.CI(v_r1_3_cry_23),.S(v_r1_3_axb_24),.LO(v_r1_3_cry_24));
  XORCY v_r1_3_s_23(.LI(v_r1_3_axb_23),.CI(v_r1_3_cry_22),.O(v_r1_3[23:23]));
  MUXCY_L v_r1_3_cry_23_cZ(.DI(r0[23:23]),.CI(v_r1_3_cry_22),.S(v_r1_3_axb_23),.LO(v_r1_3_cry_23));
  XORCY v_r1_3_s_22(.LI(v_r1_3_axb_22),.CI(v_r1_3_cry_21),.O(v_r1_3[22:22]));
  MUXCY_L v_r1_3_cry_22_cZ(.DI(r0[22:22]),.CI(v_r1_3_cry_21),.S(v_r1_3_axb_22),.LO(v_r1_3_cry_22));
  XORCY v_r1_3_s_21(.LI(v_r1_3_axb_21),.CI(v_r1_3_cry_20),.O(v_r1_3[21:21]));
  MUXCY_L v_r1_3_cry_21_cZ(.DI(r0[21:21]),.CI(v_r1_3_cry_20),.S(v_r1_3_axb_21),.LO(v_r1_3_cry_21));
  XORCY v_r1_3_s_20(.LI(v_r1_3_axb_20),.CI(v_r1_3_cry_19),.O(v_r1_3[20:20]));
  MUXCY_L v_r1_3_cry_20_cZ(.DI(r0[20:20]),.CI(v_r1_3_cry_19),.S(v_r1_3_axb_20),.LO(v_r1_3_cry_20));
  XORCY v_r1_3_s_19(.LI(v_r1_3_axb_19),.CI(v_r1_3_cry_18),.O(v_r1_3[19:19]));
  MUXCY_L v_r1_3_cry_19_cZ(.DI(r0[19:19]),.CI(v_r1_3_cry_18),.S(v_r1_3_axb_19),.LO(v_r1_3_cry_19));
  XORCY v_r1_3_s_18(.LI(v_r1_3_axb_18),.CI(v_r1_3_cry_17),.O(v_r1_3[18:18]));
  MUXCY_L v_r1_3_cry_18_cZ(.DI(r0[18:18]),.CI(v_r1_3_cry_17),.S(v_r1_3_axb_18),.LO(v_r1_3_cry_18));
  XORCY v_r1_3_s_17(.LI(v_r1_3_axb_17),.CI(v_r1_3_cry_16),.O(v_r1_3[17:17]));
  MUXCY_L v_r1_3_cry_17_cZ(.DI(r0[17:17]),.CI(v_r1_3_cry_16),.S(v_r1_3_axb_17),.LO(v_r1_3_cry_17));
  XORCY v_r1_3_s_16(.LI(v_r1_3_axb_16),.CI(v_r1_3_cry_15),.O(v_r1_3[16:16]));
  MUXCY_L v_r1_3_cry_16_cZ(.DI(r0[16:16]),.CI(v_r1_3_cry_15),.S(v_r1_3_axb_16),.LO(v_r1_3_cry_16));
  XORCY v_r1_3_s_15(.LI(v_r1_3_axb_15),.CI(v_r1_3_cry_14),.O(v_r1_3[15:15]));
  MUXCY_L v_r1_3_cry_15_cZ(.DI(r0[15:15]),.CI(v_r1_3_cry_14),.S(v_r1_3_axb_15),.LO(v_r1_3_cry_15));
  XORCY v_r1_3_s_14(.LI(v_r1_3_axb_14),.CI(v_r1_3_cry_13),.O(v_r1_3[14:14]));
  MUXCY_L v_r1_3_cry_14_cZ(.DI(r0[14:14]),.CI(v_r1_3_cry_13),.S(v_r1_3_axb_14),.LO(v_r1_3_cry_14));
  XORCY v_r1_3_s_13(.LI(v_r1_3_axb_13),.CI(v_r1_3_cry_12),.O(v_r1_3[13:13]));
  MUXCY_L v_r1_3_cry_13_cZ(.DI(r0[13:13]),.CI(v_r1_3_cry_12),.S(v_r1_3_axb_13),.LO(v_r1_3_cry_13));
  XORCY v_r1_3_s_12(.LI(v_r1_3_axb_12),.CI(v_r1_3_cry_11),.O(v_r1_3[12:12]));
  MUXCY_L v_r1_3_cry_12_cZ(.DI(r0[12:12]),.CI(v_r1_3_cry_11),.S(v_r1_3_axb_12),.LO(v_r1_3_cry_12));
  XORCY v_r1_3_s_11(.LI(v_r1_3_axb_11),.CI(v_r1_3_cry_10),.O(v_r1_3[11:11]));
  MUXCY_L v_r1_3_cry_11_cZ(.DI(r0[11:11]),.CI(v_r1_3_cry_10),.S(v_r1_3_axb_11),.LO(v_r1_3_cry_11));
  XORCY v_r1_3_s_10(.LI(v_r1_3_axb_10),.CI(v_r1_3_cry_9),.O(v_r1_3[10:10]));
  MUXCY_L v_r1_3_cry_10_cZ(.DI(r0[10:10]),.CI(v_r1_3_cry_9),.S(v_r1_3_axb_10),.LO(v_r1_3_cry_10));
  XORCY v_r1_3_s_9(.LI(v_r1_3_axb_9),.CI(v_r1_3_cry_8),.O(v_r1_3[9:9]));
  MUXCY_L v_r1_3_cry_9_cZ(.DI(r0[9:9]),.CI(v_r1_3_cry_8),.S(v_r1_3_axb_9),.LO(v_r1_3_cry_9));
  XORCY v_r1_3_s_8(.LI(v_r1_3_axb_8),.CI(v_r1_3_cry_7),.O(v_r1_3[8:8]));
  MUXCY_L v_r1_3_cry_8_cZ(.DI(r0[8:8]),.CI(v_r1_3_cry_7),.S(v_r1_3_axb_8),.LO(v_r1_3_cry_8));
  XORCY v_r1_3_s_7(.LI(v_r1_3_axb_7),.CI(v_r1_3_cry_6),.O(v_r1_3[7:7]));
  MUXCY_L v_r1_3_cry_7_cZ(.DI(r0[7:7]),.CI(v_r1_3_cry_6),.S(v_r1_3_axb_7),.LO(v_r1_3_cry_7));
  XORCY v_r1_3_s_6(.LI(v_r1_3_axb_6),.CI(v_r1_3_cry_5),.O(v_r1_3[6:6]));
  MUXCY_L v_r1_3_cry_6_cZ(.DI(r0[6:6]),.CI(v_r1_3_cry_5),.S(v_r1_3_axb_6),.LO(v_r1_3_cry_6));
  XORCY v_r1_3_s_5(.LI(v_r1_3_axb_5),.CI(v_r1_3_cry_4),.O(v_r1_3[5:5]));
  MUXCY_L v_r1_3_cry_5_cZ(.DI(r0[5:5]),.CI(v_r1_3_cry_4),.S(v_r1_3_axb_5),.LO(v_r1_3_cry_5));
  XORCY v_r1_3_s_4(.LI(v_r1_3_axb_4),.CI(v_r1_3_cry_3),.O(v_r1_3[4:4]));
  MUXCY_L v_r1_3_cry_4_cZ(.DI(r0[4:4]),.CI(v_r1_3_cry_3),.S(v_r1_3_axb_4),.LO(v_r1_3_cry_4));
  XORCY v_r1_3_s_3(.LI(v_r1_3_axb_3),.CI(v_r1_3_cry_2),.O(v_r1_3[3:3]));
  MUXCY_L v_r1_3_cry_3_cZ(.DI(r0[3:3]),.CI(v_r1_3_cry_2),.S(v_r1_3_axb_3),.LO(v_r1_3_cry_3));
  XORCY v_r1_3_s_2(.LI(v_r1_3_axb_2),.CI(v_r1_3_cry_1),.O(v_r1_3[2:2]));
  MUXCY_L v_r1_3_cry_2_cZ(.DI(r0[2:2]),.CI(v_r1_3_cry_1),.S(v_r1_3_axb_2),.LO(v_r1_3_cry_2));
  XORCY v_r1_3_s_1(.LI(v_r1_3_axb_1),.CI(v_r1_3_cry_0),.O(v_r1_3[1:1]));
  MUXCY_L v_r1_3_cry_1_cZ(.DI(r0[1:1]),.CI(v_r1_3_cry_0),.S(v_r1_3_axb_1),.LO(v_r1_3_cry_1));
  XORCY v_r1_3_s_0(.LI(v_r1_3_axb_0),.CI(un14_s_state_cry[50:50]),.O(v_r1_3[0:0]));
  MUXCY_L v_r1_3_cry_0_cZ(.DI(r0[0:0]),.CI(un14_s_state_cry[50:50]),.S(v_r1_3_axb_0),.LO(v_r1_3_cry_0));
  XORCY un33_s_count_a_5_0_s_51(.LI(un33_s_count_a_5_0_axb_51),.CI(un33_s_count_a_5_0_cry_50),.O(un33_s_count_51));
  XORCY un33_s_count_a_5_0_s_50(.LI(un33_s_count_a_5_0_axb_50),.CI(un33_s_count_a_5_0_cry_49),.O(un33_s_count_50));
  MUXCY_L un33_s_count_a_5_0_cry_50_cZ(.DI(un33_s_count_a_5_0_cry_50_RNO),.CI(un33_s_count_a_5_0_cry_49),.S(un33_s_count_a_5_0_axb_50),.LO(un33_s_count_a_5_0_cry_50));
  XORCY un33_s_count_a_5_0_s_49(.LI(un33_s_count_a_5_0_axb_49),.CI(un33_s_count_a_5_0_cry_48),.O(un33_s_count_49));
  MUXCY_L un33_s_count_a_5_0_cry_49_cZ(.DI(un33_s_count_a_5_0_cry_49_RNO),.CI(un33_s_count_a_5_0_cry_48),.S(un33_s_count_a_5_0_axb_49),.LO(un33_s_count_a_5_0_cry_49));
  XORCY un33_s_count_a_5_0_s_48(.LI(un33_s_count_a_5_0_axb_48),.CI(un33_s_count_a_5_0_cry_47),.O(un33_s_count_48));
  MUXCY_L un33_s_count_a_5_0_cry_48_cZ(.DI(un33_s_count_a_5_0_cry_48_RNO),.CI(un33_s_count_a_5_0_cry_47),.S(un33_s_count_a_5_0_axb_48),.LO(un33_s_count_a_5_0_cry_48));
  XORCY un33_s_count_a_5_0_s_47(.LI(un33_s_count_a_5_0_axb_47),.CI(un33_s_count_a_5_0_cry_46),.O(un33_s_count_47));
  MUXCY_L un33_s_count_a_5_0_cry_47_cZ(.DI(un33_s_count_a_5_0_cry_47_RNO),.CI(un33_s_count_a_5_0_cry_46),.S(un33_s_count_a_5_0_axb_47),.LO(un33_s_count_a_5_0_cry_47));
  XORCY un33_s_count_a_5_0_s_46(.LI(un33_s_count_a_5_0_axb_46),.CI(un33_s_count_a_5_0_cry_45),.O(un33_s_count_46));
  MUXCY_L un33_s_count_a_5_0_cry_46_cZ(.DI(un33_s_count_a_5_0_cry_46_RNO),.CI(un33_s_count_a_5_0_cry_45),.S(un33_s_count_a_5_0_axb_46),.LO(un33_s_count_a_5_0_cry_46));
  XORCY un33_s_count_a_5_0_s_45(.LI(un33_s_count_a_5_0_axb_45),.CI(un33_s_count_a_5_0_cry_44),.O(un33_s_count_45));
  MUXCY_L un33_s_count_a_5_0_cry_45_cZ(.DI(un33_s_count_a_5_0_cry_45_RNO),.CI(un33_s_count_a_5_0_cry_44),.S(un33_s_count_a_5_0_axb_45),.LO(un33_s_count_a_5_0_cry_45));
  XORCY un33_s_count_a_5_0_s_44(.LI(un33_s_count_a_5_0_axb_44),.CI(un33_s_count_a_5_0_cry_43),.O(un33_s_count_44));
  MUXCY_L un33_s_count_a_5_0_cry_44_cZ(.DI(un33_s_count_a_5_0_cry_44_RNO),.CI(un33_s_count_a_5_0_cry_43),.S(un33_s_count_a_5_0_axb_44),.LO(un33_s_count_a_5_0_cry_44));
  XORCY un33_s_count_a_5_0_s_43(.LI(un33_s_count_a_5_0_axb_43),.CI(un33_s_count_a_5_0_cry_42),.O(un33_s_count_43));
  MUXCY_L un33_s_count_a_5_0_cry_43_cZ(.DI(un33_s_count_a_5_0_cry_43_RNO),.CI(un33_s_count_a_5_0_cry_42),.S(un33_s_count_a_5_0_axb_43),.LO(un33_s_count_a_5_0_cry_43));
  XORCY un33_s_count_a_5_0_s_42(.LI(un33_s_count_a_5_0_axb_42),.CI(un33_s_count_a_5_0_cry_41),.O(un33_s_count_42));
  MUXCY_L un33_s_count_a_5_0_cry_42_cZ(.DI(un33_s_count_a_5_0_cry_42_RNO),.CI(un33_s_count_a_5_0_cry_41),.S(un33_s_count_a_5_0_axb_42),.LO(un33_s_count_a_5_0_cry_42));
  XORCY un33_s_count_a_5_0_s_41(.LI(un33_s_count_a_5_0_axb_41),.CI(un33_s_count_a_5_0_cry_40),.O(un33_s_count_41));
  MUXCY_L un33_s_count_a_5_0_cry_41_cZ(.DI(un33_s_count_a_5_0_cry_41_RNO),.CI(un33_s_count_a_5_0_cry_40),.S(un33_s_count_a_5_0_axb_41),.LO(un33_s_count_a_5_0_cry_41));
  XORCY un33_s_count_a_5_0_s_40(.LI(un33_s_count_a_5_0_axb_40),.CI(un33_s_count_a_5_0_cry_39),.O(un33_s_count_40));
  MUXCY_L un33_s_count_a_5_0_cry_40_cZ(.DI(un33_s_count_a_5_0_cry_40_RNO),.CI(un33_s_count_a_5_0_cry_39),.S(un33_s_count_a_5_0_axb_40),.LO(un33_s_count_a_5_0_cry_40));
  XORCY un33_s_count_a_5_0_s_39(.LI(un33_s_count_a_5_0_axb_39),.CI(un33_s_count_a_5_0_cry_38),.O(un33_s_count_39));
  MUXCY_L un33_s_count_a_5_0_cry_39_cZ(.DI(un33_s_count_a_5_0_cry_39_RNO),.CI(un33_s_count_a_5_0_cry_38),.S(un33_s_count_a_5_0_axb_39),.LO(un33_s_count_a_5_0_cry_39));
  XORCY un33_s_count_a_5_0_s_38(.LI(un33_s_count_a_5_0_axb_38),.CI(un33_s_count_a_5_0_cry_37),.O(un33_s_count_38));
  MUXCY_L un33_s_count_a_5_0_cry_38_cZ(.DI(un33_s_count_a_5_0_cry_38_RNO),.CI(un33_s_count_a_5_0_cry_37),.S(un33_s_count_a_5_0_axb_38),.LO(un33_s_count_a_5_0_cry_38));
  XORCY un33_s_count_a_5_0_s_37(.LI(un33_s_count_a_5_0_axb_37),.CI(un33_s_count_a_5_0_cry_36),.O(un33_s_count_37));
  MUXCY_L un33_s_count_a_5_0_cry_37_cZ(.DI(un33_s_count_a_5_0_cry_37_RNO),.CI(un33_s_count_a_5_0_cry_36),.S(un33_s_count_a_5_0_axb_37),.LO(un33_s_count_a_5_0_cry_37));
  XORCY un33_s_count_a_5_0_s_36(.LI(un33_s_count_a_5_0_axb_36),.CI(un33_s_count_a_5_0_cry_35),.O(un33_s_count_36));
  MUXCY_L un33_s_count_a_5_0_cry_36_cZ(.DI(un33_s_count_a_5_0_cry_36_RNO),.CI(un33_s_count_a_5_0_cry_35),.S(un33_s_count_a_5_0_axb_36),.LO(un33_s_count_a_5_0_cry_36));
  XORCY un33_s_count_a_5_0_s_35(.LI(un33_s_count_a_5_0_axb_35),.CI(un33_s_count_a_5_0_cry_34),.O(un33_s_count_35));
  MUXCY_L un33_s_count_a_5_0_cry_35_cZ(.DI(un33_s_count_a_5_0_cry_35_RNO),.CI(un33_s_count_a_5_0_cry_34),.S(un33_s_count_a_5_0_axb_35),.LO(un33_s_count_a_5_0_cry_35));
  XORCY un33_s_count_a_5_0_s_34(.LI(un33_s_count_a_5_0_axb_34),.CI(un33_s_count_a_5_0_cry_33),.O(un33_s_count_34));
  MUXCY_L un33_s_count_a_5_0_cry_34_cZ(.DI(un33_s_count_a_5_0_cry_34_RNO),.CI(un33_s_count_a_5_0_cry_33),.S(un33_s_count_a_5_0_axb_34),.LO(un33_s_count_a_5_0_cry_34));
  XORCY un33_s_count_a_5_0_s_33(.LI(un33_s_count_a_5_0_axb_33),.CI(un33_s_count_a_5_0_cry_32),.O(un33_s_count_33));
  MUXCY_L un33_s_count_a_5_0_cry_33_cZ(.DI(un33_s_count_a_5_0_cry_33_RNO),.CI(un33_s_count_a_5_0_cry_32),.S(un33_s_count_a_5_0_axb_33),.LO(un33_s_count_a_5_0_cry_33));
  XORCY un33_s_count_a_5_0_s_32(.LI(un33_s_count_a_5_0_axb_32),.CI(un33_s_count_a_5_0_cry_31),.O(un33_s_count_32));
  MUXCY_L un33_s_count_a_5_0_cry_32_cZ(.DI(un33_s_count_a_5_0_cry_32_RNO),.CI(un33_s_count_a_5_0_cry_31),.S(un33_s_count_a_5_0_axb_32),.LO(un33_s_count_a_5_0_cry_32));
  XORCY un33_s_count_a_5_0_s_31(.LI(un33_s_count_a_5_0_axb_31),.CI(un33_s_count_a_5_0_cry_30),.O(un33_s_count_31));
  MUXCY_L un33_s_count_a_5_0_cry_31_cZ(.DI(un33_s_count_a_5_0_cry_31_RNO),.CI(un33_s_count_a_5_0_cry_30),.S(un33_s_count_a_5_0_axb_31),.LO(un33_s_count_a_5_0_cry_31));
  XORCY un33_s_count_a_5_0_s_30(.LI(un33_s_count_a_5_0_axb_30),.CI(un33_s_count_a_5_0_cry_29),.O(un33_s_count_30));
  MUXCY_L un33_s_count_a_5_0_cry_30_cZ(.DI(un33_s_count_a_5_0_cry_30_RNO),.CI(un33_s_count_a_5_0_cry_29),.S(un33_s_count_a_5_0_axb_30),.LO(un33_s_count_a_5_0_cry_30));
  XORCY un33_s_count_a_5_0_s_29(.LI(un33_s_count_a_5_0_axb_29),.CI(un33_s_count_a_5_0_cry_28),.O(un33_s_count_29));
  MUXCY_L un33_s_count_a_5_0_cry_29_cZ(.DI(un33_s_count_a_5_0_cry_29_RNO),.CI(un33_s_count_a_5_0_cry_28),.S(un33_s_count_a_5_0_axb_29),.LO(un33_s_count_a_5_0_cry_29));
  XORCY un33_s_count_a_5_0_s_28(.LI(un33_s_count_a_5_0_axb_28),.CI(un33_s_count_a_5_0_cry_27),.O(un33_s_count_28));
  MUXCY_L un33_s_count_a_5_0_cry_28_cZ(.DI(un33_s_count_a_5_0_cry_28_RNO),.CI(un33_s_count_a_5_0_cry_27),.S(un33_s_count_a_5_0_axb_28),.LO(un33_s_count_a_5_0_cry_28));
  XORCY un33_s_count_a_5_0_s_27(.LI(un33_s_count_a_5_0_axb_27),.CI(un33_s_count_a_5_0_cry_26),.O(un33_s_count_27));
  MUXCY_L un33_s_count_a_5_0_cry_27_cZ(.DI(r1_RNIABVR_O5[25:25]),.CI(un33_s_count_a_5_0_cry_26),.S(un33_s_count_a_5_0_axb_27),.LO(un33_s_count_a_5_0_cry_27));
  XORCY un33_s_count_a_5_0_s_26(.LI(un33_s_count_a_5_0_axb_26),.CI(un33_s_count_a_5_0_cry_25),.O(un33_s_count_a_5[26:26]));
  MUXCY_L un33_s_count_a_5_0_cry_26_cZ(.DI(un33_s_count_a_5_0_cry_26_RNO),.CI(un33_s_count_a_5_0_cry_25),.S(un33_s_count_a_5_0_axb_26),.LO(un33_s_count_a_5_0_cry_26));
  XORCY un33_s_count_a_5_0_s_25(.LI(un33_s_count_a_5_0_axb_25),.CI(un33_s_count_a_5_0_cry_24),.O(un33_s_count_a_5[25:25]));
  MUXCY_L un33_s_count_a_5_0_cry_25_cZ(.DI(un33_s_count_a_5_0_o5_24),.CI(un33_s_count_a_5_0_cry_24),.S(un33_s_count_a_5_0_axb_25),.LO(un33_s_count_a_5_0_cry_25));
  XORCY un33_s_count_a_5_0_s_24(.LI(un33_s_count_a_5_0_axb_24),.CI(un33_s_count_a_5_0_cry_23),.O(un33_s_count_a_5[24:24]));
  MUXCY_L un33_s_count_a_5_0_cry_24_cZ(.DI(un33_s_count_a_5_0_o5_23),.CI(un33_s_count_a_5_0_cry_23),.S(un33_s_count_a_5_0_axb_24),.LO(un33_s_count_a_5_0_cry_24));
  XORCY un33_s_count_a_5_0_s_23(.LI(un33_s_count_a_5_0_axb_23),.CI(un33_s_count_a_5_0_cry_22),.O(un33_s_count_a_5[23:23]));
  MUXCY_L un33_s_count_a_5_0_cry_23_cZ(.DI(un33_s_count_a_5_0_o5_22),.CI(un33_s_count_a_5_0_cry_22),.S(un33_s_count_a_5_0_axb_23),.LO(un33_s_count_a_5_0_cry_23));
  XORCY un33_s_count_a_5_0_s_22(.LI(un33_s_count_a_5_0_axb_22),.CI(un33_s_count_a_5_0_cry_21),.O(un33_s_count_a_5[22:22]));
  MUXCY_L un33_s_count_a_5_0_cry_22_cZ(.DI(un33_s_count_a_5_0_o5_21),.CI(un33_s_count_a_5_0_cry_21),.S(un33_s_count_a_5_0_axb_22),.LO(un33_s_count_a_5_0_cry_22));
  XORCY un33_s_count_a_5_0_s_21(.LI(un33_s_count_a_5_0_axb_21),.CI(un33_s_count_a_5_0_cry_20),.O(un33_s_count_a_5[21:21]));
  MUXCY_L un33_s_count_a_5_0_cry_21_cZ(.DI(un33_s_count_a_5_0_o5_20),.CI(un33_s_count_a_5_0_cry_20),.S(un33_s_count_a_5_0_axb_21),.LO(un33_s_count_a_5_0_cry_21));
  XORCY un33_s_count_a_5_0_s_20(.LI(un33_s_count_a_5_0_axb_20),.CI(un33_s_count_a_5_0_cry_19),.O(un33_s_count_a_5[20:20]));
  MUXCY_L un33_s_count_a_5_0_cry_20_cZ(.DI(un33_s_count_a_5_0_o5_19),.CI(un33_s_count_a_5_0_cry_19),.S(un33_s_count_a_5_0_axb_20),.LO(un33_s_count_a_5_0_cry_20));
  XORCY un33_s_count_a_5_0_s_19(.LI(un33_s_count_a_5_0_axb_19),.CI(un33_s_count_a_5_0_cry_18),.O(un33_s_count_a_5[19:19]));
  MUXCY_L un33_s_count_a_5_0_cry_19_cZ(.DI(un33_s_count_a_5_0_o5_18),.CI(un33_s_count_a_5_0_cry_18),.S(un33_s_count_a_5_0_axb_19),.LO(un33_s_count_a_5_0_cry_19));
  XORCY un33_s_count_a_5_0_s_18(.LI(un33_s_count_a_5_0_axb_18),.CI(un33_s_count_a_5_0_cry_17),.O(un33_s_count_a_5[18:18]));
  MUXCY_L un33_s_count_a_5_0_cry_18_cZ(.DI(un33_s_count_a_5_0_o5_17),.CI(un33_s_count_a_5_0_cry_17),.S(un33_s_count_a_5_0_axb_18),.LO(un33_s_count_a_5_0_cry_18));
  XORCY un33_s_count_a_5_0_s_17(.LI(un33_s_count_a_5_0_axb_17),.CI(un33_s_count_a_5_0_cry_16),.O(un33_s_count_a_5[17:17]));
  MUXCY_L un33_s_count_a_5_0_cry_17_cZ(.DI(un33_s_count_a_5_0_o5_16),.CI(un33_s_count_a_5_0_cry_16),.S(un33_s_count_a_5_0_axb_17),.LO(un33_s_count_a_5_0_cry_17));
  XORCY un33_s_count_a_5_0_s_16(.LI(un33_s_count_a_5_0_axb_16),.CI(un33_s_count_a_5_0_cry_15),.O(un33_s_count_a_5[16:16]));
  MUXCY_L un33_s_count_a_5_0_cry_16_cZ(.DI(un33_s_count_a_5_0_o5_15),.CI(un33_s_count_a_5_0_cry_15),.S(un33_s_count_a_5_0_axb_16),.LO(un33_s_count_a_5_0_cry_16));
  XORCY un33_s_count_a_5_0_s_15(.LI(un33_s_count_a_5_0_axb_15),.CI(un33_s_count_a_5_0_cry_14),.O(un33_s_count_a_5[15:15]));
  MUXCY_L un33_s_count_a_5_0_cry_15_cZ(.DI(un33_s_count_a_5_0_o5_14),.CI(un33_s_count_a_5_0_cry_14),.S(un33_s_count_a_5_0_axb_15),.LO(un33_s_count_a_5_0_cry_15));
  XORCY un33_s_count_a_5_0_s_14(.LI(un33_s_count_a_5_0_axb_14),.CI(un33_s_count_a_5_0_cry_13),.O(un33_s_count_a_5[14:14]));
  MUXCY_L un33_s_count_a_5_0_cry_14_cZ(.DI(un33_s_count_a_5_0_o5_13),.CI(un33_s_count_a_5_0_cry_13),.S(un33_s_count_a_5_0_axb_14),.LO(un33_s_count_a_5_0_cry_14));
  XORCY un33_s_count_a_5_0_s_13(.LI(un33_s_count_a_5_0_axb_13),.CI(un33_s_count_a_5_0_cry_12),.O(un33_s_count_a_5[13:13]));
  MUXCY_L un33_s_count_a_5_0_cry_13_cZ(.DI(un33_s_count_a_5_0_o5_12),.CI(un33_s_count_a_5_0_cry_12),.S(un33_s_count_a_5_0_axb_13),.LO(un33_s_count_a_5_0_cry_13));
  XORCY un33_s_count_a_5_0_s_12(.LI(un33_s_count_a_5_0_axb_12),.CI(un33_s_count_a_5_0_cry_11),.O(un33_s_count_a_5[12:12]));
  MUXCY_L un33_s_count_a_5_0_cry_12_cZ(.DI(un33_s_count_a_5_0_o5_11),.CI(un33_s_count_a_5_0_cry_11),.S(un33_s_count_a_5_0_axb_12),.LO(un33_s_count_a_5_0_cry_12));
  XORCY un33_s_count_a_5_0_s_11(.LI(un33_s_count_a_5_0_axb_11),.CI(un33_s_count_a_5_0_cry_10),.O(un33_s_count_a_5[11:11]));
  MUXCY_L un33_s_count_a_5_0_cry_11_cZ(.DI(un33_s_count_a_5_0_o5_10),.CI(un33_s_count_a_5_0_cry_10),.S(un33_s_count_a_5_0_axb_11),.LO(un33_s_count_a_5_0_cry_11));
  XORCY un33_s_count_a_5_0_s_10(.LI(un33_s_count_a_5_0_axb_10),.CI(un33_s_count_a_5_0_cry_9),.O(un33_s_count_a_5[10:10]));
  MUXCY_L un33_s_count_a_5_0_cry_10_cZ(.DI(un33_s_count_a_5_0_o5_9),.CI(un33_s_count_a_5_0_cry_9),.S(un33_s_count_a_5_0_axb_10),.LO(un33_s_count_a_5_0_cry_10));
  XORCY un33_s_count_a_5_0_s_9(.LI(un33_s_count_a_5_0_axb_9),.CI(un33_s_count_a_5_0_cry_8),.O(un33_s_count_a_5[9:9]));
  MUXCY_L un33_s_count_a_5_0_cry_9_cZ(.DI(un33_s_count_a_5_0_o5_8),.CI(un33_s_count_a_5_0_cry_8),.S(un33_s_count_a_5_0_axb_9),.LO(un33_s_count_a_5_0_cry_9));
  XORCY un33_s_count_a_5_0_s_8(.LI(un33_s_count_a_5_0_axb_8),.CI(un33_s_count_a_5_0_cry_7),.O(un33_s_count_a_5[8:8]));
  MUXCY_L un33_s_count_a_5_0_cry_8_cZ(.DI(un33_s_count_a_5_0_o5_7),.CI(un33_s_count_a_5_0_cry_7),.S(un33_s_count_a_5_0_axb_8),.LO(un33_s_count_a_5_0_cry_8));
  XORCY un33_s_count_a_5_0_s_7(.LI(un33_s_count_a_5_0_axb_7),.CI(un33_s_count_a_5_0_cry_6),.O(un33_s_count_a_5[7:7]));
  MUXCY_L un33_s_count_a_5_0_cry_7_cZ(.DI(un33_s_count_a_5_0_o5_6),.CI(un33_s_count_a_5_0_cry_6),.S(un33_s_count_a_5_0_axb_7),.LO(un33_s_count_a_5_0_cry_7));
  XORCY un33_s_count_a_5_0_s_6(.LI(un33_s_count_a_5_0_axb_6),.CI(un33_s_count_a_5_0_cry_5),.O(un33_s_count_a_5[6:6]));
  MUXCY_L un33_s_count_a_5_0_cry_6_cZ(.DI(un33_s_count_a_5_0_o5_5),.CI(un33_s_count_a_5_0_cry_5),.S(un33_s_count_a_5_0_axb_6),.LO(un33_s_count_a_5_0_cry_6));
  XORCY un33_s_count_a_5_0_s_5(.LI(un33_s_count_a_5_0_axb_5),.CI(un33_s_count_a_5_0_cry_4),.O(un33_s_count_a_5[5:5]));
  MUXCY_L un33_s_count_a_5_0_cry_5_cZ(.DI(un33_s_count_a_5_0_o5_4),.CI(un33_s_count_a_5_0_cry_4),.S(un33_s_count_a_5_0_axb_5),.LO(un33_s_count_a_5_0_cry_5));
  XORCY un33_s_count_a_5_0_s_4(.LI(un33_s_count_a_5_0_axb_4),.CI(un33_s_count_a_5_0_cry_3),.O(un33_s_count_a_5[4:4]));
  MUXCY_L un33_s_count_a_5_0_cry_4_cZ(.DI(un33_s_count_a_5_0_o5_3),.CI(un33_s_count_a_5_0_cry_3),.S(un33_s_count_a_5_0_axb_4),.LO(un33_s_count_a_5_0_cry_4));
  XORCY un33_s_count_a_5_0_s_3(.LI(un33_s_count_a_5_0_axb_3),.CI(un33_s_count_a_5_0_cry_2),.O(un33_s_count_a_5[3:3]));
  MUXCY_L un33_s_count_a_5_0_cry_3_cZ(.DI(un33_s_count_a_5_0_axb_2_lut6_2_O5),.CI(un33_s_count_a_5_0_cry_2),.S(un33_s_count_a_5_0_axb_3),.LO(un33_s_count_a_5_0_cry_3));
  XORCY un33_s_count_a_5_0_s_2(.LI(un33_s_count_a_5_0_axb_2),.CI(un33_s_count_a_5_0_cry_1),.O(un33_s_count_a_5[2:2]));
  MUXCY_L un33_s_count_a_5_0_cry_2_cZ(.DI(r1_2[1:1]),.CI(un33_s_count_a_5_0_cry_1),.S(un33_s_count_a_5_0_axb_2),.LO(un33_s_count_a_5_0_cry_2));
  XORCY un33_s_count_a_5_0_s_1(.LI(un33_s_count_a_5_0_axb_1),.CI(un33_s_count_a_5_0_cry_0),.O(un33_s_count_1));
  MUXCY_L un33_s_count_a_5_0_cry_1_cZ(.DI(r1_2_i[1:1]),.CI(un33_s_count_a_5_0_cry_0),.S(un33_s_count_a_5_0_axb_1),.LO(un33_s_count_a_5_0_cry_1));
  MUXCY_L un33_s_count_a_5_0_cry_0_cZ(.DI(VCC),.CI(GND),.S(r1_2_i[0:0]),.LO(un33_s_count_a_5_0_cry_0));
  XORCY v_r1_2_3_0_s_51(.LI(v_r1_2_3_0_axb_51),.CI(v_r1_2_3_0_cry_50),.O(v_r1_2_3[51:51]));
  XORCY v_r1_2_3_0_s_50(.LI(v_r1_2_3_0_axb_50),.CI(v_r1_2_3_0_cry_49),.O(v_r1_2_3[50:50]));
  MUXCY_L v_r1_2_3_0_cry_50_cZ(.DI(v_r1_2_3_0_cry_50_RNO),.CI(v_r1_2_3_0_cry_49),.S(v_r1_2_3_0_axb_50),.LO(v_r1_2_3_0_cry_50));
  XORCY v_r1_2_3_0_s_49(.LI(v_r1_2_3_0_axb_49),.CI(v_r1_2_3_0_cry_48),.O(v_r1_2_3[49:49]));
  MUXCY_L v_r1_2_3_0_cry_49_cZ(.DI(v_r1_2_3_0_cry_49_RNO),.CI(v_r1_2_3_0_cry_48),.S(v_r1_2_3_0_axb_49),.LO(v_r1_2_3_0_cry_49));
  XORCY v_r1_2_3_0_s_48(.LI(v_r1_2_3_0_axb_48),.CI(v_r1_2_3_0_cry_47),.O(v_r1_2_3[48:48]));
  MUXCY_L v_r1_2_3_0_cry_48_cZ(.DI(v_r1_2_3_0_cry_48_RNO),.CI(v_r1_2_3_0_cry_47),.S(v_r1_2_3_0_axb_48),.LO(v_r1_2_3_0_cry_48));
  XORCY v_r1_2_3_0_s_47(.LI(v_r1_2_3_0_axb_47),.CI(v_r1_2_3_0_cry_46),.O(v_r1_2_3[47:47]));
  MUXCY_L v_r1_2_3_0_cry_47_cZ(.DI(v_r1_2_3_0_cry_47_RNO),.CI(v_r1_2_3_0_cry_46),.S(v_r1_2_3_0_axb_47),.LO(v_r1_2_3_0_cry_47));
  XORCY v_r1_2_3_0_s_46(.LI(v_r1_2_3_0_axb_46),.CI(v_r1_2_3_0_cry_45),.O(v_r1_2_3[46:46]));
  MUXCY_L v_r1_2_3_0_cry_46_cZ(.DI(v_r1_2_3_0_cry_46_RNO),.CI(v_r1_2_3_0_cry_45),.S(v_r1_2_3_0_axb_46),.LO(v_r1_2_3_0_cry_46));
  XORCY v_r1_2_3_0_s_45(.LI(v_r1_2_3_0_axb_45),.CI(v_r1_2_3_0_cry_44),.O(v_r1_2_3[45:45]));
  MUXCY_L v_r1_2_3_0_cry_45_cZ(.DI(v_r1_2_3_0_cry_45_RNO),.CI(v_r1_2_3_0_cry_44),.S(v_r1_2_3_0_axb_45),.LO(v_r1_2_3_0_cry_45));
  XORCY v_r1_2_3_0_s_44(.LI(v_r1_2_3_0_axb_44),.CI(v_r1_2_3_0_cry_43),.O(v_r1_2_3[44:44]));
  MUXCY_L v_r1_2_3_0_cry_44_cZ(.DI(v_r1_2_3_0_cry_44_RNO),.CI(v_r1_2_3_0_cry_43),.S(v_r1_2_3_0_axb_44),.LO(v_r1_2_3_0_cry_44));
  XORCY v_r1_2_3_0_s_43(.LI(v_r1_2_3_0_axb_43),.CI(v_r1_2_3_0_cry_42),.O(v_r1_2_3[43:43]));
  MUXCY_L v_r1_2_3_0_cry_43_cZ(.DI(v_r1_2_3_0_cry_43_RNO),.CI(v_r1_2_3_0_cry_42),.S(v_r1_2_3_0_axb_43),.LO(v_r1_2_3_0_cry_43));
  XORCY v_r1_2_3_0_s_42(.LI(v_r1_2_3_0_axb_42),.CI(v_r1_2_3_0_cry_41),.O(v_r1_2_3[42:42]));
  MUXCY_L v_r1_2_3_0_cry_42_cZ(.DI(v_r1_2_3_0_cry_42_RNO),.CI(v_r1_2_3_0_cry_41),.S(v_r1_2_3_0_axb_42),.LO(v_r1_2_3_0_cry_42));
  XORCY v_r1_2_3_0_s_41(.LI(v_r1_2_3_0_axb_41),.CI(v_r1_2_3_0_cry_40),.O(v_r1_2_3[41:41]));
  MUXCY_L v_r1_2_3_0_cry_41_cZ(.DI(v_r1_2_3_0_cry_41_RNO),.CI(v_r1_2_3_0_cry_40),.S(v_r1_2_3_0_axb_41),.LO(v_r1_2_3_0_cry_41));
  XORCY v_r1_2_3_0_s_40(.LI(v_r1_2_3_0_axb_40),.CI(v_r1_2_3_0_cry_39),.O(v_r1_2_3[40:40]));
  MUXCY_L v_r1_2_3_0_cry_40_cZ(.DI(v_r1_2_3_0_cry_40_RNO),.CI(v_r1_2_3_0_cry_39),.S(v_r1_2_3_0_axb_40),.LO(v_r1_2_3_0_cry_40));
  XORCY v_r1_2_3_0_s_39(.LI(v_r1_2_3_0_axb_39),.CI(v_r1_2_3_0_cry_38),.O(v_r1_2_3[39:39]));
  MUXCY_L v_r1_2_3_0_cry_39_cZ(.DI(v_r1_2_3_0_cry_39_RNO),.CI(v_r1_2_3_0_cry_38),.S(v_r1_2_3_0_axb_39),.LO(v_r1_2_3_0_cry_39));
  XORCY v_r1_2_3_0_s_38(.LI(v_r1_2_3_0_axb_38),.CI(v_r1_2_3_0_cry_37),.O(v_r1_2_3[38:38]));
  MUXCY_L v_r1_2_3_0_cry_38_cZ(.DI(v_r1_2_3_0_cry_38_RNO),.CI(v_r1_2_3_0_cry_37),.S(v_r1_2_3_0_axb_38),.LO(v_r1_2_3_0_cry_38));
  XORCY v_r1_2_3_0_s_37(.LI(v_r1_2_3_0_axb_37),.CI(v_r1_2_3_0_cry_36),.O(v_r1_2_3[37:37]));
  MUXCY_L v_r1_2_3_0_cry_37_cZ(.DI(v_r1_2_3_0_cry_37_RNO),.CI(v_r1_2_3_0_cry_36),.S(v_r1_2_3_0_axb_37),.LO(v_r1_2_3_0_cry_37));
  XORCY v_r1_2_3_0_s_36(.LI(v_r1_2_3_0_axb_36),.CI(v_r1_2_3_0_cry_35),.O(v_r1_2_3[36:36]));
  MUXCY_L v_r1_2_3_0_cry_36_cZ(.DI(v_r1_2_3_0_cry_36_RNO),.CI(v_r1_2_3_0_cry_35),.S(v_r1_2_3_0_axb_36),.LO(v_r1_2_3_0_cry_36));
  XORCY v_r1_2_3_0_s_35(.LI(v_r1_2_3_0_axb_35),.CI(v_r1_2_3_0_cry_34),.O(v_r1_2_3[35:35]));
  MUXCY_L v_r1_2_3_0_cry_35_cZ(.DI(v_r1_2_3_0_cry_35_RNO),.CI(v_r1_2_3_0_cry_34),.S(v_r1_2_3_0_axb_35),.LO(v_r1_2_3_0_cry_35));
  XORCY v_r1_2_3_0_s_34(.LI(v_r1_2_3_0_axb_34),.CI(v_r1_2_3_0_cry_33),.O(v_r1_2_3[34:34]));
  MUXCY_L v_r1_2_3_0_cry_34_cZ(.DI(v_r1_2_3_0_cry_34_RNO),.CI(v_r1_2_3_0_cry_33),.S(v_r1_2_3_0_axb_34),.LO(v_r1_2_3_0_cry_34));
  XORCY v_r1_2_3_0_s_33(.LI(v_r1_2_3_0_axb_33),.CI(v_r1_2_3_0_cry_32),.O(v_r1_2_3[33:33]));
  MUXCY_L v_r1_2_3_0_cry_33_cZ(.DI(v_r1_2_3_0_cry_33_RNO),.CI(v_r1_2_3_0_cry_32),.S(v_r1_2_3_0_axb_33),.LO(v_r1_2_3_0_cry_33));
  XORCY v_r1_2_3_0_s_32(.LI(v_r1_2_3_0_axb_32),.CI(v_r1_2_3_0_cry_31),.O(v_r1_2_3[32:32]));
  MUXCY_L v_r1_2_3_0_cry_32_cZ(.DI(v_r1_2_3_0_cry_32_RNO),.CI(v_r1_2_3_0_cry_31),.S(v_r1_2_3_0_axb_32),.LO(v_r1_2_3_0_cry_32));
  XORCY v_r1_2_3_0_s_31(.LI(v_r1_2_3_0_axb_31),.CI(v_r1_2_3_0_cry_30),.O(v_r1_2_3[31:31]));
  MUXCY_L v_r1_2_3_0_cry_31_cZ(.DI(v_r1_2_3_0_cry_31_RNO),.CI(v_r1_2_3_0_cry_30),.S(v_r1_2_3_0_axb_31),.LO(v_r1_2_3_0_cry_31));
  XORCY v_r1_2_3_0_s_30(.LI(v_r1_2_3_0_axb_30),.CI(v_r1_2_3_0_cry_29),.O(v_r1_2_3[30:30]));
  MUXCY_L v_r1_2_3_0_cry_30_cZ(.DI(v_r1_2_3_0_cry_30_RNO),.CI(v_r1_2_3_0_cry_29),.S(v_r1_2_3_0_axb_30),.LO(v_r1_2_3_0_cry_30));
  XORCY v_r1_2_3_0_s_29(.LI(v_r1_2_3_0_axb_29),.CI(v_r1_2_3_0_cry_28),.O(v_r1_2_3[29:29]));
  MUXCY_L v_r1_2_3_0_cry_29_cZ(.DI(v_r1_2_3_0_cry_29_RNO),.CI(v_r1_2_3_0_cry_28),.S(v_r1_2_3_0_axb_29),.LO(v_r1_2_3_0_cry_29));
  XORCY v_r1_2_3_0_s_28(.LI(v_r1_2_3_0_axb_28),.CI(v_r1_2_3_0_cry_27),.O(v_r1_2_3[28:28]));
  MUXCY_L v_r1_2_3_0_cry_28_cZ(.DI(v_r1_2_3_0_cry_28_RNO),.CI(v_r1_2_3_0_cry_27),.S(v_r1_2_3_0_axb_28),.LO(v_r1_2_3_0_cry_28));
  XORCY v_r1_2_3_0_s_27(.LI(v_r1_2_3_0_axb_27),.CI(v_r1_2_3_0_cry_26),.O(v_r1_2_3[27:27]));
  MUXCY_L v_r1_2_3_0_cry_27_cZ(.DI(v_r1_2_3_0_o5_26),.CI(v_r1_2_3_0_cry_26),.S(v_r1_2_3_0_axb_27),.LO(v_r1_2_3_0_cry_27));
  XORCY v_r1_2_3_0_s_26(.LI(v_r1_2_3_0_axb_26),.CI(v_r1_2_3_0_cry_25),.O(v_r1_2_3[26:26]));
  MUXCY_L v_r1_2_3_0_cry_26_cZ(.DI(v_r1_2_3_0_cry_26_RNO),.CI(v_r1_2_3_0_cry_25),.S(v_r1_2_3_0_axb_26),.LO(v_r1_2_3_0_cry_26));
  XORCY v_r1_2_3_0_s_25(.LI(v_r1_2_3_0_axb_25),.CI(v_r1_2_3_0_cry_24),.O(v_r1_2_3[25:25]));
  MUXCY_L v_r1_2_3_0_cry_25_cZ(.DI(v_r1_2_3_0_o5_24),.CI(v_r1_2_3_0_cry_24),.S(v_r1_2_3_0_axb_25),.LO(v_r1_2_3_0_cry_25));
  XORCY v_r1_2_3_0_s_24(.LI(v_r1_2_3_0_axb_24),.CI(v_r1_2_3_0_cry_23),.O(v_r1_2_3[24:24]));
  MUXCY_L v_r1_2_3_0_cry_24_cZ(.DI(v_r1_2_3_0_cry_24_RNO),.CI(v_r1_2_3_0_cry_23),.S(v_r1_2_3_0_axb_24),.LO(v_r1_2_3_0_cry_24));
  XORCY v_r1_2_3_0_s_23(.LI(v_r1_2_3_0_axb_23),.CI(v_r1_2_3_0_cry_22),.O(v_r1_2_3[23:23]));
  MUXCY_L v_r1_2_3_0_cry_23_cZ(.DI(v_r1_2_3_0_cry_23_RNO),.CI(v_r1_2_3_0_cry_22),.S(v_r1_2_3_0_axb_23),.LO(v_r1_2_3_0_cry_23));
  XORCY v_r1_2_3_0_s_22(.LI(v_r1_2_3_0_axb_22),.CI(v_r1_2_3_0_cry_21),.O(v_r1_2_3[22:22]));
  MUXCY_L v_r1_2_3_0_cry_22_cZ(.DI(v_r1_2_3_0_cry_22_RNO),.CI(v_r1_2_3_0_cry_21),.S(v_r1_2_3_0_axb_22),.LO(v_r1_2_3_0_cry_22));
  XORCY v_r1_2_3_0_s_21(.LI(v_r1_2_3_0_axb_21),.CI(v_r1_2_3_0_cry_20),.O(v_r1_2_3[21:21]));
  MUXCY_L v_r1_2_3_0_cry_21_cZ(.DI(v_r1_2_3_0_cry_21_RNO),.CI(v_r1_2_3_0_cry_20),.S(v_r1_2_3_0_axb_21),.LO(v_r1_2_3_0_cry_21));
  XORCY v_r1_2_3_0_s_20(.LI(v_r1_2_3_0_axb_20),.CI(v_r1_2_3_0_cry_19),.O(v_r1_2_3[20:20]));
  MUXCY_L v_r1_2_3_0_cry_20_cZ(.DI(v_r1_2_3_0_cry_20_RNO),.CI(v_r1_2_3_0_cry_19),.S(v_r1_2_3_0_axb_20),.LO(v_r1_2_3_0_cry_20));
  XORCY v_r1_2_3_0_s_19(.LI(v_r1_2_3_0_axb_19),.CI(v_r1_2_3_0_cry_18),.O(v_r1_2_3[19:19]));
  MUXCY_L v_r1_2_3_0_cry_19_cZ(.DI(v_r1_2_3_0_cry_19_RNO),.CI(v_r1_2_3_0_cry_18),.S(v_r1_2_3_0_axb_19),.LO(v_r1_2_3_0_cry_19));
  XORCY v_r1_2_3_0_s_18(.LI(v_r1_2_3_0_axb_18),.CI(v_r1_2_3_0_cry_17),.O(v_r1_2_3[18:18]));
  MUXCY_L v_r1_2_3_0_cry_18_cZ(.DI(v_r1_2_3_0_cry_18_RNO),.CI(v_r1_2_3_0_cry_17),.S(v_r1_2_3_0_axb_18),.LO(v_r1_2_3_0_cry_18));
  XORCY v_r1_2_3_0_s_17(.LI(v_r1_2_3_0_axb_17),.CI(v_r1_2_3_0_cry_16),.O(v_r1_2_3[17:17]));
  MUXCY_L v_r1_2_3_0_cry_17_cZ(.DI(v_r1_2_3_0_cry_17_RNO),.CI(v_r1_2_3_0_cry_16),.S(v_r1_2_3_0_axb_17),.LO(v_r1_2_3_0_cry_17));
  XORCY v_r1_2_3_0_s_16(.LI(v_r1_2_3_0_axb_16),.CI(v_r1_2_3_0_cry_15),.O(v_r1_2_3[16:16]));
  MUXCY_L v_r1_2_3_0_cry_16_cZ(.DI(v_r1_2_3_0_cry_16_RNO),.CI(v_r1_2_3_0_cry_15),.S(v_r1_2_3_0_axb_16),.LO(v_r1_2_3_0_cry_16));
  XORCY v_r1_2_3_0_s_15(.LI(v_r1_2_3_0_axb_15),.CI(v_r1_2_3_0_cry_14),.O(v_r1_2_3[15:15]));
  MUXCY_L v_r1_2_3_0_cry_15_cZ(.DI(v_r1_2_3_0_cry_15_RNO),.CI(v_r1_2_3_0_cry_14),.S(v_r1_2_3_0_axb_15),.LO(v_r1_2_3_0_cry_15));
  XORCY v_r1_2_3_0_s_14(.LI(v_r1_2_3_0_axb_14),.CI(v_r1_2_3_0_cry_13),.O(v_r1_2_3[14:14]));
  MUXCY_L v_r1_2_3_0_cry_14_cZ(.DI(v_r1_2_3_0_cry_14_RNO),.CI(v_r1_2_3_0_cry_13),.S(v_r1_2_3_0_axb_14),.LO(v_r1_2_3_0_cry_14));
  XORCY v_r1_2_3_0_s_13(.LI(v_r1_2_3_0_axb_13),.CI(v_r1_2_3_0_cry_12),.O(v_r1_2_3[13:13]));
  MUXCY_L v_r1_2_3_0_cry_13_cZ(.DI(v_r1_2_3_0_cry_13_RNO),.CI(v_r1_2_3_0_cry_12),.S(v_r1_2_3_0_axb_13),.LO(v_r1_2_3_0_cry_13));
  XORCY v_r1_2_3_0_s_12(.LI(v_r1_2_3_0_axb_12),.CI(v_r1_2_3_0_cry_11),.O(v_r1_2_3[12:12]));
  MUXCY_L v_r1_2_3_0_cry_12_cZ(.DI(v_r1_2_3_0_cry_12_RNO),.CI(v_r1_2_3_0_cry_11),.S(v_r1_2_3_0_axb_12),.LO(v_r1_2_3_0_cry_12));
  XORCY v_r1_2_3_0_s_11(.LI(v_r1_2_3_0_axb_11),.CI(v_r1_2_3_0_cry_10),.O(v_r1_2_3[11:11]));
  MUXCY_L v_r1_2_3_0_cry_11_cZ(.DI(v_r1_2_3_0_cry_11_RNO),.CI(v_r1_2_3_0_cry_10),.S(v_r1_2_3_0_axb_11),.LO(v_r1_2_3_0_cry_11));
  XORCY v_r1_2_3_0_s_10(.LI(v_r1_2_3_0_axb_10),.CI(v_r1_2_3_0_cry_9),.O(v_r1_2_3[10:10]));
  MUXCY_L v_r1_2_3_0_cry_10_cZ(.DI(v_r1_2_3_0_cry_10_RNO),.CI(v_r1_2_3_0_cry_9),.S(v_r1_2_3_0_axb_10),.LO(v_r1_2_3_0_cry_10));
  XORCY v_r1_2_3_0_s_9(.LI(v_r1_2_3_0_axb_9),.CI(v_r1_2_3_0_cry_8),.O(v_r1_2_3[9:9]));
  MUXCY_L v_r1_2_3_0_cry_9_cZ(.DI(v_r1_2_3_0_cry_9_RNO),.CI(v_r1_2_3_0_cry_8),.S(v_r1_2_3_0_axb_9),.LO(v_r1_2_3_0_cry_9));
  XORCY v_r1_2_3_0_s_8(.LI(v_r1_2_3_0_axb_8),.CI(v_r1_2_3_0_cry_7),.O(v_r1_2_3[8:8]));
  MUXCY_L v_r1_2_3_0_cry_8_cZ(.DI(v_r1_2_3_0_cry_8_RNO),.CI(v_r1_2_3_0_cry_7),.S(v_r1_2_3_0_axb_8),.LO(v_r1_2_3_0_cry_8));
  XORCY v_r1_2_3_0_s_7(.LI(v_r1_2_3_0_axb_7),.CI(v_r1_2_3_0_cry_6),.O(v_r1_2_3[7:7]));
  MUXCY_L v_r1_2_3_0_cry_7_cZ(.DI(v_r1_2_3_0_cry_7_RNO),.CI(v_r1_2_3_0_cry_6),.S(v_r1_2_3_0_axb_7),.LO(v_r1_2_3_0_cry_7));
  XORCY v_r1_2_3_0_s_6(.LI(v_r1_2_3_0_axb_6),.CI(v_r1_2_3_0_cry_5),.O(v_r1_2_3[6:6]));
  MUXCY_L v_r1_2_3_0_cry_6_cZ(.DI(v_r1_2_3_0_cry_6_RNO),.CI(v_r1_2_3_0_cry_5),.S(v_r1_2_3_0_axb_6),.LO(v_r1_2_3_0_cry_6));
  XORCY v_r1_2_3_0_s_5(.LI(v_r1_2_3_0_axb_5),.CI(v_r1_2_3_0_cry_4),.O(v_r1_2_3[5:5]));
  MUXCY_L v_r1_2_3_0_cry_5_cZ(.DI(v_r1_2_3_0_cry_5_RNO),.CI(v_r1_2_3_0_cry_4),.S(v_r1_2_3_0_axb_5),.LO(v_r1_2_3_0_cry_5));
  XORCY v_r1_2_3_0_s_4(.LI(v_r1_2_3_0_axb_4),.CI(v_r1_2_3_0_cry_3),.O(v_r1_2_3[4:4]));
  MUXCY_L v_r1_2_3_0_cry_4_cZ(.DI(v_r1_2_3_0_cry_4_RNO),.CI(v_r1_2_3_0_cry_3),.S(v_r1_2_3_0_axb_4),.LO(v_r1_2_3_0_cry_4));
  XORCY v_r1_2_3_0_s_3(.LI(v_r1_2_3_0_axb_3),.CI(v_r1_2_3_0_cry_2),.O(v_r1_2_3[3:3]));
  MUXCY_L v_r1_2_3_0_cry_3_cZ(.DI(v_r1_2_3_0_cry_3_RNO),.CI(v_r1_2_3_0_cry_2),.S(v_r1_2_3_0_axb_3),.LO(v_r1_2_3_0_cry_3));
  XORCY v_r1_2_3_0_s_2(.LI(v_r1_2_3_0_axb_2),.CI(v_r1_2_3_0_cry_1),.O(v_r1_2_3[2:2]));
  MUXCY_L v_r1_2_3_0_cry_2_cZ(.DI(v_r1_2_3_0_cry_2_RNO),.CI(v_r1_2_3_0_cry_1),.S(v_r1_2_3_0_axb_2),.LO(v_r1_2_3_0_cry_2));
  XORCY v_r1_2_3_0_s_1(.LI(v_r1_2_3_0_axb_1),.CI(v_r1_2_3_0_cry_0),.O(v_r1_2_3[1:1]));
  MUXCY_L v_r1_2_3_0_cry_1_cZ(.DI(v_r1_2_3_0_cry_1_RNO),.CI(v_r1_2_3_0_cry_0),.S(v_r1_2_3_0_axb_1),.LO(v_r1_2_3_0_cry_1));
  XORCY v_r1_2_3_0_s_0(.LI(v_r1_2_3_0_axb_0),.CI(v_r1_2_3_0_cry_0_cy),.O(v_r1_2_3[0:0]));
  MUXCY_L v_r1_2_3_0_cry_0_cZ(.DI(un14_s_state_cry[50:50]),.CI(v_r1_2_3_0_cry_0_cy),.S(v_r1_2_3_0_axb_0),.LO(v_r1_2_3_0_cry_0));
  MUXCY_L desc3002(.DI(un27_s_count_lt48),.CI(un27_s_count_cry[46:46]),.S(un27_s_count_df48),.LO(un27_s_count_cry[48:48]));
  MUXCY_L desc3003(.DI(un27_s_count_lt46),.CI(un27_s_count_cry[44:44]),.S(un27_s_count_df46),.LO(un27_s_count_cry[46:46]));
  MUXCY_L desc3004(.DI(un27_s_count_lt44),.CI(un27_s_count_cry[42:42]),.S(un27_s_count_df44),.LO(un27_s_count_cry[44:44]));
  MUXCY_L desc3005(.DI(un27_s_count_lt42),.CI(un27_s_count_cry[40:40]),.S(un27_s_count_df42),.LO(un27_s_count_cry[42:42]));
  MUXCY_L desc3006(.DI(un27_s_count_lt40),.CI(un27_s_count_cry[38:38]),.S(un27_s_count_df40),.LO(un27_s_count_cry[40:40]));
  MUXCY_L desc3007(.DI(un27_s_count_lt38),.CI(un27_s_count_cry[36:36]),.S(un27_s_count_df38),.LO(un27_s_count_cry[38:38]));
  MUXCY_L desc3008(.DI(un27_s_count_lt36),.CI(un27_s_count_cry[34:34]),.S(un27_s_count_df36),.LO(un27_s_count_cry[36:36]));
  MUXCY_L desc3009(.DI(un27_s_count_lt34),.CI(un27_s_count_cry[32:32]),.S(un27_s_count_df34),.LO(un27_s_count_cry[34:34]));
  MUXCY_L desc3010(.DI(un27_s_count_lt32),.CI(un27_s_count_cry[30:30]),.S(un27_s_count_df32),.LO(un27_s_count_cry[32:32]));
  MUXCY_L desc3011(.DI(un27_s_count_lt30),.CI(un27_s_count_cry[28:28]),.S(un27_s_count_df30),.LO(un27_s_count_cry[30:30]));
  MUXCY_L desc3012(.DI(un27_s_count_lt28),.CI(un27_s_count_cry[26:26]),.S(un27_s_count_df28),.LO(un27_s_count_cry[28:28]));
  MUXCY_L desc3013(.DI(un27_s_count_lt26),.CI(un27_s_count_cry[24:24]),.S(un27_s_count_df26),.LO(un27_s_count_cry[26:26]));
  MUXCY_L desc3014(.DI(un27_s_count_lt24),.CI(un27_s_count_cry[22:22]),.S(un27_s_count_df24),.LO(un27_s_count_cry[24:24]));
  MUXCY_L desc3015(.DI(un27_s_count_lt22),.CI(un27_s_count_cry[20:20]),.S(un27_s_count_df22),.LO(un27_s_count_cry[22:22]));
  MUXCY_L desc3016(.DI(un27_s_count_lt20),.CI(un27_s_count_cry[18:18]),.S(un27_s_count_df20),.LO(un27_s_count_cry[20:20]));
  MUXCY_L desc3017(.DI(un27_s_count_lt18),.CI(un27_s_count_cry[16:16]),.S(un27_s_count_df18),.LO(un27_s_count_cry[18:18]));
  MUXCY_L desc3018(.DI(un27_s_count_lt16),.CI(un27_s_count_cry[14:14]),.S(un27_s_count_df16),.LO(un27_s_count_cry[16:16]));
  MUXCY_L desc3019(.DI(un27_s_count_lt14),.CI(un27_s_count_cry[12:12]),.S(un27_s_count_df14),.LO(un27_s_count_cry[14:14]));
  MUXCY_L desc3020(.DI(un27_s_count_lt12),.CI(un27_s_count_cry[10:10]),.S(un27_s_count_df12),.LO(un27_s_count_cry[12:12]));
  MUXCY_L desc3021(.DI(un27_s_count_lt10),.CI(un27_s_count_cry[8:8]),.S(un27_s_count_df10),.LO(un27_s_count_cry[10:10]));
  MUXCY_L desc3022(.DI(un27_s_count_lt8),.CI(un27_s_count_cry[6:6]),.S(un27_s_count_df8),.LO(un27_s_count_cry[8:8]));
  MUXCY_L desc3023(.DI(un27_s_count_lt6),.CI(un27_s_count_cry[4:4]),.S(un27_s_count_df6),.LO(un27_s_count_cry[6:6]));
  MUXCY_L desc3024(.DI(un27_s_count_lt4),.CI(un27_s_count_cry[2:2]),.S(un27_s_count_df4),.LO(un27_s_count_cry[4:4]));
  MUXCY_L desc3025(.DI(un27_s_count_lt2),.CI(un27_s_count_cry[0:0]),.S(un27_s_count_df2),.LO(un27_s_count_cry[2:2]));
  MUXCY_L desc3026(.DI(un27_s_count_lt0),.CI(GND),.S(un27_s_count_df0),.LO(un27_s_count_cry[0:0]));
  MUXCY_L desc3027(.DI(un14_s_state_lt48),.CI(un14_s_state_cry[46:46]),.S(un14_s_state_df48),.LO(un14_s_state_cry[48:48]));
  MUXCY_L desc3028(.DI(un14_s_state_lt46),.CI(un14_s_state_cry[44:44]),.S(un14_s_state_df46),.LO(un14_s_state_cry[46:46]));
  MUXCY_L desc3029(.DI(un14_s_state_lt44),.CI(un14_s_state_cry[42:42]),.S(un14_s_state_df44),.LO(un14_s_state_cry[44:44]));
  MUXCY_L desc3030(.DI(un14_s_state_lt42),.CI(un14_s_state_cry[40:40]),.S(un14_s_state_df42),.LO(un14_s_state_cry[42:42]));
  MUXCY_L desc3031(.DI(un14_s_state_lt40),.CI(un14_s_state_cry[38:38]),.S(un14_s_state_df40),.LO(un14_s_state_cry[40:40]));
  MUXCY_L desc3032(.DI(un14_s_state_lt38),.CI(un14_s_state_cry[36:36]),.S(un14_s_state_df38),.LO(un14_s_state_cry[38:38]));
  MUXCY_L desc3033(.DI(un14_s_state_lt36),.CI(un14_s_state_cry[34:34]),.S(un14_s_state_df36),.LO(un14_s_state_cry[36:36]));
  MUXCY_L desc3034(.DI(un14_s_state_lt34),.CI(un14_s_state_cry[32:32]),.S(un14_s_state_df34),.LO(un14_s_state_cry[34:34]));
  MUXCY_L desc3035(.DI(un14_s_state_lt32),.CI(un14_s_state_cry[30:30]),.S(un14_s_state_df32),.LO(un14_s_state_cry[32:32]));
  MUXCY_L desc3036(.DI(un14_s_state_lt30),.CI(un14_s_state_cry[28:28]),.S(un14_s_state_df30),.LO(un14_s_state_cry[30:30]));
  MUXCY_L desc3037(.DI(un14_s_state_lt28),.CI(un14_s_state_cry[26:26]),.S(un14_s_state_df28),.LO(un14_s_state_cry[28:28]));
  MUXCY_L desc3038(.DI(un14_s_state_lt26),.CI(un14_s_state_cry[24:24]),.S(un14_s_state_df26),.LO(un14_s_state_cry[26:26]));
  MUXCY_L desc3039(.DI(un14_s_state_lt24),.CI(un14_s_state_cry[22:22]),.S(un14_s_state_df24),.LO(un14_s_state_cry[24:24]));
  MUXCY_L desc3040(.DI(un14_s_state_lt22),.CI(un14_s_state_cry[20:20]),.S(un14_s_state_df22),.LO(un14_s_state_cry[22:22]));
  MUXCY_L desc3041(.DI(un14_s_state_lt20),.CI(un14_s_state_cry[18:18]),.S(un14_s_state_df20),.LO(un14_s_state_cry[20:20]));
  MUXCY_L desc3042(.DI(un14_s_state_lt18),.CI(un14_s_state_cry[16:16]),.S(un14_s_state_df18),.LO(un14_s_state_cry[18:18]));
  MUXCY_L desc3043(.DI(un14_s_state_lt16),.CI(un14_s_state_cry[14:14]),.S(un14_s_state_df16),.LO(un14_s_state_cry[16:16]));
  MUXCY_L desc3044(.DI(un14_s_state_lt14),.CI(un14_s_state_cry[12:12]),.S(un14_s_state_df14),.LO(un14_s_state_cry[14:14]));
  MUXCY_L desc3045(.DI(un14_s_state_lt12),.CI(un14_s_state_cry[10:10]),.S(un14_s_state_df12),.LO(un14_s_state_cry[12:12]));
  MUXCY_L desc3046(.DI(un14_s_state_lt10),.CI(un14_s_state_cry[8:8]),.S(un14_s_state_df10),.LO(un14_s_state_cry[10:10]));
  MUXCY_L desc3047(.DI(un14_s_state_lt8),.CI(un14_s_state_cry[6:6]),.S(un14_s_state_df8),.LO(un14_s_state_cry[8:8]));
  MUXCY_L desc3048(.DI(un14_s_state_lt6),.CI(un14_s_state_cry[4:4]),.S(un14_s_state_df6),.LO(un14_s_state_cry[6:6]));
  MUXCY_L desc3049(.DI(un14_s_state_lt4),.CI(un14_s_state_cry[2:2]),.S(un14_s_state_df4),.LO(un14_s_state_cry[4:4]));
  MUXCY_L desc3050(.DI(un14_s_state_lt2),.CI(un14_s_state_cry[0:0]),.S(un14_s_state_df2),.LO(un14_s_state_cry[2:2]));
  MUXCY_L desc3051(.DI(un14_s_state_lt0),.CI(GND),.S(un14_s_state_df0),.LO(un14_s_state_cry[0:0]));
  LUT2 un14_s_state_lt0_cZ(.I0(r0_2[1:1]),.I1(r0_2[0:0]),.O(un14_s_state_lt0));
defparam un14_s_state_lt0_cZ.INIT=4'hE;
  MUXCY_L un31_s_count_0_I_131(.DI(GND),.CI(un31_s_count_0_data_tmp[15:15]),.S(un31_s_count_0_N_4),.LO(un31_s_count_0_data_tmp[16:16]));
  MUXCY_L un31_s_count_0_I_123(.DI(GND),.CI(un31_s_count_0_data_tmp[14:14]),.S(un31_s_count_0_N_11),.LO(un31_s_count_0_data_tmp[15:15]));
  MUXCY_L un31_s_count_0_I_115(.DI(GND),.CI(un31_s_count_0_data_tmp[13:13]),.S(un31_s_count_0_N_18),.LO(un31_s_count_0_data_tmp[14:14]));
  MUXCY_L un31_s_count_0_I_107(.DI(GND),.CI(un31_s_count_0_data_tmp[12:12]),.S(un31_s_count_0_N_25),.LO(un31_s_count_0_data_tmp[13:13]));
  MUXCY_L un31_s_count_0_I_99(.DI(GND),.CI(un31_s_count_0_data_tmp[11:11]),.S(un31_s_count_0_N_32),.LO(un31_s_count_0_data_tmp[12:12]));
  MUXCY_L un31_s_count_0_I_91(.DI(GND),.CI(un31_s_count_0_data_tmp[10:10]),.S(un31_s_count_0_N_39),.LO(un31_s_count_0_data_tmp[11:11]));
  MUXCY_L un31_s_count_0_I_83(.DI(GND),.CI(un31_s_count_0_data_tmp[9:9]),.S(un31_s_count_0_N_46),.LO(un31_s_count_0_data_tmp[10:10]));
  MUXCY_L un31_s_count_0_I_75(.DI(GND),.CI(un31_s_count_0_data_tmp[8:8]),.S(un31_s_count_0_N_53),.LO(un31_s_count_0_data_tmp[9:9]));
  MUXCY_L un31_s_count_0_I_67(.DI(GND),.CI(un31_s_count_0_data_tmp[7:7]),.S(un31_s_count_0_N_60),.LO(un31_s_count_0_data_tmp[8:8]));
  MUXCY_L un31_s_count_0_I_59(.DI(GND),.CI(un31_s_count_0_data_tmp[6:6]),.S(un31_s_count_0_N_67),.LO(un31_s_count_0_data_tmp[7:7]));
  MUXCY_L un31_s_count_0_I_51(.DI(GND),.CI(un31_s_count_0_data_tmp[5:5]),.S(un31_s_count_0_N_74),.LO(un31_s_count_0_data_tmp[6:6]));
  MUXCY_L un31_s_count_0_I_43(.DI(GND),.CI(un31_s_count_0_data_tmp[4:4]),.S(un31_s_count_0_N_81),.LO(un31_s_count_0_data_tmp[5:5]));
  MUXCY_L un31_s_count_0_I_35(.DI(GND),.CI(un31_s_count_0_data_tmp[3:3]),.S(un31_s_count_0_N_88),.LO(un31_s_count_0_data_tmp[4:4]));
  MUXCY_L un31_s_count_0_I_27(.DI(GND),.CI(un31_s_count_0_data_tmp[2:2]),.S(un31_s_count_0_N_95),.LO(un31_s_count_0_data_tmp[3:3]));
  MUXCY_L un31_s_count_0_I_19(.DI(GND),.CI(un31_s_count_0_data_tmp[1:1]),.S(un31_s_count_0_N_102),.LO(un31_s_count_0_data_tmp[2:2]));
  MUXCY_L un31_s_count_0_I_11(.DI(GND),.CI(un31_s_count_0_data_tmp[0:0]),.S(un31_s_count_0_N_109),.LO(un31_s_count_0_data_tmp[1:1]));
  MUXCY_L un31_s_count_0_I_1(.DI(GND),.CI(VCC),.S(un31_s_count_0_N_116),.LO(un31_s_count_0_data_tmp[0:0]));
  FDR desc3052(.Q(b_2[40:40]),.D(b_2[42:42]),.C(clk_i),.R(s_start_i));
  FDR desc3053(.Q(b_2[42:42]),.D(b_2[44:44]),.C(clk_i),.R(s_start_i));
  FDR desc3054(.Q(b_2[44:44]),.D(b_2[46:46]),.C(clk_i),.R(s_start_i));
  FDR desc3055(.Q(b_2[46:46]),.D(b_2[48:48]),.C(clk_i),.R(s_start_i));
  FDR desc3056(.Q(b_2[48:48]),.D(b_2[50:50]),.C(clk_i),.R(s_start_i));
  FDR desc3057(.Q(b_2[38:38]),.D(b_2[40:40]),.C(clk_i),.R(s_start_i));
  FDR desc3058(.Q(b_2[36:36]),.D(b_2[38:38]),.C(clk_i),.R(s_start_i));
  FDR desc3059(.Q(b_2[34:34]),.D(b_2[36:36]),.C(clk_i),.R(s_start_i));
  FDR desc3060(.Q(b_2[32:32]),.D(b_2[34:34]),.C(clk_i),.R(s_start_i));
  FDR desc3061(.Q(b_2[30:30]),.D(b_2[32:32]),.C(clk_i),.R(s_start_i));
  FDR desc3062(.Q(b_2[28:28]),.D(b_2[30:30]),.C(clk_i),.R(s_start_i));
  FDR desc3063(.Q(b_2[26:26]),.D(b_2[28:28]),.C(clk_i),.R(s_start_i));
  FDR desc3064(.Q(b_2[24:24]),.D(b_2[26:26]),.C(clk_i),.R(s_start_i));
  FDR desc3065(.Q(b_2[22:22]),.D(b_2[24:24]),.C(clk_i),.R(s_start_i));
  FDR desc3066(.Q(b_2[20:20]),.D(b_2[22:22]),.C(clk_i),.R(s_start_i));
  FDR desc3067(.Q(b_2[18:18]),.D(b_2[20:20]),.C(clk_i),.R(s_start_i));
  FDR desc3068(.Q(b_2[16:16]),.D(b_2[18:18]),.C(clk_i),.R(s_start_i));
  FDR desc3069(.Q(b_2[14:14]),.D(b_2[16:16]),.C(clk_i),.R(s_start_i));
  FDR desc3070(.Q(b_2[12:12]),.D(b_2[14:14]),.C(clk_i),.R(s_start_i));
  FDR desc3071(.Q(b_2[10:10]),.D(b_2[12:12]),.C(clk_i),.R(s_start_i));
  FDR desc3072(.Q(b_2[8:8]),.D(b_2[10:10]),.C(clk_i),.R(s_start_i));
  FDR desc3073(.Q(b_2[6:6]),.D(b_2[8:8]),.C(clk_i),.R(s_start_i));
  FDR desc3074(.Q(b_2[4:4]),.D(b_2[6:6]),.C(clk_i),.R(s_start_i));
  FDR desc3075(.Q(b_2[2:2]),.D(b_2[4:4]),.C(clk_i),.R(s_start_i));
  FDR desc3076(.Q(b_2[0:0]),.D(b_2[2:2]),.C(clk_i),.R(s_start_i));
  FDS desc3077(.Q(b[25:25]),.D(GND),.C(clk_i),.S(s_start_i));
  FDR desc3078(.Q(b[24:24]),.D(b[25:25]),.C(clk_i),.R(s_start_i));
  FDR desc3079(.Q(b[23:23]),.D(b[24:24]),.C(clk_i),.R(s_start_i));
  FDR desc3080(.Q(b[22:22]),.D(b[23:23]),.C(clk_i),.R(s_start_i));
  FDR desc3081(.Q(b[21:21]),.D(b[22:22]),.C(clk_i),.R(s_start_i));
  FDR desc3082(.Q(b[20:20]),.D(b[21:21]),.C(clk_i),.R(s_start_i));
  FDR desc3083(.Q(b[19:19]),.D(b[20:20]),.C(clk_i),.R(s_start_i));
  FDR desc3084(.Q(b[18:18]),.D(b[19:19]),.C(clk_i),.R(s_start_i));
  FDR desc3085(.Q(b[17:17]),.D(b[18:18]),.C(clk_i),.R(s_start_i));
  FDR desc3086(.Q(b[16:16]),.D(b[17:17]),.C(clk_i),.R(s_start_i));
  FDR desc3087(.Q(b[15:15]),.D(b[16:16]),.C(clk_i),.R(s_start_i));
  FDR desc3088(.Q(b[14:14]),.D(b[15:15]),.C(clk_i),.R(s_start_i));
  FDR desc3089(.Q(b[13:13]),.D(b[14:14]),.C(clk_i),.R(s_start_i));
  FDR desc3090(.Q(b[12:12]),.D(b[13:13]),.C(clk_i),.R(s_start_i));
  FDR desc3091(.Q(b[11:11]),.D(b[12:12]),.C(clk_i),.R(s_start_i));
  FDR desc3092(.Q(b[10:10]),.D(b[11:11]),.C(clk_i),.R(s_start_i));
  FDR desc3093(.Q(b[9:9]),.D(b[10:10]),.C(clk_i),.R(s_start_i));
  FDR desc3094(.Q(b[8:8]),.D(b[9:9]),.C(clk_i),.R(s_start_i));
  FDR desc3095(.Q(b[7:7]),.D(b[8:8]),.C(clk_i),.R(s_start_i));
  FDR desc3096(.Q(b[6:6]),.D(b[7:7]),.C(clk_i),.R(s_start_i));
  FDR desc3097(.Q(b[5:5]),.D(b[6:6]),.C(clk_i),.R(s_start_i));
  FDR desc3098(.Q(b[4:4]),.D(b[5:5]),.C(clk_i),.R(s_start_i));
  FDR desc3099(.Q(b[3:3]),.D(b[4:4]),.C(clk_i),.R(s_start_i));
  FDR desc3100(.Q(b[2:2]),.D(b[3:3]),.C(clk_i),.R(s_start_i));
  FDR desc3101(.Q(b[1:1]),.D(b[2:2]),.C(clk_i),.R(s_start_i));
  FDR desc3102(.Q(b[0:0]),.D(b[1:1]),.C(clk_i),.R(s_start_i));
  FDS desc3103(.Q(c[4:4]),.D(m154_lut6_2_O6),.C(clk_i),.S(s_start_i));
  FDS desc3104(.Q(c[3:3]),.D(m154_lut6_2_O5),.C(clk_i),.S(s_start_i));
  FDR desc3105(.Q(c[2:2]),.D(m127_lut6_2_O5),.C(clk_i),.R(s_start_i));
  FDS desc3106(.Q(c[1:1]),.D(N_2),.C(clk_i),.S(s_start_i));
  FDR desc3107(.Q(c[0:0]),.D(c_i),.C(clk_i),.R(s_start_i));
  FDRE desc3108(.Q(s_sqr_o[24:24]),.D(un1_r1_s_24),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3109(.Q(s_sqr_o[23:23]),.D(un1_r1_s_23),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3110(.Q(s_sqr_o[22:22]),.D(un1_r1_s_22),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3111(.Q(s_sqr_o[21:21]),.D(un1_r1_s_21),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3112(.Q(s_sqr_o[20:20]),.D(un1_r1_s_20),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3113(.Q(s_sqr_o[19:19]),.D(un1_r1_s_19),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3114(.Q(s_sqr_o[18:18]),.D(un1_r1_s_18),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3115(.Q(s_sqr_o[17:17]),.D(un1_r1_s_17),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3116(.Q(s_sqr_o[16:16]),.D(un1_r1_s_16),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3117(.Q(s_sqr_o[15:15]),.D(un1_r1_s_15),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3118(.Q(s_sqr_o[14:14]),.D(un1_r1_s_14),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3119(.Q(s_sqr_o[13:13]),.D(un1_r1_s_13),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3120(.Q(s_sqr_o[12:12]),.D(un1_r1_s_12),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3121(.Q(s_sqr_o[11:11]),.D(un1_r1_s_11),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3122(.Q(s_sqr_o[10:10]),.D(un1_r1_s_10),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3123(.Q(s_sqr_o[9:9]),.D(un1_r1_s_9),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3124(.Q(s_sqr_o[8:8]),.D(un1_r1_s_8),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3125(.Q(s_sqr_o[7:7]),.D(un1_r1_s_7),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3126(.Q(s_sqr_o[6:6]),.D(un1_r1_s_6),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3127(.Q(s_sqr_o[5:5]),.D(un1_r1_s_5),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3128(.Q(s_sqr_o[4:4]),.D(un1_r1_s_4),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3129(.Q(s_sqr_o[3:3]),.D(un1_r1_s_3),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3130(.Q(s_sqr_o[2:2]),.D(un1_r1_s_2),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3131(.Q(s_sqr_o[1:1]),.D(un1_r1_s_1),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3132(.Q(s_sqr_o[0:0]),.D(un1_r1_axb_0),.C(clk_i),.R(s_start_i),.CE(un3_s_count_0_a2_lut6_2_O6));
  FDRE desc3133(.Q(r0[25:25]),.D(v_r1_3[25:25]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3134(.Q(r0[24:24]),.D(v_r1_3[24:24]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3135(.Q(r0[23:23]),.D(v_r1_3[23:23]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3136(.Q(r0[22:22]),.D(v_r1_3[22:22]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3137(.Q(r0[21:21]),.D(v_r1_3[21:21]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3138(.Q(r0[20:20]),.D(v_r1_3[20:20]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3139(.Q(r0[19:19]),.D(v_r1_3[19:19]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3140(.Q(r0[18:18]),.D(v_r1_3[18:18]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3141(.Q(r0[17:17]),.D(v_r1_3[17:17]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3142(.Q(r0[16:16]),.D(v_r1_3[16:16]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3143(.Q(r0[15:15]),.D(v_r1_3[15:15]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3144(.Q(r0[14:14]),.D(v_r1_3[14:14]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3145(.Q(r0[13:13]),.D(v_r1_3[13:13]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3146(.Q(r0[12:12]),.D(v_r1_3[12:12]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3147(.Q(r0[11:11]),.D(v_r1_3[11:11]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3148(.Q(r0[10:10]),.D(v_r1_3[10:10]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3149(.Q(r0[9:9]),.D(v_r1_3[9:9]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3150(.Q(r0[8:8]),.D(v_r1_3[8:8]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3151(.Q(r0[7:7]),.D(v_r1_3[7:7]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3152(.Q(r0[6:6]),.D(v_r1_3[6:6]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3153(.Q(r0[5:5]),.D(v_r1_3[5:5]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3154(.Q(r0[4:4]),.D(v_r1_3[4:4]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3155(.Q(r0[3:3]),.D(v_r1_3[3:3]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3156(.Q(r0[2:2]),.D(v_r1_3[2:2]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3157(.Q(r0[1:1]),.D(v_r1_3[1:1]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3158(.Q(r0[0:0]),.D(v_r1_3[0:0]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3159(.Q(r0_2[51:51]),.D(v_r1_2_3[51:51]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3160(.Q(r0_2[50:50]),.D(v_r1_2_3[50:50]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3161(.Q(r0_2[49:49]),.D(v_r1_2_3[49:49]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3162(.Q(r0_2[48:48]),.D(v_r1_2_3[48:48]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3163(.Q(r0_2[47:47]),.D(v_r1_2_3[47:47]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3164(.Q(r0_2[46:46]),.D(v_r1_2_3[46:46]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3165(.Q(r0_2[45:45]),.D(v_r1_2_3[45:45]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3166(.Q(r0_2[44:44]),.D(v_r1_2_3[44:44]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3167(.Q(r0_2[43:43]),.D(v_r1_2_3[43:43]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3168(.Q(r0_2[42:42]),.D(v_r1_2_3[42:42]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3169(.Q(r0_2[41:41]),.D(v_r1_2_3[41:41]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3170(.Q(r0_2[40:40]),.D(v_r1_2_3[40:40]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3171(.Q(r0_2[39:39]),.D(v_r1_2_3[39:39]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3172(.Q(r0_2[38:38]),.D(v_r1_2_3[38:38]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3173(.Q(r0_2[37:37]),.D(v_r1_2_3[37:37]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3174(.Q(r0_2[36:36]),.D(v_r1_2_3[36:36]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3175(.Q(r0_2[35:35]),.D(v_r1_2_3[35:35]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3176(.Q(r0_2[34:34]),.D(v_r1_2_3[34:34]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3177(.Q(r0_2[33:33]),.D(v_r1_2_3[33:33]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3178(.Q(r0_2[32:32]),.D(v_r1_2_3[32:32]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3179(.Q(r0_2[31:31]),.D(v_r1_2_3[31:31]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3180(.Q(r0_2[30:30]),.D(v_r1_2_3[30:30]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3181(.Q(r0_2[29:29]),.D(v_r1_2_3[29:29]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3182(.Q(r0_2[28:28]),.D(v_r1_2_3[28:28]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3183(.Q(r0_2[27:27]),.D(v_r1_2_3[27:27]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3184(.Q(r0_2[26:26]),.D(v_r1_2_3[26:26]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3185(.Q(r0_2[25:25]),.D(v_r1_2_3[25:25]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3186(.Q(r0_2[24:24]),.D(v_r1_2_3[24:24]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3187(.Q(r0_2[23:23]),.D(v_r1_2_3[23:23]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3188(.Q(r0_2[22:22]),.D(v_r1_2_3[22:22]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3189(.Q(r0_2[21:21]),.D(v_r1_2_3[21:21]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3190(.Q(r0_2[20:20]),.D(v_r1_2_3[20:20]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3191(.Q(r0_2[19:19]),.D(v_r1_2_3[19:19]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3192(.Q(r0_2[18:18]),.D(v_r1_2_3[18:18]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3193(.Q(r0_2[17:17]),.D(v_r1_2_3[17:17]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3194(.Q(r0_2[16:16]),.D(v_r1_2_3[16:16]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3195(.Q(r0_2[15:15]),.D(v_r1_2_3[15:15]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3196(.Q(r0_2[14:14]),.D(v_r1_2_3[14:14]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3197(.Q(r0_2[13:13]),.D(v_r1_2_3[13:13]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3198(.Q(r0_2[12:12]),.D(v_r1_2_3[12:12]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3199(.Q(r0_2[11:11]),.D(v_r1_2_3[11:11]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3200(.Q(r0_2[10:10]),.D(v_r1_2_3[10:10]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3201(.Q(r0_2[9:9]),.D(v_r1_2_3[9:9]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3202(.Q(r0_2[8:8]),.D(v_r1_2_3[8:8]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3203(.Q(r0_2[7:7]),.D(v_r1_2_3[7:7]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3204(.Q(r0_2[6:6]),.D(v_r1_2_3[6:6]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3205(.Q(r0_2[5:5]),.D(v_r1_2_3[5:5]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3206(.Q(r0_2[4:4]),.D(v_r1_2_3[4:4]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3207(.Q(r0_2[3:3]),.D(v_r1_2_3[3:3]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3208(.Q(r0_2[2:2]),.D(v_r1_2_3[2:2]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3209(.Q(r0_2[1:1]),.D(v_r1_2_3[1:1]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  FDRE desc3210(.Q(r0_2[0:0]),.D(v_r1_2_3[0:0]),.C(clk_i),.R(s_start_i),.CE(s_state_0));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT5 desc3211(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_964_i));
defparam desc3211.INIT=32'hE1E1E1E0;
  LUT5 desc3212(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_963_i));
defparam desc3212.INIT=32'h55555554;
  LUT4 desc3213(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.O(N_980_i));
defparam desc3213.INIT=16'hFE01;
  LUT5 desc3214(.I0(s_count[0:0]),.I1(s_count[1:1]),.I2(s_count[2:2]),.I3(s_count[3:3]),.I4(s_count[4:4]),.O(N_981_i));
defparam desc3214.INIT=32'hFFFE0001;
  LUT2 v_r1_2_3_21_2_RNIQ1CU_o6(.I0(r0_2[8:8]),.I1(r0_2[7:7]),.O(v_r1_2_3_27_0));
defparam v_r1_2_3_21_2_RNIQ1CU_o6.INIT=4'h8;
  LUT5 v_r1_2_3_21_2_RNIQ1CU_o5(.I0(b_2[8:8]),.I1(r0_2[8:8]),.I2(r0_2[7:7]),.I3(r0_2[9:9]),.I4(v_r1_2_3_21_2),.O(v_r1_2_3_21_2_RNIQ1CU_O5));
defparam v_r1_2_3_21_2_RNIQ1CU_o5.INIT=32'hE8008800;
  LUT4 desc3215(.I0(r0_2[14:14]),.I1(r0_2[13:13]),.I2(r0_2[16:16]),.I3(r0_2[15:15]),.O(g0_0_a3_0_2));
defparam desc3215.INIT=16'h8000;
  LUT3 desc3216(.I0(b_2[14:14]),.I1(r0_2[16:16]),.I2(r0_2[15:15]),.O(g1_1_1));
defparam desc3216.INIT=8'h80;
  LUT2 desc3217(.I0(r0_2[10:10]),.I1(r0_2[9:9]),.O(g4_0_0_1));
defparam desc3217.INIT=4'h8;
  LUT2 desc3218(.I0(r0_2[10:10]),.I1(r0_2[9:9]),.O(v_r1_2_3_34_0));
defparam desc3218.INIT=4'h8;
  LUT4 desc3219(.I0(r0_2[21:21]),.I1(c[4:4]),.I2(m191),.I3(m176),.O(r0_2_RNI9011F_O6[22:22]));
defparam desc3219.INIT=16'h6A59;
  LUT2 desc3220(.I0(r0_2[22:22]),.I1(r0_2[21:21]),.O(g0_0_2));
defparam desc3220.INIT=4'h8;
  LUT2 desc3221(.I0(b_2[18:18]),.I1(r0_2[19:19]),.O(g4_0_1));
defparam desc3221.INIT=4'h8;
  LUT2 desc3222(.I0(r0_2[19:19]),.I1(r0_2[18:18]),.O(g0_6_0));
defparam desc3222.INIT=4'h8;
  LUT2 desc3223(.I0(b_2[18:18]),.I1(r0_2[19:19]),.O(g4_0_0));
defparam desc3223.INIT=4'h8;
  LUT2 desc3224(.I0(b_2[18:18]),.I1(r0_2[19:19]),.O(g1_0_0_1));
defparam desc3224.INIT=4'h8;
  LUT2 desc3225(.I0(b_2[14:14]),.I1(r0_2[15:15]),.O(g1_0_0_2));
defparam desc3225.INIT=4'h8;
  LUT3 desc3226(.I0(r0_2[16:16]),.I1(r0_2[17:17]),.I2(r0_2[15:15]),.O(g0_0_a4_0_1));
defparam desc3226.INIT=8'h80;
  LUT2 v_r1_2_3_35_0_RNI40J52_o6(.I0(r0_2[10:10]),.I1(r0_2[9:9]),.O(g0_0_a4_0_2));
defparam v_r1_2_3_35_0_RNI40J52_o6.INIT=4'h8;
  LUT5 v_r1_2_3_35_0_RNI40J52_o5(.I0(r0_2[10:10]),.I1(r0_2[11:11]),.I2(r0_2[9:9]),.I3(v_r1_2_3_35_0),.I4(v_r1_2_3_21_2_RNIMLGQ),.O(v_r1_2_3_35_0_RNI40J52_O5));
defparam v_r1_2_3_35_0_RNI40J52_o5.INIT=32'hCC80CC00;
  LUT2 v_r1_2_3_73_0_lut6_2_o6(.I0(b_2[22:22]),.I1(r0_2[22:22]),.O(v_r1_2_3_73_0));
defparam v_r1_2_3_73_0_lut6_2_o6.INIT=4'h6;
  LUT5 v_r1_2_3_73_0_lut6_2_o5(.I0(r0_2[23:23]),.I1(b_2[22:22]),.I2(r0_2[22:22]),.I3(r0_2[21:21]),.I4(r0_2[20:20]),.O(v_r1_2_3_73_0_lut6_2_O5));
defparam v_r1_2_3_73_0_lut6_2_o5.INIT=32'hA8808080;
  LUT2 v_r1_2_3_59_0_lut6_2_o6(.I0(b_2[18:18]),.I1(r0_2[18:18]),.O(v_r1_2_3_59_0));
defparam v_r1_2_3_59_0_lut6_2_o6.INIT=4'h6;
  LUT5 v_r1_2_3_59_0_lut6_2_o5(.I0(b_2[18:18]),.I1(r0_2[20:20]),.I2(r0_2[19:19]),.I3(r0_2[18:18]),.I4(r0_2[17:17]),.O(g0_i_1));
defparam v_r1_2_3_59_0_lut6_2_o5.INIT=32'hC0808000;
  LUT2 v_r1_2_3_52_0_lut6_2_o6(.I0(b_2[16:16]),.I1(r0_2[16:16]),.O(v_r1_2_3_52_0));
defparam v_r1_2_3_52_0_lut6_2_o6.INIT=4'h6;
  LUT2 v_r1_2_3_52_0_lut6_2_o5(.I0(b_2[16:16]),.I1(r0_2[17:17]),.O(g0_0_a4_0));
defparam v_r1_2_3_52_0_lut6_2_o5.INIT=4'h8;
  LUT5 v_r1_2_3_44_lut6_2_o6(.I0(r0_2[12:12]),.I1(r0_2[11:11]),.I2(r0_2[13:13]),.I3(b_2_RNIMF314[10:10]),.I4(v_r1_2_3_42_0),.O(v_r1_2_3_44_lut6_2_O6));
defparam v_r1_2_3_44_lut6_2_o6.INIT=32'hF0F08000;
  LUT2 v_r1_2_3_44_lut6_2_o5(.I0(r0_2[12:12]),.I1(r0_2[11:11]),.O(v_r1_2_3_41_0));
defparam v_r1_2_3_44_lut6_2_o5.INIT=4'h8;
  LUT2 desc3227(.I0(r0_2[10:10]),.I1(r0_2[9:9]),.O(g4_0_2));
defparam desc3227.INIT=4'h8;
  LUT2 desc3228(.I0(b_2[10:10]),.I1(r0_2[10:10]),.O(v_r1_2_3_31_0));
defparam desc3228.INIT=4'h6;
  LUT2 un12_s_state_0_a2_lut6_2_o6(.I0(s_state_0),.I1(s_start_i),.O(un12_s_state_0_a2_lut6_2_O6));
defparam un12_s_state_0_a2_lut6_2_o6.INIT=4'h2;
  LUT2 un12_s_state_0_a2_lut6_2_o5(.I0(s_state),.I1(s_start_i),.O(un12_s_state_0_a2_lut6_2_O5));
defparam un12_s_state_0_a2_lut6_2_o5.INIT=4'h2;
  LUT3 un33_s_count_a_5_0_axb_2_lut6_2_o6(.I0(r1[1:1]),.I1(r1_2[2:2]),.I2(r1_2[1:1]),.O(un33_s_count_a_5_0_axb_2));
defparam un33_s_count_a_5_0_axb_2_lut6_2_o6.INIT=8'h96;
  LUT2 un33_s_count_a_5_0_axb_2_lut6_2_o5(.I0(r1[1:1]),.I1(r1_2[2:2]),.O(un33_s_count_a_5_0_axb_2_lut6_2_O5));
defparam un33_s_count_a_5_0_axb_2_lut6_2_o5.INIT=4'hD;
  LUT4 desc3229(.I0(r1[25:25]),.I1(r1[24:24]),.I2(r1_2[26:26]),.I3(r1_2[25:25]),.O(un33_s_count_a_5_0_axb_26));
defparam desc3229.INIT=16'hA569;
  LUT2 desc3230(.I0(r1[25:25]),.I1(r1_2[26:26]),.O(r1_RNIABVR_O5[25:25]));
defparam desc3230.INIT=4'hD;
  LUT4 desc3231(.I0(r0[4:4]),.I1(r0[3:3]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m55_lut6_2_O6));
defparam desc3231.INIT=16'h35CA;
  LUT4 desc3232(.I0(r0[4:4]),.I1(r0[5:5]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m55_lut6_2_O5));
defparam desc3232.INIT=16'h53AC;
  LUT4 desc3233(.I0(r0[20:20]),.I1(r0[19:19]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(N_18_1));
defparam desc3233.INIT=16'h35CA;
  LUT4 desc3234(.I0(r0[20:20]),.I1(r0[21:21]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m17_lut6_2_O5));
defparam desc3234.INIT=16'h53AC;
  LUT4 desc3235(.I0(r0[23:23]),.I1(r0[24:24]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(N_10_1));
defparam desc3235.INIT=16'h53AC;
  LUT4 desc3236(.I0(r0[24:24]),.I1(r0[25:25]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m9_lut6_2_O5));
defparam desc3236.INIT=16'h53AC;
  LUT4 desc3237(.I0(r0[16:16]),.I1(r0[15:15]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m24_lut6_2_O6));
defparam desc3237.INIT=16'h35CA;
  LUT3 desc3238(.I0(r0[25:25]),.I1(c[0:0]),.I2(un14_s_state_cry[50:50]),.O(m24_lut6_2_O5));
defparam desc3238.INIT=8'h78;
  LUT4 desc3239(.I0(r0[1:1]),.I1(r0[0:0]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m138_lut6_2_O6));
defparam desc3239.INIT=16'h35CA;
  LUT5 desc3240(.I0(r0[1:1]),.I1(r0[0:0]),.I2(c[1:1]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.O(m138_lut6_2_O5));
defparam desc3240.INIT=32'h0C0AF3F5;
  LUT5 desc3241(.I0(c[1:1]),.I1(c[2:2]),.I2(c[0:0]),.I3(c[3:3]),.I4(c[4:4]),.O(m154_lut6_2_O6));
defparam desc3241.INIT=32'hFFFE0001;
  LUT4 desc3242(.I0(c[1:1]),.I1(c[2:2]),.I2(c[0:0]),.I3(c[3:3]),.O(m154_lut6_2_O5));
defparam desc3242.INIT=16'hFE01;
  LUT4 desc3243(.I0(r0[0:0]),.I1(c[1:1]),.I2(c[0:0]),.I3(un14_s_state_cry[50:50]),.O(m127_lut6_2_O6));
defparam desc3243.INIT=16'h02FD;
  LUT3 desc3244(.I0(c[1:1]),.I1(c[2:2]),.I2(c[0:0]),.O(m127_lut6_2_O5));
defparam desc3244.INIT=8'hC9;
  LUT5 un3_s_count_0_a2_lut6_2_o6(.I0(s_count[4:4]),.I1(s_count[2:2]),.I2(s_count[3:3]),.I3(s_count[0:0]),.I4(s_count[1:1]),.O(un3_s_count_0_a2_lut6_2_O6));
defparam un3_s_count_0_a2_lut6_2_o6.INIT=32'h00000001;
  LUT2 un3_s_count_0_a2_lut6_2_o5(.I0(s_count[0:0]),.I1(s_count[1:1]),.O(N_22_i_i));
defparam un3_s_count_0_a2_lut6_2_o5.INIT=4'h9;
  LUT5 desc3245(.I0(r0[25:25]),.I1(c[1:1]),.I2(c[2:2]),.I3(c[0:0]),.I4(un14_s_state_cry[50:50]),.O(N_83_0));
defparam desc3245.INIT=32'h7FFF8000;
  LUT2 desc3246(.I0(c[1:1]),.I1(c[0:0]),.O(N_2));
defparam desc3246.INIT=4'h9;
  LUT3 desc3247(.I0(c[2:2]),.I1(N_19_1),.I2(m25),.O(m26_lut6_2_O6));
defparam desc3247.INIT=8'hE4;
  LUT3 desc3248(.I0(c[2:2]),.I1(N_84_0),.I2(m84),.O(N_86_0));
defparam desc3248.INIT=8'hE4;
  LUT5 desc3249(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m136),.I4(m139),.O(m141_lut6_2_O6));
defparam desc3249.INIT=32'h0C1D2E3F;
  LUT4 desc3250(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m139),.O(m141_lut6_2_O5));
defparam desc3250.INIT=16'h0E1F;
  LUT5 desc3251(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m65),.I4(m56),.O(m73_lut6_2_O6));
defparam desc3251.INIT=32'h2E0C3F1D;
  LUT4 desc3252(.I0(c[2:2]),.I1(c[3:3]),.I2(un14_s_state_cry[50:50]),.I3(m65),.O(m73_lut6_2_O5));
defparam desc3252.INIT=16'h1F0E;
  LUT3 desc3253(.I0(c[4:4]),.I1(m189),.I2(m171),.O(m190_lut6_2_O6));
defparam desc3253.INIT=8'h8D;
  LUT3 desc3254(.I0(c[4:4]),.I1(un14_s_state_cry[50:50]),.I2(m171),.O(m190_lut6_2_O5));
defparam desc3254.INIT=8'hE4;
  LUT3 desc3255(.I0(c[4:4]),.I1(m186),.I2(m166),.O(m187_lut6_2_O6));
defparam desc3255.INIT=8'h8D;
  LUT3 desc3256(.I0(c[4:4]),.I1(un14_s_state_cry[50:50]),.I2(m166),.O(m187_lut6_2_O5));
defparam desc3256.INIT=8'hE4;
  LUT5 desc3257(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m47),.I4(N_50_0),.O(m168_lut6_2_O6));
defparam desc3257.INIT=32'hFCB87430;
  LUT4 desc3258(.I0(c[3:3]),.I1(c[4:4]),.I2(un14_s_state_cry[50:50]),.I3(m47),.O(m168_lut6_2_O5));
defparam desc3258.INIT=16'hF870;
  LUT3 desc3259(.I0(c[4:4]),.I1(m143),.I2(m121),.O(N_48_i));
defparam desc3259.INIT=8'h72;
  LUT3 desc3260(.I0(c[4:4]),.I1(m159),.I2(m180),.O(N_48_i_lut6_2_O5));
defparam desc3260.INIT=8'hE4;
  LUT4 un27_s_count_df50_lut6_2_o6(.I0(r1_2[51:51]),.I1(r1_2[50:50]),.I2(s_rad_i[51:51]),.I3(s_rad_i[50:50]),.O(un27_s_count_df50));
defparam un27_s_count_df50_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df50_lut6_2_o5(.I0(r1_2[51:51]),.I1(r1_2[50:50]),.I2(s_rad_i[51:51]),.I3(s_rad_i[50:50]),.O(un27_s_count_lt50));
defparam un27_s_count_df50_lut6_2_o5.INIT=16'h0A8E;
  LUT4 un27_s_count_df48_lut6_2_o6(.I0(r1_2[48:48]),.I1(r1_2[49:49]),.I2(s_rad_i[48:48]),.I3(s_rad_i[49:49]),.O(un27_s_count_df48));
defparam un27_s_count_df48_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df48_lut6_2_o5(.I0(r1_2[48:48]),.I1(r1_2[49:49]),.I2(s_rad_i[48:48]),.I3(s_rad_i[49:49]),.O(un27_s_count_lt48));
defparam un27_s_count_df48_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df46_lut6_2_o6(.I0(r1_2[46:46]),.I1(r1_2[47:47]),.I2(s_rad_i[46:46]),.I3(s_rad_i[47:47]),.O(un27_s_count_df46));
defparam un27_s_count_df46_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df46_lut6_2_o5(.I0(r1_2[46:46]),.I1(r1_2[47:47]),.I2(s_rad_i[46:46]),.I3(s_rad_i[47:47]),.O(un27_s_count_lt46));
defparam un27_s_count_df46_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df44_lut6_2_o6(.I0(r1_2[44:44]),.I1(r1_2[45:45]),.I2(s_rad_i[44:44]),.I3(s_rad_i[45:45]),.O(un27_s_count_df44));
defparam un27_s_count_df44_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df44_lut6_2_o5(.I0(r1_2[44:44]),.I1(r1_2[45:45]),.I2(s_rad_i[44:44]),.I3(s_rad_i[45:45]),.O(un27_s_count_lt44));
defparam un27_s_count_df44_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df42_lut6_2_o6(.I0(r1_2[42:42]),.I1(r1_2[43:43]),.I2(s_rad_i[42:42]),.I3(s_rad_i[43:43]),.O(un27_s_count_df42));
defparam un27_s_count_df42_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df42_lut6_2_o5(.I0(r1_2[42:42]),.I1(r1_2[43:43]),.I2(s_rad_i[42:42]),.I3(s_rad_i[43:43]),.O(un27_s_count_lt42));
defparam un27_s_count_df42_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df40_lut6_2_o6(.I0(r1_2[40:40]),.I1(r1_2[41:41]),.I2(s_rad_i[40:40]),.I3(s_rad_i[41:41]),.O(un27_s_count_df40));
defparam un27_s_count_df40_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df40_lut6_2_o5(.I0(r1_2[40:40]),.I1(r1_2[41:41]),.I2(s_rad_i[40:40]),.I3(s_rad_i[41:41]),.O(un27_s_count_lt40));
defparam un27_s_count_df40_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df38_lut6_2_o6(.I0(r1_2[38:38]),.I1(r1_2[39:39]),.I2(s_rad_i[38:38]),.I3(s_rad_i[39:39]),.O(un27_s_count_df38));
defparam un27_s_count_df38_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df38_lut6_2_o5(.I0(r1_2[38:38]),.I1(r1_2[39:39]),.I2(s_rad_i[38:38]),.I3(s_rad_i[39:39]),.O(un27_s_count_lt38));
defparam un27_s_count_df38_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df36_lut6_2_o6(.I0(r1_2[36:36]),.I1(r1_2[37:37]),.I2(s_rad_i[36:36]),.I3(s_rad_i[37:37]),.O(un27_s_count_df36));
defparam un27_s_count_df36_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df36_lut6_2_o5(.I0(r1_2[36:36]),.I1(r1_2[37:37]),.I2(s_rad_i[36:36]),.I3(s_rad_i[37:37]),.O(un27_s_count_lt36));
defparam un27_s_count_df36_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df34_lut6_2_o6(.I0(r1_2[34:34]),.I1(r1_2[35:35]),.I2(s_rad_i[34:34]),.I3(s_rad_i[35:35]),.O(un27_s_count_df34));
defparam un27_s_count_df34_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df34_lut6_2_o5(.I0(r1_2[34:34]),.I1(r1_2[35:35]),.I2(s_rad_i[34:34]),.I3(s_rad_i[35:35]),.O(un27_s_count_lt34));
defparam un27_s_count_df34_lut6_2_o5.INIT=16'h08CE;
  LUT4 un27_s_count_df32_lut6_2_o6(.I0(s_rad_i[32:32]),.I1(s_rad_i[33:33]),.I2(r1_2[32:32]),.I3(r1_2[33:33]),.O(un27_s_count_df32));
defparam un27_s_count_df32_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df32_lut6_2_o5(.I0(s_rad_i[32:32]),.I1(s_rad_i[33:33]),.I2(r1_2[32:32]),.I3(r1_2[33:33]),.O(un27_s_count_lt32));
defparam un27_s_count_df32_lut6_2_o5.INIT=16'h7310;
  LUT4 un27_s_count_df30_lut6_2_o6(.I0(s_rad_i[30:30]),.I1(s_rad_i[31:31]),.I2(r1_2[30:30]),.I3(r1_2[31:31]),.O(un27_s_count_df30));
defparam un27_s_count_df30_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df30_lut6_2_o5(.I0(s_rad_i[30:30]),.I1(s_rad_i[31:31]),.I2(r1_2[30:30]),.I3(r1_2[31:31]),.O(un27_s_count_lt30));
defparam un27_s_count_df30_lut6_2_o5.INIT=16'h7310;
  LUT4 un27_s_count_df28_lut6_2_o6(.I0(s_rad_i[29:29]),.I1(r1_2[28:28]),.I2(r1_2[29:29]),.I3(s_rad_i[28:28]),.O(un27_s_count_df28));
defparam un27_s_count_df28_lut6_2_o6.INIT=16'h8421;
  LUT4 un27_s_count_df28_lut6_2_o5(.I0(s_rad_i[29:29]),.I1(r1_2[28:28]),.I2(r1_2[29:29]),.I3(s_rad_i[28:28]),.O(un27_s_count_lt28));
defparam un27_s_count_df28_lut6_2_o5.INIT=16'h50D4;
  LUT3 un27_s_count_df26_lut6_2_o6(.I0(r1_2[26:26]),.I1(r1_2[27:27]),.I2(s_rad_i[27:27]),.O(un27_s_count_df26));
defparam un27_s_count_df26_lut6_2_o6.INIT=8'h41;
  LUT3 un27_s_count_df26_lut6_2_o5(.I0(r1_2[26:26]),.I1(r1_2[27:27]),.I2(s_rad_i[27:27]),.O(un27_s_count_lt26));
defparam un27_s_count_df26_lut6_2_o5.INIT=8'h8E;
  LUT2 un27_s_count_df24_lut6_2_o6(.I0(r1_2[24:24]),.I1(r1_2[25:25]),.O(un27_s_count_df24));
defparam un27_s_count_df24_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df24_lut6_2_o5(.I0(r1_2[24:24]),.I1(r1_2[25:25]),.O(un27_s_count_lt24));
defparam un27_s_count_df24_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df22_lut6_2_o6(.I0(r1_2[22:22]),.I1(r1_2[23:23]),.O(un27_s_count_df22));
defparam un27_s_count_df22_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df22_lut6_2_o5(.I0(r1_2[22:22]),.I1(r1_2[23:23]),.O(un27_s_count_lt22));
defparam un27_s_count_df22_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df20_lut6_2_o6(.I0(r1_2[20:20]),.I1(r1_2[21:21]),.O(un27_s_count_df20));
defparam un27_s_count_df20_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df20_lut6_2_o5(.I0(r1_2[20:20]),.I1(r1_2[21:21]),.O(un27_s_count_lt20));
defparam un27_s_count_df20_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df18_lut6_2_o6(.I0(r1_2[18:18]),.I1(r1_2[19:19]),.O(un27_s_count_df18));
defparam un27_s_count_df18_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df18_lut6_2_o5(.I0(r1_2[18:18]),.I1(r1_2[19:19]),.O(un27_s_count_lt18));
defparam un27_s_count_df18_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df16_lut6_2_o6(.I0(r1_2[16:16]),.I1(r1_2[17:17]),.O(un27_s_count_df16));
defparam un27_s_count_df16_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df16_lut6_2_o5(.I0(r1_2[16:16]),.I1(r1_2[17:17]),.O(un27_s_count_lt16));
defparam un27_s_count_df16_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df14_lut6_2_o6(.I0(r1_2[14:14]),.I1(r1_2[15:15]),.O(un27_s_count_df14));
defparam un27_s_count_df14_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df14_lut6_2_o5(.I0(r1_2[14:14]),.I1(r1_2[15:15]),.O(un27_s_count_lt14));
defparam un27_s_count_df14_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df12_lut6_2_o6(.I0(r1_2[12:12]),.I1(r1_2[13:13]),.O(un27_s_count_df12));
defparam un27_s_count_df12_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df12_lut6_2_o5(.I0(r1_2[12:12]),.I1(r1_2[13:13]),.O(un27_s_count_lt12));
defparam un27_s_count_df12_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df10_lut6_2_o6(.I0(r1_2[10:10]),.I1(r1_2[11:11]),.O(un27_s_count_df10));
defparam un27_s_count_df10_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df10_lut6_2_o5(.I0(r1_2[10:10]),.I1(r1_2[11:11]),.O(un27_s_count_lt10));
defparam un27_s_count_df10_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df8_lut6_2_o6(.I0(r1_2[8:8]),.I1(r1_2[9:9]),.O(un27_s_count_df8));
defparam un27_s_count_df8_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df8_lut6_2_o5(.I0(r1_2[8:8]),.I1(r1_2[9:9]),.O(un27_s_count_lt8));
defparam un27_s_count_df8_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df6_lut6_2_o6(.I0(r1_2[6:6]),.I1(r1_2[7:7]),.O(un27_s_count_df6));
defparam un27_s_count_df6_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df6_lut6_2_o5(.I0(r1_2[6:6]),.I1(r1_2[7:7]),.O(un27_s_count_lt6));
defparam un27_s_count_df6_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df4_lut6_2_o6(.I0(r1_2[4:4]),.I1(r1_2[5:5]),.O(un27_s_count_df4));
defparam un27_s_count_df4_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df4_lut6_2_o5(.I0(r1_2[4:4]),.I1(r1_2[5:5]),.O(un27_s_count_lt4));
defparam un27_s_count_df4_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df2_lut6_2_o6(.I0(r1_2[2:2]),.I1(r1_2[3:3]),.O(un27_s_count_df2));
defparam un27_s_count_df2_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df2_lut6_2_o5(.I0(r1_2[2:2]),.I1(r1_2[3:3]),.O(un27_s_count_lt2));
defparam un27_s_count_df2_lut6_2_o5.INIT=4'hE;
  LUT2 un27_s_count_df0_lut6_2_o6(.I0(r1_2[0:0]),.I1(r1_2[1:1]),.O(un27_s_count_df0));
defparam un27_s_count_df0_lut6_2_o6.INIT=4'h1;
  LUT2 un27_s_count_df0_lut6_2_o5(.I0(r1_2[0:0]),.I1(r1_2[1:1]),.O(un27_s_count_lt0));
defparam un27_s_count_df0_lut6_2_o5.INIT=4'hE;
  LUT4 un14_s_state_df50_lut6_2_o6(.I0(r0_2[51:51]),.I1(r0_2[50:50]),.I2(s_rad_i[51:51]),.I3(s_rad_i[50:50]),.O(un14_s_state_df50));
defparam un14_s_state_df50_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df50_lut6_2_o5(.I0(r0_2[51:51]),.I1(r0_2[50:50]),.I2(s_rad_i[51:51]),.I3(s_rad_i[50:50]),.O(un14_s_state_lt50));
defparam un14_s_state_df50_lut6_2_o5.INIT=16'h0A8E;
  LUT4 un14_s_state_df48_lut6_2_o6(.I0(r0_2[48:48]),.I1(r0_2[49:49]),.I2(s_rad_i[48:48]),.I3(s_rad_i[49:49]),.O(un14_s_state_df48));
defparam un14_s_state_df48_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df48_lut6_2_o5(.I0(r0_2[48:48]),.I1(r0_2[49:49]),.I2(s_rad_i[48:48]),.I3(s_rad_i[49:49]),.O(un14_s_state_lt48));
defparam un14_s_state_df48_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df46_lut6_2_o6(.I0(r0_2[46:46]),.I1(r0_2[47:47]),.I2(s_rad_i[46:46]),.I3(s_rad_i[47:47]),.O(un14_s_state_df46));
defparam un14_s_state_df46_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df46_lut6_2_o5(.I0(r0_2[46:46]),.I1(r0_2[47:47]),.I2(s_rad_i[46:46]),.I3(s_rad_i[47:47]),.O(un14_s_state_lt46));
defparam un14_s_state_df46_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df44_lut6_2_o6(.I0(r0_2[44:44]),.I1(r0_2[45:45]),.I2(s_rad_i[44:44]),.I3(s_rad_i[45:45]),.O(un14_s_state_df44));
defparam un14_s_state_df44_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df44_lut6_2_o5(.I0(r0_2[44:44]),.I1(r0_2[45:45]),.I2(s_rad_i[44:44]),.I3(s_rad_i[45:45]),.O(un14_s_state_lt44));
defparam un14_s_state_df44_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df42_lut6_2_o6(.I0(r0_2[42:42]),.I1(r0_2[43:43]),.I2(s_rad_i[42:42]),.I3(s_rad_i[43:43]),.O(un14_s_state_df42));
defparam un14_s_state_df42_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df42_lut6_2_o5(.I0(r0_2[42:42]),.I1(r0_2[43:43]),.I2(s_rad_i[42:42]),.I3(s_rad_i[43:43]),.O(un14_s_state_lt42));
defparam un14_s_state_df42_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df40_lut6_2_o6(.I0(r0_2[40:40]),.I1(r0_2[41:41]),.I2(s_rad_i[40:40]),.I3(s_rad_i[41:41]),.O(un14_s_state_df40));
defparam un14_s_state_df40_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df40_lut6_2_o5(.I0(r0_2[40:40]),.I1(r0_2[41:41]),.I2(s_rad_i[40:40]),.I3(s_rad_i[41:41]),.O(un14_s_state_lt40));
defparam un14_s_state_df40_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df38_lut6_2_o6(.I0(r0_2[38:38]),.I1(r0_2[39:39]),.I2(s_rad_i[38:38]),.I3(s_rad_i[39:39]),.O(un14_s_state_df38));
defparam un14_s_state_df38_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df38_lut6_2_o5(.I0(r0_2[38:38]),.I1(r0_2[39:39]),.I2(s_rad_i[38:38]),.I3(s_rad_i[39:39]),.O(un14_s_state_lt38));
defparam un14_s_state_df38_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df36_lut6_2_o6(.I0(r0_2[36:36]),.I1(r0_2[37:37]),.I2(s_rad_i[36:36]),.I3(s_rad_i[37:37]),.O(un14_s_state_df36));
defparam un14_s_state_df36_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df36_lut6_2_o5(.I0(r0_2[36:36]),.I1(r0_2[37:37]),.I2(s_rad_i[36:36]),.I3(s_rad_i[37:37]),.O(un14_s_state_lt36));
defparam un14_s_state_df36_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df34_lut6_2_o6(.I0(r0_2[34:34]),.I1(r0_2[35:35]),.I2(s_rad_i[34:34]),.I3(s_rad_i[35:35]),.O(un14_s_state_df34));
defparam un14_s_state_df34_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df34_lut6_2_o5(.I0(r0_2[34:34]),.I1(r0_2[35:35]),.I2(s_rad_i[34:34]),.I3(s_rad_i[35:35]),.O(un14_s_state_lt34));
defparam un14_s_state_df34_lut6_2_o5.INIT=16'h08CE;
  LUT4 un14_s_state_df32_lut6_2_o6(.I0(s_rad_i[32:32]),.I1(s_rad_i[33:33]),.I2(r0_2[32:32]),.I3(r0_2[33:33]),.O(un14_s_state_df32));
defparam un14_s_state_df32_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df32_lut6_2_o5(.I0(s_rad_i[32:32]),.I1(s_rad_i[33:33]),.I2(r0_2[32:32]),.I3(r0_2[33:33]),.O(un14_s_state_lt32));
defparam un14_s_state_df32_lut6_2_o5.INIT=16'h7310;
  LUT4 un14_s_state_df30_lut6_2_o6(.I0(s_rad_i[30:30]),.I1(s_rad_i[31:31]),.I2(r0_2[30:30]),.I3(r0_2[31:31]),.O(un14_s_state_df30));
defparam un14_s_state_df30_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df30_lut6_2_o5(.I0(s_rad_i[30:30]),.I1(s_rad_i[31:31]),.I2(r0_2[30:30]),.I3(r0_2[31:31]),.O(un14_s_state_lt30));
defparam un14_s_state_df30_lut6_2_o5.INIT=16'h7310;
  LUT4 un14_s_state_df28_lut6_2_o6(.I0(s_rad_i[29:29]),.I1(r0_2[28:28]),.I2(r0_2[29:29]),.I3(s_rad_i[28:28]),.O(un14_s_state_df28));
defparam un14_s_state_df28_lut6_2_o6.INIT=16'h8421;
  LUT4 un14_s_state_df28_lut6_2_o5(.I0(s_rad_i[29:29]),.I1(r0_2[28:28]),.I2(r0_2[29:29]),.I3(s_rad_i[28:28]),.O(un14_s_state_lt28));
defparam un14_s_state_df28_lut6_2_o5.INIT=16'h50D4;
  LUT3 un14_s_state_df26_lut6_2_o6(.I0(r0_2[26:26]),.I1(r0_2[27:27]),.I2(s_rad_i[27:27]),.O(un14_s_state_df26));
defparam un14_s_state_df26_lut6_2_o6.INIT=8'h41;
  LUT3 un14_s_state_df26_lut6_2_o5(.I0(r0_2[26:26]),.I1(r0_2[27:27]),.I2(s_rad_i[27:27]),.O(un14_s_state_lt26));
defparam un14_s_state_df26_lut6_2_o5.INIT=8'h8E;
  LUT2 un14_s_state_df24_lut6_2_o6(.I0(r0_2[25:25]),.I1(r0_2[24:24]),.O(un14_s_state_df24));
defparam un14_s_state_df24_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df24_lut6_2_o5(.I0(r0_2[25:25]),.I1(r0_2[24:24]),.O(un14_s_state_lt24));
defparam un14_s_state_df24_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df22_lut6_2_o6(.I0(r0_2[23:23]),.I1(r0_2[22:22]),.O(un14_s_state_df22));
defparam un14_s_state_df22_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df22_lut6_2_o5(.I0(r0_2[23:23]),.I1(r0_2[22:22]),.O(un14_s_state_lt22));
defparam un14_s_state_df22_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df20_lut6_2_o6(.I0(r0_2[21:21]),.I1(r0_2[20:20]),.O(un14_s_state_df20));
defparam un14_s_state_df20_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df20_lut6_2_o5(.I0(r0_2[21:21]),.I1(r0_2[20:20]),.O(un14_s_state_lt20));
defparam un14_s_state_df20_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df18_lut6_2_o6(.I0(r0_2[19:19]),.I1(r0_2[18:18]),.O(un14_s_state_df18));
defparam un14_s_state_df18_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df18_lut6_2_o5(.I0(r0_2[19:19]),.I1(r0_2[18:18]),.O(un14_s_state_lt18));
defparam un14_s_state_df18_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df16_lut6_2_o6(.I0(r0_2[16:16]),.I1(r0_2[17:17]),.O(un14_s_state_df16));
defparam un14_s_state_df16_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df16_lut6_2_o5(.I0(r0_2[16:16]),.I1(r0_2[17:17]),.O(un14_s_state_lt16));
defparam un14_s_state_df16_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df14_lut6_2_o6(.I0(r0_2[14:14]),.I1(r0_2[15:15]),.O(un14_s_state_df14));
defparam un14_s_state_df14_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df14_lut6_2_o5(.I0(r0_2[14:14]),.I1(r0_2[15:15]),.O(un14_s_state_lt14));
defparam un14_s_state_df14_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df12_lut6_2_o6(.I0(r0_2[12:12]),.I1(r0_2[13:13]),.O(un14_s_state_df12));
defparam un14_s_state_df12_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df12_lut6_2_o5(.I0(r0_2[12:12]),.I1(r0_2[13:13]),.O(un14_s_state_lt12));
defparam un14_s_state_df12_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df10_lut6_2_o6(.I0(r0_2[10:10]),.I1(r0_2[11:11]),.O(un14_s_state_df10));
defparam un14_s_state_df10_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df10_lut6_2_o5(.I0(r0_2[10:10]),.I1(r0_2[11:11]),.O(un14_s_state_lt10));
defparam un14_s_state_df10_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df8_lut6_2_o6(.I0(r0_2[8:8]),.I1(r0_2[9:9]),.O(un14_s_state_df8));
defparam un14_s_state_df8_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df8_lut6_2_o5(.I0(r0_2[8:8]),.I1(r0_2[9:9]),.O(un14_s_state_lt8));
defparam un14_s_state_df8_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df6_lut6_2_o6(.I0(r0_2[6:6]),.I1(r0_2[7:7]),.O(un14_s_state_df6));
defparam un14_s_state_df6_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df6_lut6_2_o5(.I0(r0_2[6:6]),.I1(r0_2[7:7]),.O(un14_s_state_lt6));
defparam un14_s_state_df6_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df4_lut6_2_o6(.I0(r0_2[4:4]),.I1(r0_2[5:5]),.O(un14_s_state_df4));
defparam un14_s_state_df4_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df4_lut6_2_o5(.I0(r0_2[4:4]),.I1(r0_2[5:5]),.O(un14_s_state_lt4));
defparam un14_s_state_df4_lut6_2_o5.INIT=4'hE;
  LUT2 un14_s_state_df2_lut6_2_o6(.I0(r0_2[3:3]),.I1(r0_2[2:2]),.O(un14_s_state_df2));
defparam un14_s_state_df2_lut6_2_o6.INIT=4'h1;
  LUT2 un14_s_state_df2_lut6_2_o5(.I0(r0_2[3:3]),.I1(r0_2[2:2]),.O(un14_s_state_lt2));
defparam un14_s_state_df2_lut6_2_o5.INIT=4'hE;
endmodule
module post_norm_sqrt_inj (sqrt_sqr_o,pre_norm_sqrt_exp_o,s_rmode_i,post_norm_sqrt_output,s_signb_i,s_signa_i,un1_s_infa,result_4,N_6_i,un1_s_nan_a,clk_i,sqrt_ine_o,post_norm_sqrt_ine_o);
input [24:0] sqrt_sqr_o ;
input [7:0] pre_norm_sqrt_exp_o ;
input [1:0] s_rmode_i ;
output [31:0] post_norm_sqrt_output ;
input s_signb_i ;
input s_signa_i ;
input un1_s_infa ;
input result_4 ;
output N_6_i ;
input un1_s_nan_a ;
input clk_i ;
input sqrt_ine_o ;
output post_norm_sqrt_ine_o ;
wire s_signb_i ;
wire s_signa_i ;
wire un1_s_infa ;
wire result_4 ;
wire N_6_i ;
wire un1_s_nan_a ;
wire clk_i ;
wire sqrt_ine_o ;
wire post_norm_sqrt_ine_o ;
wire [22:0] s_frac_rnd ;
wire [22:22] s_output_o_0 ;
wire [22:0] s_frac_rnd_3 ;
wire [24:0] s_fract_26_i ;
wire [7:0] s_exp_i ;
wire GND ;
wire VCC ;
wire un2_s_ine_o ;
wire s_ine_i ;
wire N_959_i ;
wire s_frac_rnd_3_cry_0_cy ;
wire s_frac_rnd_3_axb_22 ;
wire s_frac_rnd_3_axb_21 ;
wire s_frac_rnd_3_axb_20 ;
wire s_frac_rnd_3_axb_19 ;
wire s_frac_rnd_3_axb_18 ;
wire s_frac_rnd_3_axb_17 ;
wire s_frac_rnd_3_axb_16 ;
wire s_frac_rnd_3_axb_15 ;
wire s_frac_rnd_3_axb_14 ;
wire s_frac_rnd_3_axb_13 ;
wire s_frac_rnd_3_axb_12 ;
wire s_frac_rnd_3_axb_11 ;
wire s_frac_rnd_3_axb_10 ;
wire s_frac_rnd_3_axb_9 ;
wire s_frac_rnd_3_axb_8 ;
wire s_frac_rnd_3_axb_7 ;
wire s_frac_rnd_3_axb_6 ;
wire s_frac_rnd_3_axb_5 ;
wire s_frac_rnd_3_axb_4 ;
wire s_frac_rnd_3_axb_3 ;
wire s_frac_rnd_3_axb_2 ;
wire s_frac_rnd_3_axb_1 ;
wire s_frac_rnd_3_axb_0 ;
wire N_959_1 ;
wire s_frac_rnd_3_cry_21 ;
wire s_frac_rnd_3_cry_20 ;
wire s_frac_rnd_3_cry_19 ;
wire s_frac_rnd_3_cry_18 ;
wire s_frac_rnd_3_cry_17 ;
wire s_frac_rnd_3_cry_16 ;
wire s_frac_rnd_3_cry_15 ;
wire s_frac_rnd_3_cry_14 ;
wire s_frac_rnd_3_cry_13 ;
wire s_frac_rnd_3_cry_12 ;
wire s_frac_rnd_3_cry_11 ;
wire s_frac_rnd_3_cry_10 ;
wire s_frac_rnd_3_cry_9 ;
wire s_frac_rnd_3_cry_8 ;
wire s_frac_rnd_3_cry_7 ;
wire s_frac_rnd_3_cry_6 ;
wire s_frac_rnd_3_cry_5 ;
wire s_frac_rnd_3_cry_4 ;
wire s_frac_rnd_3_cry_3 ;
wire s_frac_rnd_3_cry_2 ;
wire s_frac_rnd_3_cry_1 ;
wire s_frac_rnd_3_cry_0 ;
// instances
  LUT5 desc3261(.I0(s_signa_i),.I1(result_4),.I2(un1_s_infa),.I3(un1_s_nan_a),.I4(s_frac_rnd[22:22]),.O(s_output_o_0[22:22]));
defparam desc3261.INIT=32'hFF8FFF88;
  FD desc3262(.Q(s_frac_rnd[18:18]),.D(s_frac_rnd_3[18:18]),.C(clk_i));
  FD desc3263(.Q(s_frac_rnd[19:19]),.D(s_frac_rnd_3[19:19]),.C(clk_i));
  FD desc3264(.Q(s_frac_rnd[20:20]),.D(s_frac_rnd_3[20:20]),.C(clk_i));
  FD desc3265(.Q(s_frac_rnd[21:21]),.D(s_frac_rnd_3[21:21]),.C(clk_i));
  FD desc3266(.Q(s_frac_rnd[22:22]),.D(s_frac_rnd_3[22:22]),.C(clk_i));
  FD desc3267(.Q(s_frac_rnd[3:3]),.D(s_frac_rnd_3[3:3]),.C(clk_i));
  FD desc3268(.Q(s_frac_rnd[4:4]),.D(s_frac_rnd_3[4:4]),.C(clk_i));
  FD desc3269(.Q(s_frac_rnd[5:5]),.D(s_frac_rnd_3[5:5]),.C(clk_i));
  FD desc3270(.Q(s_frac_rnd[6:6]),.D(s_frac_rnd_3[6:6]),.C(clk_i));
  FD desc3271(.Q(s_frac_rnd[7:7]),.D(s_frac_rnd_3[7:7]),.C(clk_i));
  FD desc3272(.Q(s_frac_rnd[8:8]),.D(s_frac_rnd_3[8:8]),.C(clk_i));
  FD desc3273(.Q(s_frac_rnd[9:9]),.D(s_frac_rnd_3[9:9]),.C(clk_i));
  FD desc3274(.Q(s_frac_rnd[10:10]),.D(s_frac_rnd_3[10:10]),.C(clk_i));
  FD desc3275(.Q(s_frac_rnd[11:11]),.D(s_frac_rnd_3[11:11]),.C(clk_i));
  FD desc3276(.Q(s_frac_rnd[12:12]),.D(s_frac_rnd_3[12:12]),.C(clk_i));
  FD desc3277(.Q(s_frac_rnd[13:13]),.D(s_frac_rnd_3[13:13]),.C(clk_i));
  FD desc3278(.Q(s_frac_rnd[14:14]),.D(s_frac_rnd_3[14:14]),.C(clk_i));
  FD desc3279(.Q(s_frac_rnd[15:15]),.D(s_frac_rnd_3[15:15]),.C(clk_i));
  FD desc3280(.Q(s_frac_rnd[16:16]),.D(s_frac_rnd_3[16:16]),.C(clk_i));
  FD desc3281(.Q(s_frac_rnd[17:17]),.D(s_frac_rnd_3[17:17]),.C(clk_i));
  FD desc3282(.Q(s_frac_rnd[0:0]),.D(s_frac_rnd_3[0:0]),.C(clk_i));
  FD desc3283(.Q(s_frac_rnd[1:1]),.D(s_frac_rnd_3[1:1]),.C(clk_i));
  FD desc3284(.Q(s_frac_rnd[2:2]),.D(s_frac_rnd_3[2:2]),.C(clk_i));
  FD desc3285(.Q(s_fract_26_i[14:14]),.D(sqrt_sqr_o[14:14]),.C(clk_i));
  FD desc3286(.Q(s_fract_26_i[15:15]),.D(sqrt_sqr_o[15:15]),.C(clk_i));
  FD desc3287(.Q(s_fract_26_i[16:16]),.D(sqrt_sqr_o[16:16]),.C(clk_i));
  FD desc3288(.Q(s_fract_26_i[17:17]),.D(sqrt_sqr_o[17:17]),.C(clk_i));
  FD desc3289(.Q(s_fract_26_i[18:18]),.D(sqrt_sqr_o[18:18]),.C(clk_i));
  FD desc3290(.Q(s_fract_26_i[19:19]),.D(sqrt_sqr_o[19:19]),.C(clk_i));
  FD desc3291(.Q(s_fract_26_i[20:20]),.D(sqrt_sqr_o[20:20]),.C(clk_i));
  FD desc3292(.Q(s_fract_26_i[21:21]),.D(sqrt_sqr_o[21:21]),.C(clk_i));
  FD desc3293(.Q(s_fract_26_i[22:22]),.D(sqrt_sqr_o[22:22]),.C(clk_i));
  FD desc3294(.Q(s_fract_26_i[23:23]),.D(sqrt_sqr_o[23:23]),.C(clk_i));
  FD desc3295(.Q(s_fract_26_i[24:24]),.D(sqrt_sqr_o[24:24]),.C(clk_i));
  FD desc3296(.Q(s_exp_i[7:7]),.D(pre_norm_sqrt_exp_o[7:7]),.C(clk_i));
  FD desc3297(.Q(s_fract_26_i[0:0]),.D(sqrt_sqr_o[0:0]),.C(clk_i));
  FD desc3298(.Q(s_fract_26_i[1:1]),.D(sqrt_sqr_o[1:1]),.C(clk_i));
  FD desc3299(.Q(s_fract_26_i[2:2]),.D(sqrt_sqr_o[2:2]),.C(clk_i));
  FD desc3300(.Q(s_fract_26_i[3:3]),.D(sqrt_sqr_o[3:3]),.C(clk_i));
  FD desc3301(.Q(s_fract_26_i[4:4]),.D(sqrt_sqr_o[4:4]),.C(clk_i));
  FD desc3302(.Q(s_fract_26_i[5:5]),.D(sqrt_sqr_o[5:5]),.C(clk_i));
  FD desc3303(.Q(s_fract_26_i[6:6]),.D(sqrt_sqr_o[6:6]),.C(clk_i));
  FD desc3304(.Q(s_fract_26_i[7:7]),.D(sqrt_sqr_o[7:7]),.C(clk_i));
  FD desc3305(.Q(s_fract_26_i[8:8]),.D(sqrt_sqr_o[8:8]),.C(clk_i));
  FD desc3306(.Q(s_fract_26_i[9:9]),.D(sqrt_sqr_o[9:9]),.C(clk_i));
  FD desc3307(.Q(s_fract_26_i[10:10]),.D(sqrt_sqr_o[10:10]),.C(clk_i));
  FD desc3308(.Q(s_fract_26_i[11:11]),.D(sqrt_sqr_o[11:11]),.C(clk_i));
  FD desc3309(.Q(s_fract_26_i[12:12]),.D(sqrt_sqr_o[12:12]),.C(clk_i));
  FD desc3310(.Q(s_fract_26_i[13:13]),.D(sqrt_sqr_o[13:13]),.C(clk_i));
  FD desc3311(.Q(post_norm_sqrt_output[31:31]),.D(s_signa_i),.C(clk_i));
  FD desc3312(.Q(s_exp_i[0:0]),.D(pre_norm_sqrt_exp_o[0:0]),.C(clk_i));
  FD desc3313(.Q(s_exp_i[1:1]),.D(pre_norm_sqrt_exp_o[1:1]),.C(clk_i));
  FD desc3314(.Q(s_exp_i[2:2]),.D(pre_norm_sqrt_exp_o[2:2]),.C(clk_i));
  FD desc3315(.Q(s_exp_i[3:3]),.D(pre_norm_sqrt_exp_o[3:3]),.C(clk_i));
  FD desc3316(.Q(s_exp_i[4:4]),.D(pre_norm_sqrt_exp_o[4:4]),.C(clk_i));
  FD desc3317(.Q(s_exp_i[5:5]),.D(pre_norm_sqrt_exp_o[5:5]),.C(clk_i));
  FD desc3318(.Q(s_exp_i[6:6]),.D(pre_norm_sqrt_exp_o[6:6]),.C(clk_i));
  FD desc3319(.Q(post_norm_sqrt_output[22:22]),.D(s_output_o_0[22:22]),.C(clk_i));
  FD s_ine_i_Z(.Q(s_ine_i),.D(sqrt_ine_o),.C(clk_i));
  FDR desc3320(.Q(post_norm_sqrt_output[11:11]),.D(s_frac_rnd[11:11]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3321(.Q(post_norm_sqrt_output[12:12]),.D(s_frac_rnd[12:12]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3322(.Q(post_norm_sqrt_output[13:13]),.D(s_frac_rnd[13:13]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3323(.Q(post_norm_sqrt_output[14:14]),.D(s_frac_rnd[14:14]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3324(.Q(post_norm_sqrt_output[15:15]),.D(s_frac_rnd[15:15]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3325(.Q(post_norm_sqrt_output[16:16]),.D(s_frac_rnd[16:16]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3326(.Q(post_norm_sqrt_output[17:17]),.D(s_frac_rnd[17:17]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3327(.Q(post_norm_sqrt_output[18:18]),.D(s_frac_rnd[18:18]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3328(.Q(post_norm_sqrt_output[19:19]),.D(s_frac_rnd[19:19]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3329(.Q(post_norm_sqrt_output[20:20]),.D(s_frac_rnd[20:20]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3330(.Q(post_norm_sqrt_output[21:21]),.D(s_frac_rnd[21:21]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3331(.Q(post_norm_sqrt_output[0:0]),.D(s_frac_rnd[0:0]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3332(.Q(post_norm_sqrt_output[1:1]),.D(s_frac_rnd[1:1]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3333(.Q(post_norm_sqrt_output[2:2]),.D(s_frac_rnd[2:2]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3334(.Q(post_norm_sqrt_output[3:3]),.D(s_frac_rnd[3:3]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3335(.Q(post_norm_sqrt_output[4:4]),.D(s_frac_rnd[4:4]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3336(.Q(post_norm_sqrt_output[5:5]),.D(s_frac_rnd[5:5]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3337(.Q(post_norm_sqrt_output[6:6]),.D(s_frac_rnd[6:6]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3338(.Q(post_norm_sqrt_output[7:7]),.D(s_frac_rnd[7:7]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3339(.Q(post_norm_sqrt_output[8:8]),.D(s_frac_rnd[8:8]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3340(.Q(post_norm_sqrt_output[9:9]),.D(s_frac_rnd[9:9]),.C(clk_i),.R(un2_s_ine_o));
  FDR desc3341(.Q(post_norm_sqrt_output[10:10]),.D(s_frac_rnd[10:10]),.C(clk_i),.R(un2_s_ine_o));
  FDR ine_o_Z(.Q(post_norm_sqrt_ine_o),.D(s_ine_i),.C(clk_i),.R(un2_s_ine_o));
  MUXCY_L s_frac_rnd_3_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(N_959_i),.LO(s_frac_rnd_3_cry_0_cy));
  LUT1_L s_frac_rnd_3_axb_22_cZ(.I0(s_fract_26_i[24:24]),.LO(s_frac_rnd_3_axb_22));
defparam s_frac_rnd_3_axb_22_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_21_cZ(.I0(s_fract_26_i[23:23]),.LO(s_frac_rnd_3_axb_21));
defparam s_frac_rnd_3_axb_21_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_20_cZ(.I0(s_fract_26_i[22:22]),.LO(s_frac_rnd_3_axb_20));
defparam s_frac_rnd_3_axb_20_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_19_cZ(.I0(s_fract_26_i[21:21]),.LO(s_frac_rnd_3_axb_19));
defparam s_frac_rnd_3_axb_19_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_18_cZ(.I0(s_fract_26_i[20:20]),.LO(s_frac_rnd_3_axb_18));
defparam s_frac_rnd_3_axb_18_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_17_cZ(.I0(s_fract_26_i[19:19]),.LO(s_frac_rnd_3_axb_17));
defparam s_frac_rnd_3_axb_17_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_16_cZ(.I0(s_fract_26_i[18:18]),.LO(s_frac_rnd_3_axb_16));
defparam s_frac_rnd_3_axb_16_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_15_cZ(.I0(s_fract_26_i[17:17]),.LO(s_frac_rnd_3_axb_15));
defparam s_frac_rnd_3_axb_15_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_14_cZ(.I0(s_fract_26_i[16:16]),.LO(s_frac_rnd_3_axb_14));
defparam s_frac_rnd_3_axb_14_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_13_cZ(.I0(s_fract_26_i[15:15]),.LO(s_frac_rnd_3_axb_13));
defparam s_frac_rnd_3_axb_13_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_12_cZ(.I0(s_fract_26_i[14:14]),.LO(s_frac_rnd_3_axb_12));
defparam s_frac_rnd_3_axb_12_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_11_cZ(.I0(s_fract_26_i[13:13]),.LO(s_frac_rnd_3_axb_11));
defparam s_frac_rnd_3_axb_11_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_10_cZ(.I0(s_fract_26_i[12:12]),.LO(s_frac_rnd_3_axb_10));
defparam s_frac_rnd_3_axb_10_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_9_cZ(.I0(s_fract_26_i[11:11]),.LO(s_frac_rnd_3_axb_9));
defparam s_frac_rnd_3_axb_9_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_8_cZ(.I0(s_fract_26_i[10:10]),.LO(s_frac_rnd_3_axb_8));
defparam s_frac_rnd_3_axb_8_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_7_cZ(.I0(s_fract_26_i[9:9]),.LO(s_frac_rnd_3_axb_7));
defparam s_frac_rnd_3_axb_7_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_6_cZ(.I0(s_fract_26_i[8:8]),.LO(s_frac_rnd_3_axb_6));
defparam s_frac_rnd_3_axb_6_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_5_cZ(.I0(s_fract_26_i[7:7]),.LO(s_frac_rnd_3_axb_5));
defparam s_frac_rnd_3_axb_5_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_4_cZ(.I0(s_fract_26_i[6:6]),.LO(s_frac_rnd_3_axb_4));
defparam s_frac_rnd_3_axb_4_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_3_cZ(.I0(s_fract_26_i[5:5]),.LO(s_frac_rnd_3_axb_3));
defparam s_frac_rnd_3_axb_3_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_2_cZ(.I0(s_fract_26_i[4:4]),.LO(s_frac_rnd_3_axb_2));
defparam s_frac_rnd_3_axb_2_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_1_cZ(.I0(s_fract_26_i[3:3]),.LO(s_frac_rnd_3_axb_1));
defparam s_frac_rnd_3_axb_1_cZ.INIT=2'h2;
  LUT1_L s_frac_rnd_3_axb_0_cZ(.I0(s_fract_26_i[2:2]),.LO(s_frac_rnd_3_axb_0));
defparam s_frac_rnd_3_axb_0_cZ.INIT=2'h2;
  LUT5_L s_roundup_3_i_1(.I0(s_fract_26_i[0:0]),.I1(s_fract_26_i[1:1]),.I2(s_fract_26_i[3:3]),.I3(s_ine_i),.I4(s_rmode_i[1:1]),.LO(N_959_1));
defparam s_roundup_3_i_1.INIT=32'h00110015;
  LUT5 s_frac_rnd_3_cry_0_cy_RNO(.I0(s_fract_26_i[1:1]),.I1(s_rmode_i[0:0]),.I2(s_rmode_i[1:1]),.I3(s_signa_i),.I4(N_959_1),.O(N_959_i));
defparam s_frac_rnd_3_cry_0_cy_RNO.INIT=32'h0000C232;
  XORCY s_frac_rnd_3_s_22(.LI(s_frac_rnd_3_axb_22),.CI(s_frac_rnd_3_cry_21),.O(s_frac_rnd_3[22:22]));
  XORCY s_frac_rnd_3_s_21(.LI(s_frac_rnd_3_axb_21),.CI(s_frac_rnd_3_cry_20),.O(s_frac_rnd_3[21:21]));
  MUXCY_L s_frac_rnd_3_cry_21_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_20),.S(s_frac_rnd_3_axb_21),.LO(s_frac_rnd_3_cry_21));
  XORCY s_frac_rnd_3_s_20(.LI(s_frac_rnd_3_axb_20),.CI(s_frac_rnd_3_cry_19),.O(s_frac_rnd_3[20:20]));
  MUXCY_L s_frac_rnd_3_cry_20_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_19),.S(s_frac_rnd_3_axb_20),.LO(s_frac_rnd_3_cry_20));
  XORCY s_frac_rnd_3_s_19(.LI(s_frac_rnd_3_axb_19),.CI(s_frac_rnd_3_cry_18),.O(s_frac_rnd_3[19:19]));
  MUXCY_L s_frac_rnd_3_cry_19_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_18),.S(s_frac_rnd_3_axb_19),.LO(s_frac_rnd_3_cry_19));
  XORCY s_frac_rnd_3_s_18(.LI(s_frac_rnd_3_axb_18),.CI(s_frac_rnd_3_cry_17),.O(s_frac_rnd_3[18:18]));
  MUXCY_L s_frac_rnd_3_cry_18_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_17),.S(s_frac_rnd_3_axb_18),.LO(s_frac_rnd_3_cry_18));
  XORCY s_frac_rnd_3_s_17(.LI(s_frac_rnd_3_axb_17),.CI(s_frac_rnd_3_cry_16),.O(s_frac_rnd_3[17:17]));
  MUXCY_L s_frac_rnd_3_cry_17_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_16),.S(s_frac_rnd_3_axb_17),.LO(s_frac_rnd_3_cry_17));
  XORCY s_frac_rnd_3_s_16(.LI(s_frac_rnd_3_axb_16),.CI(s_frac_rnd_3_cry_15),.O(s_frac_rnd_3[16:16]));
  MUXCY_L s_frac_rnd_3_cry_16_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_15),.S(s_frac_rnd_3_axb_16),.LO(s_frac_rnd_3_cry_16));
  XORCY s_frac_rnd_3_s_15(.LI(s_frac_rnd_3_axb_15),.CI(s_frac_rnd_3_cry_14),.O(s_frac_rnd_3[15:15]));
  MUXCY_L s_frac_rnd_3_cry_15_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_14),.S(s_frac_rnd_3_axb_15),.LO(s_frac_rnd_3_cry_15));
  XORCY s_frac_rnd_3_s_14(.LI(s_frac_rnd_3_axb_14),.CI(s_frac_rnd_3_cry_13),.O(s_frac_rnd_3[14:14]));
  MUXCY_L s_frac_rnd_3_cry_14_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_13),.S(s_frac_rnd_3_axb_14),.LO(s_frac_rnd_3_cry_14));
  XORCY s_frac_rnd_3_s_13(.LI(s_frac_rnd_3_axb_13),.CI(s_frac_rnd_3_cry_12),.O(s_frac_rnd_3[13:13]));
  MUXCY_L s_frac_rnd_3_cry_13_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_12),.S(s_frac_rnd_3_axb_13),.LO(s_frac_rnd_3_cry_13));
  XORCY s_frac_rnd_3_s_12(.LI(s_frac_rnd_3_axb_12),.CI(s_frac_rnd_3_cry_11),.O(s_frac_rnd_3[12:12]));
  MUXCY_L s_frac_rnd_3_cry_12_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_11),.S(s_frac_rnd_3_axb_12),.LO(s_frac_rnd_3_cry_12));
  XORCY s_frac_rnd_3_s_11(.LI(s_frac_rnd_3_axb_11),.CI(s_frac_rnd_3_cry_10),.O(s_frac_rnd_3[11:11]));
  MUXCY_L s_frac_rnd_3_cry_11_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_10),.S(s_frac_rnd_3_axb_11),.LO(s_frac_rnd_3_cry_11));
  XORCY s_frac_rnd_3_s_10(.LI(s_frac_rnd_3_axb_10),.CI(s_frac_rnd_3_cry_9),.O(s_frac_rnd_3[10:10]));
  MUXCY_L s_frac_rnd_3_cry_10_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_9),.S(s_frac_rnd_3_axb_10),.LO(s_frac_rnd_3_cry_10));
  XORCY s_frac_rnd_3_s_9(.LI(s_frac_rnd_3_axb_9),.CI(s_frac_rnd_3_cry_8),.O(s_frac_rnd_3[9:9]));
  MUXCY_L s_frac_rnd_3_cry_9_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_8),.S(s_frac_rnd_3_axb_9),.LO(s_frac_rnd_3_cry_9));
  XORCY s_frac_rnd_3_s_8(.LI(s_frac_rnd_3_axb_8),.CI(s_frac_rnd_3_cry_7),.O(s_frac_rnd_3[8:8]));
  MUXCY_L s_frac_rnd_3_cry_8_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_7),.S(s_frac_rnd_3_axb_8),.LO(s_frac_rnd_3_cry_8));
  XORCY s_frac_rnd_3_s_7(.LI(s_frac_rnd_3_axb_7),.CI(s_frac_rnd_3_cry_6),.O(s_frac_rnd_3[7:7]));
  MUXCY_L s_frac_rnd_3_cry_7_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_6),.S(s_frac_rnd_3_axb_7),.LO(s_frac_rnd_3_cry_7));
  XORCY s_frac_rnd_3_s_6(.LI(s_frac_rnd_3_axb_6),.CI(s_frac_rnd_3_cry_5),.O(s_frac_rnd_3[6:6]));
  MUXCY_L s_frac_rnd_3_cry_6_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_5),.S(s_frac_rnd_3_axb_6),.LO(s_frac_rnd_3_cry_6));
  XORCY s_frac_rnd_3_s_5(.LI(s_frac_rnd_3_axb_5),.CI(s_frac_rnd_3_cry_4),.O(s_frac_rnd_3[5:5]));
  MUXCY_L s_frac_rnd_3_cry_5_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_4),.S(s_frac_rnd_3_axb_5),.LO(s_frac_rnd_3_cry_5));
  XORCY s_frac_rnd_3_s_4(.LI(s_frac_rnd_3_axb_4),.CI(s_frac_rnd_3_cry_3),.O(s_frac_rnd_3[4:4]));
  MUXCY_L s_frac_rnd_3_cry_4_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_3),.S(s_frac_rnd_3_axb_4),.LO(s_frac_rnd_3_cry_4));
  XORCY s_frac_rnd_3_s_3(.LI(s_frac_rnd_3_axb_3),.CI(s_frac_rnd_3_cry_2),.O(s_frac_rnd_3[3:3]));
  MUXCY_L s_frac_rnd_3_cry_3_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_2),.S(s_frac_rnd_3_axb_3),.LO(s_frac_rnd_3_cry_3));
  XORCY s_frac_rnd_3_s_2(.LI(s_frac_rnd_3_axb_2),.CI(s_frac_rnd_3_cry_1),.O(s_frac_rnd_3[2:2]));
  MUXCY_L s_frac_rnd_3_cry_2_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_1),.S(s_frac_rnd_3_axb_2),.LO(s_frac_rnd_3_cry_2));
  XORCY s_frac_rnd_3_s_1(.LI(s_frac_rnd_3_axb_1),.CI(s_frac_rnd_3_cry_0),.O(s_frac_rnd_3[1:1]));
  MUXCY_L s_frac_rnd_3_cry_1_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_0),.S(s_frac_rnd_3_axb_1),.LO(s_frac_rnd_3_cry_1));
  XORCY s_frac_rnd_3_s_0(.LI(s_frac_rnd_3_axb_0),.CI(s_frac_rnd_3_cry_0_cy),.O(s_frac_rnd_3[0:0]));
  MUXCY_L s_frac_rnd_3_cry_0_cZ(.DI(GND),.CI(s_frac_rnd_3_cry_0_cy),.S(s_frac_rnd_3_axb_0),.LO(s_frac_rnd_3_cry_0));
  FDS desc3342(.Q(post_norm_sqrt_output[26:26]),.D(s_exp_i[3:3]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3343(.Q(post_norm_sqrt_output[27:27]),.D(s_exp_i[4:4]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3344(.Q(post_norm_sqrt_output[28:28]),.D(s_exp_i[5:5]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3345(.Q(post_norm_sqrt_output[29:29]),.D(s_exp_i[6:6]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3346(.Q(post_norm_sqrt_output[30:30]),.D(s_exp_i[7:7]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3347(.Q(post_norm_sqrt_output[23:23]),.D(s_exp_i[0:0]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3348(.Q(post_norm_sqrt_output[24:24]),.D(s_exp_i[1:1]),.C(clk_i),.S(un2_s_ine_o));
  FDS desc3349(.Q(post_norm_sqrt_output[25:25]),.D(s_exp_i[2:2]),.C(clk_i),.S(un2_s_ine_o));
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  LUT3 un2_s_ine_o_lut6_2_o6(.I0(s_signa_i),.I1(un1_s_infa),.I2(result_4),.O(un2_s_ine_o));
defparam un2_s_ine_o_lut6_2_o6.INIT=8'hEC;
  LUT2 un2_s_ine_o_lut6_2_o5(.I0(s_signb_i),.I1(s_signa_i),.O(N_6_i));
defparam un2_s_ine_o_lut6_2_o5.INIT=4'h6;
endmodule
module fpu_inj (clk_i,opa_i,opb_i,fpu_op_i,rmode_i,output_o,start_i,ready_o,ine_o,overflow_o,underflow_o,div_zero_o,inf_o,zero_o,qnan_o,snan_o,p_desc595_p_O_FDpre_norm_mul_,p_desc596_p_O_FDpre_norm_mul_,p_desc597_p_O_FDpre_norm_mul_,p_desc598_p_O_FDpre_norm_mul_,p_desc599_p_O_FDpre_norm_mul_,p_desc600_p_O_FDpre_norm_mul_,p_desc601_p_O_FDpre_norm_mul_,p_desc602_p_O_FDpre_norm_mul_,p_desc603_p_O_FDpre_norm_mul_,p_desc604_p_O_FDpre_norm_mul_,p_desc1070_p_O_FDpost_norm_mul_,p_desc1071_p_O_FDpost_norm_mul_,p_desc1072_p_O_FDpost_norm_mul_,p_desc1073_p_O_FDpost_norm_mul_,p_desc1074_p_O_FDpost_norm_mul_,p_desc1075_p_O_FDpost_norm_mul_,p_desc1076_p_O_FDpost_norm_mul_,p_desc1077_p_O_FDpost_norm_mul_,p_desc1078_p_O_FDpost_norm_mul_,p_desc1079_p_O_FDpost_norm_mul_,p_desc1080_p_O_FDpost_norm_mul_,p_desc1081_p_O_FDpost_norm_mul_,p_desc1082_p_O_FDpost_norm_mul_,p_desc1083_p_O_FDpost_norm_mul_,p_desc1084_p_O_FDpost_norm_mul_,p_desc1085_p_O_FDpost_norm_mul_,p_desc1086_p_O_FDpost_norm_mul_,p_desc1087_p_O_FDpost_norm_mul_,p_desc1088_p_O_FDpost_norm_mul_,p_desc1089_p_O_FDpost_norm_mul_,p_desc1090_p_O_FDpost_norm_mul_,p_desc1091_p_O_FDpost_norm_mul_,p_desc1092_p_O_FDpost_norm_mul_,p_desc1163_p_O_FDpost_norm_mul_,p_desc1164_p_O_FDpost_norm_mul_,p_desc1165_p_O_FDpost_norm_mul_,p_desc1166_p_O_FDpost_norm_mul_,p_desc1167_p_O_FDpost_norm_mul_,p_desc1168_p_O_FDpost_norm_mul_,p_desc1169_p_O_FDpost_norm_mul_,p_desc1170_p_O_FDpost_norm_mul_,p_desc1171_p_O_FDpost_norm_mul_,p_desc1172_p_O_FDpost_norm_mul_,p_desc1173_p_O_FDpost_norm_mul_,p_desc1174_p_O_FDpost_norm_mul_,p_desc1175_p_O_FDpost_norm_mul_,p_desc1176_p_O_FDpost_norm_mul_,p_desc1177_p_O_FDpost_norm_mul_,p_desc1178_p_O_FDpost_norm_mul_,p_desc1179_p_O_FDpost_norm_mul_,p_desc1180_p_O_FDpost_norm_mul_,p_desc1181_p_O_FDpost_norm_mul_,p_desc1182_p_O_FDpost_norm_mul_,p_desc1183_p_O_FDpost_norm_mul_,p_desc1184_p_O_FDpost_norm_mul_,p_desc1185_p_O_FDpost_norm_mul_,p_desc1186_p_O_FDpost_norm_mul_,p_desc1187_p_O_FDpost_norm_mul_,p_desc1188_p_O_FDpost_norm_mul_,p_desc1189_p_O_FDpost_norm_mul_,p_desc1190_p_O_FDpost_norm_mul_,p_desc1191_p_O_FDpost_norm_mul_,p_desc1192_p_O_FDpost_norm_mul_,p_desc1193_p_O_FDpost_norm_mul_,p_desc1194_p_O_FDpost_norm_mul_,p_desc1195_p_O_FDpost_norm_mul_,p_desc1196_p_O_FDpost_norm_mul_,p_desc1197_p_O_FDpost_norm_mul_,p_desc1198_p_O_FDpost_norm_mul_,p_desc1199_p_O_FDpost_norm_mul_,p_desc1200_p_O_FDpost_norm_mul_,p_desc1201_p_O_FDpost_norm_mul_,p_desc1202_p_O_FDpost_norm_mul_,p_desc1203_p_O_FDpost_norm_mul_,p_desc1204_p_O_FDpost_norm_mul_,p_desc1205_p_O_FDpost_norm_mul_,p_desc1206_p_O_FDpost_norm_mul_,p_desc1207_p_O_FDpost_norm_mul_,p_desc1208_p_O_FDpost_norm_mul_,p_desc1209_p_O_FDpost_norm_mul_,p_desc1210_p_O_FDpost_norm_mul_,p_desc1211_p_O_FDpost_norm_mul_,p_desc1212_p_O_FDpost_norm_mul_,p_desc1213_p_O_FDpost_norm_mul_,p_desc1214_p_O_FDpost_norm_mul_,p_desc1215_p_O_FDpost_norm_mul_,p_desc1216_p_O_FDpost_norm_mul_,p_desc1217_p_O_FDpost_norm_mul_,p_desc1218_p_O_FDpost_norm_mul_,p_desc1219_p_O_FDpost_norm_mul_,p_desc1220_p_O_FDpost_norm_mul_,p_desc1221_p_O_FDpost_norm_mul_,p_s_sign_i_Z_p_O_FDpost_norm_mul_,p_ine_o_Z_p_O_FDpost_norm_mul_,p_desc1244_p_O_FDpost_norm_mul_,p_desc1245_p_O_FDpost_norm_mul_,p_desc1246_p_O_FDpost_norm_mul_,p_desc1247_p_O_FDpost_norm_mul_,p_desc1248_p_O_FDpost_norm_mul_,p_desc1249_p_O_FDpost_norm_mul_,p_desc1250_p_O_FDpost_norm_mul_,p_desc1251_p_O_FDpost_norm_mul_,p_desc1252_p_O_FDpost_norm_mul_,p_desc1253_p_O_FDpost_norm_mul_,p_desc1254_p_O_FDpost_norm_mul_,p_desc1255_p_O_FDpost_norm_mul_,p_desc1256_p_O_FDpost_norm_mul_,p_desc1257_p_O_FDpost_norm_mul_,p_desc1258_p_O_FDpost_norm_mul_,p_desc1259_p_O_FDpost_norm_mul_,p_desc1260_p_O_FDpost_norm_mul_,p_desc1261_p_O_FDpost_norm_mul_,p_desc1262_p_O_FDpost_norm_mul_,p_desc1263_p_O_FDpost_norm_mul_,p_desc1264_p_O_FDpost_norm_mul_,p_desc1265_p_O_FDpost_norm_mul_,p_desc1266_p_O_FDpost_norm_mul_,p_desc1267_p_O_FDpost_norm_mul_,p_desc1268_p_O_FDpost_norm_mul_,p_desc1269_p_O_FDpost_norm_mul_,p_desc1270_p_O_FDpost_norm_mul_,p_desc1271_p_O_FDpost_norm_mul_,p_desc1272_p_O_FDpost_norm_mul_,p_desc1273_p_O_FDpost_norm_mul_,p_desc1274_p_O_FDpost_norm_mul_,p_desc1275_p_O_FDpost_norm_mul_,p_desc1276_p_O_FDpost_norm_mul_,p_desc1277_p_O_FDpost_norm_mul_,p_desc1278_p_O_FDpost_norm_mul_,p_desc1279_p_O_FDpost_norm_mul_,p_desc1280_p_O_FDpost_norm_mul_,p_desc1281_p_O_FDpost_norm_mul_,p_desc1282_p_O_FDpost_norm_mul_,p_desc1283_p_O_FDpost_norm_mul_,p_desc1284_p_O_FDpost_norm_mul_,p_desc1285_p_O_FDpost_norm_mul_,p_desc1286_p_O_FDpost_norm_mul_,p_desc1287_p_O_FDpost_norm_mul_,p_desc1288_p_O_FDpost_norm_mul_,p_desc1289_p_O_FDpost_norm_mul_,p_desc1290_p_O_FDpost_norm_mul_,p_desc1291_p_O_FDpost_norm_mul_);
input clk_i ;
input [31:0] opa_i ;
input [31:0] opb_i ;
input [2:0] fpu_op_i ;
input [1:0] rmode_i ;
output [31:0] output_o ;
input start_i ;
output ready_o ;
output ine_o ;
output overflow_o ;
output underflow_o ;
output div_zero_o ;
output inf_o ;
output zero_o ;
output qnan_o ;
output snan_o ;
wire clk_i ;
wire start_i ;
wire ready_o ;
wire ine_o ;
wire overflow_o ;
wire underflow_o ;
wire div_zero_o ;
wire inf_o ;
wire zero_o ;
wire qnan_o ;
wire snan_o ;
wire [31:0] s_opa_i ;
wire [31:0] s_opb_i ;
wire [26:0] prenorm_addsub_fracta_28_o ;
wire [26:0] prenorm_addsub_fractb_28_o ;
wire [7:0] prenorm_addsub_exp_o ;
wire [2:0] s_fpu_op_i ;
wire [27:0] addsub_fract_o ;
wire [1:0] s_rmode_i ;
wire [31:0] postnorm_addsub_output_o ;
wire [9:0] pre_norm_mul_exp_10 ;
wire [31:0] post_norm_mul_output ;
wire [48:34] pre_norm_div_dvdnd ;
wire [22:5] pre_norm_div_dvsor ;
wire [26:0] serial_div_qutnt ;
wire [26:0] serial_div_rmndr ;
wire [31:0] post_norm_div_output ;
wire [50:27] pre_norm_sqrt_fracta_o ;
wire [7:0] pre_norm_sqrt_exp_o ;
wire [24:0] sqrt_sqr_o ;
wire [31:0] post_norm_sqrt_output ;
wire [31:0] s_count ;
wire [31:0] s_output1 ;
wire s_state ;
wire [23:23] s_output_o ;
wire [4:0] \i_pre_norm_sqrt.v_count  ;
wire [1:0] \i_post_norm_mul.s_rmode_i  ;
wire [30:24] \i_post_norm_mul.s_opa_i  ;
wire [30:24] \i_post_norm_mul.s_opb_i  ;
wire \i_serial_div.s_state  ;
wire [22:0] \i_mul_24.s_fracta_i  ;
wire [22:0] \i_mul_24.s_fractb_i  ;
wire s_count_RNIS5BE1 ;
wire s_count_RNIME821 ;
wire [21:21] s_count_RNIM79LF ;
wire [7:6] s_output1_6_2_i_m2 ;
wire [4:4] \i_pre_norm_div.v_count_2_0  ;
wire [47:0] mul_24_fract_48 ;
wire [1:0] \i_pre_norm_mul.s_exp_10_o_0  ;
wire [1:0] \i_pre_norm_mul.s_exp_10_o  ;
wire [9:1] \i_pre_norm_div.un11_s_exp_10_o_0  ;
wire \i_pre_norm_div.v_count_1_0_2  ;
wire [1:1] \i_pre_norm_div.v_count_1_0_0_a2_0  ;
wire [29:28] s_opa_i_i ;
wire \i_pre_norm_sqrt.v_count_i  ;
wire [4:4] \i_prenorm_addsub.v_count_56_0_2  ;
wire \i_pre_norm_div.v_count_1_0_a2_7_i_0  ;
wire \i_pre_norm_div.v_count_1_0_1  ;
wire [51:51] pre_norm_sqrt_fracta_o_0 ;
wire [31:22] s_output_o_0 ;
wire [49:49] pre_norm_div_dvdnd_0 ;
wire [23:23] pre_norm_div_dvsor_0 ;
wire [33:29] \i_pre_norm_sqrt.s_fracta_52_o_0_e  ;
wire addsub_sign_o ;
wire postnorm_addsub_ine_o ;
wire post_norm_mul_ine ;
wire post_norm_div_ine ;
wire sqrt_ine_o ;
wire post_norm_sqrt_ine_o ;
wire VCC ;
wire GND ;
wire s_ine_o ;
wire un3_s_snan_o_0 ;
wire \i_sqrt.s_start_i  ;
wire \i_post_norm_mul.or_reduce.result_5  ;
wire un12_s_state_0_a2_lut6_2_O5 ;
wire \i_mul_24.s_signa_i  ;
wire \i_mul_24.s_signb_i  ;
wire \i_prenorm_addsub.s_expa_lt_expb  ;
wire N_6_i ;
wire \or_reduce.result_1_i_o3  ;
wire \or_reduce.result_i_o3_lut6_2_O6  ;
wire un4_s_expb_in_2_i_o2_2_lut6_2_O5 ;
wire \i_post_norm_mul.un3_s_op_0  ;
wire div_zero_o_0 ;
wire i155_mux ;
wire un1_s_count_4_cry_0_cy_RNO ;
wire s_ine_o_5 ;
wire \i_post_norm_mul.s_infb  ;
wire \i_post_norm_mul.un1_s_infa  ;
wire \i_post_norm_mul.or_reduce.result_4  ;
wire N_536 ;
wire N_537 ;
wire N_538 ;
wire N_541 ;
wire N_542 ;
wire N_543 ;
wire N_544 ;
wire N_545 ;
wire N_546 ;
wire N_547 ;
wire N_548 ;
wire N_549 ;
wire N_550 ;
wire N_551 ;
wire N_552 ;
wire N_553 ;
wire N_554 ;
wire N_555 ;
wire N_556 ;
wire N_557 ;
wire N_558 ;
wire N_559 ;
wire N_560 ;
wire N_561 ;
wire N_562 ;
wire N_563 ;
wire N_564 ;
wire \i_post_norm_sqrt.or_reduce.result_11  ;
wire \i_post_norm_mul.un1_s_nan_a  ;
wire \i_post_norm_mul.un1_s_nan_b  ;
wire N_1979 ;
wire N_1948 ;
wire un2_s_snan_o_22 ;
wire \i_pre_norm_div.s_dvdnd_50_o.N_59  ;
wire un2_s_snan_o_8 ;
wire N_1166 ;
wire N_1087 ;
wire N_1227 ;
wire N_1174 ;
wire N_987 ;
wire N_1041 ;
wire un2_s_snan_o_20 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_44  ;
wire N_1241 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_88  ;
wire N_2103 ;
wire N_1620 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_53  ;
wire N_1619 ;
wire N_1624 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_46  ;
wire N_1238 ;
wire N_1242 ;
wire N_1617 ;
wire N_1245 ;
wire N_48_0 ;
wire N_36_0 ;
wire un1_s_infb ;
wire \i_postnorm_addsub.or_reduce.result_2  ;
wire N_1941 ;
wire \i_pre_norm_div.N_396  ;
wire \i_pre_norm_div.N_399  ;
wire N_1051 ;
wire N_2220 ;
wire N_1077 ;
wire \i_pre_norm_div.s_dvdnd_50_o.N_63  ;
wire \i_pre_norm_div.s_dvdnd_50_o.N_55  ;
wire N_1264 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_41  ;
wire N_1628 ;
wire N_27_0 ;
wire N_30_0 ;
wire N_38_0 ;
wire N_1236 ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_43  ;
wire N_1630 ;
wire \i_pre_norm_div.s_dvdnd_50_o.N_95  ;
wire \i_pre_norm_div.s_dvdnd_50_o.N_70  ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.N_45  ;
wire \i_postnorm_addsub.or_reduce.result_2_10  ;
wire N_1050 ;
wire N_143_mux ;
wire N_1083 ;
wire N_1055 ;
wire un4_s_infa ;
wire \i_pre_norm_div.s_dvsor_27_o.N_54  ;
wire \i_postnorm_addsub.or_reduce.result_2_16  ;
wire N_2240 ;
wire N_1170 ;
wire N_1140 ;
wire s_start_i ;
wire un1_s_count_4_s_0 ;
wire un1_s_count_4_s_1 ;
wire un1_s_count_4_s_2 ;
wire un1_s_count_4_s_3 ;
wire un1_s_count_4_s_4 ;
wire un1_s_count_4_s_5 ;
wire un1_s_count_4_s_6 ;
wire un1_s_count_4_s_7 ;
wire un1_s_count_4_s_8 ;
wire un1_s_count_4_s_9 ;
wire un1_s_count_4_s_10 ;
wire un1_s_count_4_s_11 ;
wire un1_s_count_4_s_12 ;
wire un1_s_count_4_s_13 ;
wire un1_s_count_4_s_14 ;
wire un1_s_count_4_s_15 ;
wire un1_s_count_4_s_16 ;
wire un1_s_count_4_s_17 ;
wire un1_s_count_4_s_18 ;
wire un1_s_count_4_s_19 ;
wire un1_s_count_4_s_20 ;
wire un1_s_count_4_s_21 ;
wire un1_s_count_4_s_22 ;
wire un1_s_count_4_s_23 ;
wire un1_s_count_4_s_24 ;
wire un1_s_count_4_s_25 ;
wire un1_s_count_4_s_26 ;
wire un1_s_count_4_s_27 ;
wire un1_s_count_4_s_28 ;
wire un1_s_count_4_s_29 ;
wire un1_s_count_4_s_30 ;
wire un1_s_count_4_s_31 ;
wire un1_s_count_4_axb_0 ;
wire un1_s_count_4_cry_0 ;
wire un1_s_count_4_axb_1 ;
wire un1_s_count_4_cry_1 ;
wire un1_s_count_4_axb_2 ;
wire un1_s_count_4_cry_2 ;
wire un1_s_count_4_axb_3 ;
wire un1_s_count_4_cry_3 ;
wire un1_s_count_4_axb_4 ;
wire un1_s_count_4_cry_4 ;
wire un1_s_count_4_axb_5 ;
wire un1_s_count_4_cry_5 ;
wire un1_s_count_4_axb_6 ;
wire un1_s_count_4_cry_6 ;
wire un1_s_count_4_axb_7 ;
wire un1_s_count_4_cry_7 ;
wire un1_s_count_4_axb_8 ;
wire un1_s_count_4_cry_8 ;
wire un1_s_count_4_axb_9 ;
wire un1_s_count_4_cry_9 ;
wire un1_s_count_4_axb_10 ;
wire un1_s_count_4_cry_10 ;
wire un1_s_count_4_axb_11 ;
wire un1_s_count_4_cry_11 ;
wire un1_s_count_4_axb_12 ;
wire un1_s_count_4_cry_12 ;
wire un1_s_count_4_axb_13 ;
wire un1_s_count_4_cry_13 ;
wire un1_s_count_4_axb_14 ;
wire un1_s_count_4_cry_14 ;
wire un1_s_count_4_axb_15 ;
wire un1_s_count_4_cry_15 ;
wire un1_s_count_4_axb_16 ;
wire un1_s_count_4_cry_16 ;
wire un1_s_count_4_axb_17 ;
wire un1_s_count_4_cry_17 ;
wire un1_s_count_4_axb_18 ;
wire un1_s_count_4_cry_18 ;
wire un1_s_count_4_axb_19 ;
wire un1_s_count_4_cry_19 ;
wire un1_s_count_4_axb_20 ;
wire un1_s_count_4_cry_20 ;
wire un1_s_count_4_axb_21 ;
wire un1_s_count_4_cry_21 ;
wire un1_s_count_4_axb_22 ;
wire un1_s_count_4_cry_22 ;
wire un1_s_count_4_axb_23 ;
wire un1_s_count_4_cry_23 ;
wire un1_s_count_4_axb_24 ;
wire un1_s_count_4_cry_24 ;
wire un1_s_count_4_axb_25 ;
wire un1_s_count_4_cry_25 ;
wire un1_s_count_4_axb_26 ;
wire un1_s_count_4_cry_26 ;
wire un1_s_count_4_axb_27 ;
wire un1_s_count_4_cry_27 ;
wire un1_s_count_4_axb_28 ;
wire un1_s_count_4_cry_28 ;
wire un1_s_count_4_axb_29 ;
wire un1_s_count_4_cry_29 ;
wire un1_s_count_4_axb_30 ;
wire un1_s_count_4_cry_30 ;
wire un1_s_count_4_axb_31 ;
wire N_1084_i ;
wire N_2637_i ;
wire N_503_i ;
wire N_502_i ;
wire N_501_i ;
wire N_1257_i ;
wire N_1278_i ;
wire N_1942_i ;
wire N_772_i ;
wire N_771_i ;
wire N_770_i ;
wire N_769_i ;
wire N_768_i ;
wire N_767_i ;
wire N_766_i ;
wire N_764_i ;
wire N_20_i ;
wire N_18_i ;
wire N_14_i ;
wire N_780_i ;
wire N_779_i ;
wire N_778_i ;
wire N_777_i ;
wire N_776_i ;
wire N_775_i ;
wire N_774_i ;
wire N_378_i ;
wire N_1232_i ;
wire \i_pre_norm_div.un4_s_expb_in_2_i_o2_0  ;
wire \i_pre_norm_div.un4_s_expb_in_2_i_o2_1  ;
wire \i_pre_norm_div.un4_s_expb_in_2_i_o2_2  ;
wire \i_post_norm_mul.or_reduce.result_3_21_1  ;
wire \i_post_norm_mul.or_reduce.result_3_21_3  ;
wire \i_prenorm_addsub.un4_s_infa_1  ;
wire \i_postnorm_addsub.or_reduce.result_2_2  ;
wire m16_0_0 ;
wire m16_0_1 ;
wire m16_0_3 ;
wire m16_0_4 ;
wire m16_0_2_3 ;
wire ready_o_0 ;
wire un1_s_count_4_cry_0_cy ;
wire \i_pre_norm_div.un11_s_exp_10_o_axb_0_i  ;
wire N_2715_0 ;
wire N_2745_0 ;
wire N_80_0_0 ;
wire N_81_0_0 ;
wire N_2746_0 ;
wire div_zero_o_0_0 ;
wire \or_reduce.result_i_0_0  ;
wire un3_s_underflow_o_0 ;
wire \i_pre_norm_div.un4_s_expb_in_2_i_0_e  ;
wire \i_pre_norm_div.or_reduce.result_1_i_o3_0_e  ;
wire \i_postnorm_addsub.un2_s_qnan_o_0_a2_0_e  ;
wire \i_postnorm_addsub.N_6_i_0_e  ;
wire \i_postnorm_addsub.N_9_i_0_e  ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_106_0_e  ;
wire \i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_107_0_e  ;
wire \i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_108_0_e  ;
wire \i_prenorm_addsub.m49_0_e  ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_105_0_e  ;
wire \i_prenorm_addsub.m46_0_e  ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_109_0_e  ;
wire \i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_102_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_108_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_104_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_106_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_102_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_105_0_e  ;
wire \i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_103_0_e  ;
wire \i_postnorm_addsub.N_773_i_0_e  ;
wire \i_postnorm_addsub.N_12_i_0_e  ;
wire \i_postnorm_addsub.N_763_i_0_e  ;
wire \i_postnorm_addsub.N_765_i_0_e  ;
wire \i_postnorm_addsub.or_reduce.result_3_0_0_i  ;
input p_desc595_p_O_FDpre_norm_mul_ ;
input p_desc596_p_O_FDpre_norm_mul_ ;
input p_desc597_p_O_FDpre_norm_mul_ ;
input p_desc598_p_O_FDpre_norm_mul_ ;
input p_desc599_p_O_FDpre_norm_mul_ ;
input p_desc600_p_O_FDpre_norm_mul_ ;
input p_desc601_p_O_FDpre_norm_mul_ ;
input p_desc602_p_O_FDpre_norm_mul_ ;
input p_desc603_p_O_FDpre_norm_mul_ ;
input p_desc604_p_O_FDpre_norm_mul_ ;
input p_desc1070_p_O_FDpost_norm_mul_ ;
input p_desc1071_p_O_FDpost_norm_mul_ ;
input p_desc1072_p_O_FDpost_norm_mul_ ;
input p_desc1073_p_O_FDpost_norm_mul_ ;
input p_desc1074_p_O_FDpost_norm_mul_ ;
input p_desc1075_p_O_FDpost_norm_mul_ ;
input p_desc1076_p_O_FDpost_norm_mul_ ;
input p_desc1077_p_O_FDpost_norm_mul_ ;
input p_desc1078_p_O_FDpost_norm_mul_ ;
input p_desc1079_p_O_FDpost_norm_mul_ ;
input p_desc1080_p_O_FDpost_norm_mul_ ;
input p_desc1081_p_O_FDpost_norm_mul_ ;
input p_desc1082_p_O_FDpost_norm_mul_ ;
input p_desc1083_p_O_FDpost_norm_mul_ ;
input p_desc1084_p_O_FDpost_norm_mul_ ;
input p_desc1085_p_O_FDpost_norm_mul_ ;
input p_desc1086_p_O_FDpost_norm_mul_ ;
input p_desc1087_p_O_FDpost_norm_mul_ ;
input p_desc1088_p_O_FDpost_norm_mul_ ;
input p_desc1089_p_O_FDpost_norm_mul_ ;
input p_desc1090_p_O_FDpost_norm_mul_ ;
input p_desc1091_p_O_FDpost_norm_mul_ ;
input p_desc1092_p_O_FDpost_norm_mul_ ;
input p_desc1163_p_O_FDpost_norm_mul_ ;
input p_desc1164_p_O_FDpost_norm_mul_ ;
input p_desc1165_p_O_FDpost_norm_mul_ ;
input p_desc1166_p_O_FDpost_norm_mul_ ;
input p_desc1167_p_O_FDpost_norm_mul_ ;
input p_desc1168_p_O_FDpost_norm_mul_ ;
input p_desc1169_p_O_FDpost_norm_mul_ ;
input p_desc1170_p_O_FDpost_norm_mul_ ;
input p_desc1171_p_O_FDpost_norm_mul_ ;
input p_desc1172_p_O_FDpost_norm_mul_ ;
input p_desc1173_p_O_FDpost_norm_mul_ ;
input p_desc1174_p_O_FDpost_norm_mul_ ;
input p_desc1175_p_O_FDpost_norm_mul_ ;
input p_desc1176_p_O_FDpost_norm_mul_ ;
input p_desc1177_p_O_FDpost_norm_mul_ ;
input p_desc1178_p_O_FDpost_norm_mul_ ;
input p_desc1179_p_O_FDpost_norm_mul_ ;
input p_desc1180_p_O_FDpost_norm_mul_ ;
input p_desc1181_p_O_FDpost_norm_mul_ ;
input p_desc1182_p_O_FDpost_norm_mul_ ;
input p_desc1183_p_O_FDpost_norm_mul_ ;
input p_desc1184_p_O_FDpost_norm_mul_ ;
input p_desc1185_p_O_FDpost_norm_mul_ ;
input p_desc1186_p_O_FDpost_norm_mul_ ;
input p_desc1187_p_O_FDpost_norm_mul_ ;
input p_desc1188_p_O_FDpost_norm_mul_ ;
input p_desc1189_p_O_FDpost_norm_mul_ ;
input p_desc1190_p_O_FDpost_norm_mul_ ;
input p_desc1191_p_O_FDpost_norm_mul_ ;
input p_desc1192_p_O_FDpost_norm_mul_ ;
input p_desc1193_p_O_FDpost_norm_mul_ ;
input p_desc1194_p_O_FDpost_norm_mul_ ;
input p_desc1195_p_O_FDpost_norm_mul_ ;
input p_desc1196_p_O_FDpost_norm_mul_ ;
input p_desc1197_p_O_FDpost_norm_mul_ ;
input p_desc1198_p_O_FDpost_norm_mul_ ;
input p_desc1199_p_O_FDpost_norm_mul_ ;
input p_desc1200_p_O_FDpost_norm_mul_ ;
input p_desc1201_p_O_FDpost_norm_mul_ ;
input p_desc1202_p_O_FDpost_norm_mul_ ;
input p_desc1203_p_O_FDpost_norm_mul_ ;
input p_desc1204_p_O_FDpost_norm_mul_ ;
input p_desc1205_p_O_FDpost_norm_mul_ ;
input p_desc1206_p_O_FDpost_norm_mul_ ;
input p_desc1207_p_O_FDpost_norm_mul_ ;
input p_desc1208_p_O_FDpost_norm_mul_ ;
input p_desc1209_p_O_FDpost_norm_mul_ ;
input p_desc1210_p_O_FDpost_norm_mul_ ;
input p_desc1211_p_O_FDpost_norm_mul_ ;
input p_desc1212_p_O_FDpost_norm_mul_ ;
input p_desc1213_p_O_FDpost_norm_mul_ ;
input p_desc1214_p_O_FDpost_norm_mul_ ;
input p_desc1215_p_O_FDpost_norm_mul_ ;
input p_desc1216_p_O_FDpost_norm_mul_ ;
input p_desc1217_p_O_FDpost_norm_mul_ ;
input p_desc1218_p_O_FDpost_norm_mul_ ;
input p_desc1219_p_O_FDpost_norm_mul_ ;
input p_desc1220_p_O_FDpost_norm_mul_ ;
input p_desc1221_p_O_FDpost_norm_mul_ ;
input p_s_sign_i_Z_p_O_FDpost_norm_mul_ ;
input p_ine_o_Z_p_O_FDpost_norm_mul_ ;
input p_desc1244_p_O_FDpost_norm_mul_ ;
input p_desc1245_p_O_FDpost_norm_mul_ ;
input p_desc1246_p_O_FDpost_norm_mul_ ;
input p_desc1247_p_O_FDpost_norm_mul_ ;
input p_desc1248_p_O_FDpost_norm_mul_ ;
input p_desc1249_p_O_FDpost_norm_mul_ ;
input p_desc1250_p_O_FDpost_norm_mul_ ;
input p_desc1251_p_O_FDpost_norm_mul_ ;
input p_desc1252_p_O_FDpost_norm_mul_ ;
input p_desc1253_p_O_FDpost_norm_mul_ ;
input p_desc1254_p_O_FDpost_norm_mul_ ;
input p_desc1255_p_O_FDpost_norm_mul_ ;
input p_desc1256_p_O_FDpost_norm_mul_ ;
input p_desc1257_p_O_FDpost_norm_mul_ ;
input p_desc1258_p_O_FDpost_norm_mul_ ;
input p_desc1259_p_O_FDpost_norm_mul_ ;
input p_desc1260_p_O_FDpost_norm_mul_ ;
input p_desc1261_p_O_FDpost_norm_mul_ ;
input p_desc1262_p_O_FDpost_norm_mul_ ;
input p_desc1263_p_O_FDpost_norm_mul_ ;
input p_desc1264_p_O_FDpost_norm_mul_ ;
input p_desc1265_p_O_FDpost_norm_mul_ ;
input p_desc1266_p_O_FDpost_norm_mul_ ;
input p_desc1267_p_O_FDpost_norm_mul_ ;
input p_desc1268_p_O_FDpost_norm_mul_ ;
input p_desc1269_p_O_FDpost_norm_mul_ ;
input p_desc1270_p_O_FDpost_norm_mul_ ;
input p_desc1271_p_O_FDpost_norm_mul_ ;
input p_desc1272_p_O_FDpost_norm_mul_ ;
input p_desc1273_p_O_FDpost_norm_mul_ ;
input p_desc1274_p_O_FDpost_norm_mul_ ;
input p_desc1275_p_O_FDpost_norm_mul_ ;
input p_desc1276_p_O_FDpost_norm_mul_ ;
input p_desc1277_p_O_FDpost_norm_mul_ ;
input p_desc1278_p_O_FDpost_norm_mul_ ;
input p_desc1279_p_O_FDpost_norm_mul_ ;
input p_desc1280_p_O_FDpost_norm_mul_ ;
input p_desc1281_p_O_FDpost_norm_mul_ ;
input p_desc1282_p_O_FDpost_norm_mul_ ;
input p_desc1283_p_O_FDpost_norm_mul_ ;
input p_desc1284_p_O_FDpost_norm_mul_ ;
input p_desc1285_p_O_FDpost_norm_mul_ ;
input p_desc1286_p_O_FDpost_norm_mul_ ;
input p_desc1287_p_O_FDpost_norm_mul_ ;
input p_desc1288_p_O_FDpost_norm_mul_ ;
input p_desc1289_p_O_FDpost_norm_mul_ ;
input p_desc1290_p_O_FDpost_norm_mul_ ;
input p_desc1291_p_O_FDpost_norm_mul_ ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  FD desc3350(.Q(output_o[14:14]),.D(\i_postnorm_addsub.N_773_i_0_e ),.C(clk_i));
  FD desc3351(.Q(output_o[0:0]),.D(\i_postnorm_addsub.N_12_i_0_e ),.C(clk_i));
  FD desc3352(.Q(output_o[2:2]),.D(\i_postnorm_addsub.N_763_i_0_e ),.C(clk_i));
  FD desc3353(.Q(output_o[6:6]),.D(\i_postnorm_addsub.N_765_i_0_e ),.C(clk_i));
  FD qnan_o_Z(.Q(qnan_o),.D(\i_postnorm_addsub.un2_s_qnan_o_0_a2_0_e ),.C(clk_i));
  FD overflow_o_Z(.Q(overflow_o),.D(\i_postnorm_addsub.N_6_i_0_e ),.C(clk_i));
  FD inf_o_Z(.Q(inf_o),.D(\i_postnorm_addsub.N_9_i_0_e ),.C(clk_i));
  FDSE desc3354(.Q(s_state),.D(GND),.C(clk_i),.S(s_start_i),.CE(s_count_RNIM79LF[21:21]));
  FDR desc3355(.Q(s_count[0:0]),.D(N_2746_0),.C(clk_i),.R(s_start_i));
  FDR desc3356(.Q(s_count[2:2]),.D(N_81_0_0),.C(clk_i),.R(s_start_i));
  FDR desc3357(.Q(s_count[3:3]),.D(N_80_0_0),.C(clk_i),.R(s_start_i));
  FDR desc3358(.Q(s_count[5:5]),.D(N_2745_0),.C(clk_i),.R(s_start_i));
  FDR desc3359(.Q(s_count[1:1]),.D(N_2715_0),.C(clk_i),.R(s_start_i));
  LUT1 un1_s_count_4_axb_0_cZ(.I0(s_count[0:0]),.O(un1_s_count_4_axb_0));
defparam un1_s_count_4_axb_0_cZ.INIT=2'h2;
  LUT1 un1_s_count_4_axb_1_cZ(.I0(s_count[1:1]),.O(un1_s_count_4_axb_1));
defparam un1_s_count_4_axb_1_cZ.INIT=2'h2;
  LUT1 un1_s_count_4_axb_2_cZ(.I0(s_count[2:2]),.O(un1_s_count_4_axb_2));
defparam un1_s_count_4_axb_2_cZ.INIT=2'h2;
  LUT1 un1_s_count_4_axb_3_cZ(.I0(s_count[3:3]),.O(un1_s_count_4_axb_3));
defparam un1_s_count_4_axb_3_cZ.INIT=2'h2;
  LUT1 un1_s_count_4_axb_5_cZ(.I0(s_count[5:5]),.O(un1_s_count_4_axb_5));
defparam un1_s_count_4_axb_5_cZ.INIT=2'h2;
  LUT2 un1_s_count_4_cry_0_cy_RNO_cZ(.I0(s_count_RNIM79LF[21:21]),.I1(s_state),.O(un1_s_count_4_cry_0_cy_RNO));
defparam un1_s_count_4_cry_0_cy_RNO_cZ.INIT=4'h4;
  FD ready_o_Z(.Q(ready_o),.D(ready_o_0),.C(clk_i));
  FD desc3360(.Q(s_opb_i[18:18]),.D(opb_i[18:18]),.C(clk_i));
  FD desc3361(.Q(s_opb_i[19:19]),.D(opb_i[19:19]),.C(clk_i));
  FD desc3362(.Q(s_opb_i[20:20]),.D(opb_i[20:20]),.C(clk_i));
  FD desc3363(.Q(s_opb_i[21:21]),.D(opb_i[21:21]),.C(clk_i));
  FD desc3364(.Q(s_opb_i[22:22]),.D(opb_i[22:22]),.C(clk_i));
  FD desc3365(.Q(s_opb_i[23:23]),.D(opb_i[23:23]),.C(clk_i));
  FD desc3366(.Q(s_opb_i[24:24]),.D(opb_i[24:24]),.C(clk_i));
  FD desc3367(.Q(s_opb_i[25:25]),.D(opb_i[25:25]),.C(clk_i));
  FD desc3368(.Q(s_opb_i[26:26]),.D(opb_i[26:26]),.C(clk_i));
  FD desc3369(.Q(s_opb_i[27:27]),.D(opb_i[27:27]),.C(clk_i));
  FD desc3370(.Q(s_opb_i[28:28]),.D(opb_i[28:28]),.C(clk_i));
  FD desc3371(.Q(s_opb_i[29:29]),.D(opb_i[29:29]),.C(clk_i));
  FD desc3372(.Q(s_opb_i[30:30]),.D(opb_i[30:30]),.C(clk_i));
  FD desc3373(.Q(s_opb_i[31:31]),.D(opb_i[31:31]),.C(clk_i));
  FD desc3374(.Q(s_opb_i[3:3]),.D(opb_i[3:3]),.C(clk_i));
  FD desc3375(.Q(s_opb_i[4:4]),.D(opb_i[4:4]),.C(clk_i));
  FD desc3376(.Q(s_opb_i[5:5]),.D(opb_i[5:5]),.C(clk_i));
  FD desc3377(.Q(s_opb_i[6:6]),.D(opb_i[6:6]),.C(clk_i));
  FD desc3378(.Q(s_opb_i[7:7]),.D(opb_i[7:7]),.C(clk_i));
  FD desc3379(.Q(s_opb_i[8:8]),.D(opb_i[8:8]),.C(clk_i));
  FD desc3380(.Q(s_opb_i[9:9]),.D(opb_i[9:9]),.C(clk_i));
  FD desc3381(.Q(s_opb_i[10:10]),.D(opb_i[10:10]),.C(clk_i));
  FD desc3382(.Q(s_opb_i[11:11]),.D(opb_i[11:11]),.C(clk_i));
  FD desc3383(.Q(s_opb_i[12:12]),.D(opb_i[12:12]),.C(clk_i));
  FD desc3384(.Q(s_opb_i[13:13]),.D(opb_i[13:13]),.C(clk_i));
  FD desc3385(.Q(s_opb_i[14:14]),.D(opb_i[14:14]),.C(clk_i));
  FD desc3386(.Q(s_opb_i[15:15]),.D(opb_i[15:15]),.C(clk_i));
  FD desc3387(.Q(s_opb_i[16:16]),.D(opb_i[16:16]),.C(clk_i));
  FD desc3388(.Q(s_opb_i[17:17]),.D(opb_i[17:17]),.C(clk_i));
  FD desc3389(.Q(s_opa_i[20:20]),.D(opa_i[20:20]),.C(clk_i));
  FD desc3390(.Q(s_opa_i[21:21]),.D(opa_i[21:21]),.C(clk_i));
  FD desc3391(.Q(s_opa_i[22:22]),.D(opa_i[22:22]),.C(clk_i));
  FD desc3392(.Q(s_opa_i[23:23]),.D(opa_i[23:23]),.C(clk_i));
  FD desc3393(.Q(s_opa_i[24:24]),.D(opa_i[24:24]),.C(clk_i));
  FD desc3394(.Q(s_opa_i[25:25]),.D(opa_i[25:25]),.C(clk_i));
  FD desc3395(.Q(s_opa_i[26:26]),.D(opa_i[26:26]),.C(clk_i));
  FD desc3396(.Q(s_opa_i[27:27]),.D(opa_i[27:27]),.C(clk_i));
  FD desc3397(.Q(s_opa_i[28:28]),.D(opa_i[28:28]),.C(clk_i));
  FD desc3398(.Q(s_opa_i[29:29]),.D(opa_i[29:29]),.C(clk_i));
  FD desc3399(.Q(s_opa_i[30:30]),.D(opa_i[30:30]),.C(clk_i));
  FD desc3400(.Q(s_opa_i[31:31]),.D(opa_i[31:31]),.C(clk_i));
  FD desc3401(.Q(s_opb_i[0:0]),.D(opb_i[0:0]),.C(clk_i));
  FD desc3402(.Q(s_opb_i[1:1]),.D(opb_i[1:1]),.C(clk_i));
  FD desc3403(.Q(s_opb_i[2:2]),.D(opb_i[2:2]),.C(clk_i));
  FD desc3404(.Q(s_opa_i[5:5]),.D(opa_i[5:5]),.C(clk_i));
  FD desc3405(.Q(s_opa_i[6:6]),.D(opa_i[6:6]),.C(clk_i));
  FD desc3406(.Q(s_opa_i[7:7]),.D(opa_i[7:7]),.C(clk_i));
  FD desc3407(.Q(s_opa_i[8:8]),.D(opa_i[8:8]),.C(clk_i));
  FD desc3408(.Q(s_opa_i[9:9]),.D(opa_i[9:9]),.C(clk_i));
  FD desc3409(.Q(s_opa_i[10:10]),.D(opa_i[10:10]),.C(clk_i));
  FD desc3410(.Q(s_opa_i[11:11]),.D(opa_i[11:11]),.C(clk_i));
  FD desc3411(.Q(s_opa_i[12:12]),.D(opa_i[12:12]),.C(clk_i));
  FD desc3412(.Q(s_opa_i[13:13]),.D(opa_i[13:13]),.C(clk_i));
  FD desc3413(.Q(s_opa_i[14:14]),.D(opa_i[14:14]),.C(clk_i));
  FD desc3414(.Q(s_opa_i[15:15]),.D(opa_i[15:15]),.C(clk_i));
  FD desc3415(.Q(s_opa_i[16:16]),.D(opa_i[16:16]),.C(clk_i));
  FD desc3416(.Q(s_opa_i[17:17]),.D(opa_i[17:17]),.C(clk_i));
  FD desc3417(.Q(s_opa_i[18:18]),.D(opa_i[18:18]),.C(clk_i));
  FD desc3418(.Q(s_opa_i[19:19]),.D(opa_i[19:19]),.C(clk_i));
  FD desc3419(.Q(s_rmode_i[0:0]),.D(rmode_i[0:0]),.C(clk_i));
  FD desc3420(.Q(s_rmode_i[1:1]),.D(rmode_i[1:1]),.C(clk_i));
  FD desc3421(.Q(s_fpu_op_i[0:0]),.D(fpu_op_i[0:0]),.C(clk_i));
  FD desc3422(.Q(s_fpu_op_i[1:1]),.D(fpu_op_i[1:1]),.C(clk_i));
  FD desc3423(.Q(s_fpu_op_i[2:2]),.D(fpu_op_i[2:2]),.C(clk_i));
  FD desc3424(.Q(s_opa_i[0:0]),.D(opa_i[0:0]),.C(clk_i));
  FD desc3425(.Q(s_opa_i[1:1]),.D(opa_i[1:1]),.C(clk_i));
  FD desc3426(.Q(s_opa_i[2:2]),.D(opa_i[2:2]),.C(clk_i));
  FD desc3427(.Q(s_opa_i[3:3]),.D(opa_i[3:3]),.C(clk_i));
  FD desc3428(.Q(s_opa_i[4:4]),.D(opa_i[4:4]),.C(clk_i));
  FD desc3429(.Q(output_o[29:29]),.D(s_output1[29:29]),.C(clk_i));
  FD desc3430(.Q(output_o[30:30]),.D(s_output1[30:30]),.C(clk_i));
  FD desc3431(.Q(output_o[31:31]),.D(s_output_o_0[31:31]),.C(clk_i));
  FD desc3432(.Q(output_o[15:15]),.D(N_774_i),.C(clk_i));
  FD desc3433(.Q(output_o[16:16]),.D(N_775_i),.C(clk_i));
  FD desc3434(.Q(output_o[17:17]),.D(N_776_i),.C(clk_i));
  FD desc3435(.Q(output_o[18:18]),.D(N_777_i),.C(clk_i));
  FD desc3436(.Q(output_o[19:19]),.D(N_778_i),.C(clk_i));
  FD desc3437(.Q(output_o[20:20]),.D(N_779_i),.C(clk_i));
  FD desc3438(.Q(output_o[21:21]),.D(N_780_i),.C(clk_i));
  FD desc3439(.Q(output_o[22:22]),.D(s_output_o_0[22:22]),.C(clk_i));
  FD desc3440(.Q(output_o[23:23]),.D(s_output_o[23:23]),.C(clk_i));
  FD desc3441(.Q(output_o[24:24]),.D(s_output1[24:24]),.C(clk_i));
  FD desc3442(.Q(output_o[25:25]),.D(s_output1[25:25]),.C(clk_i));
  FD desc3443(.Q(output_o[26:26]),.D(s_output1[26:26]),.C(clk_i));
  FD desc3444(.Q(output_o[27:27]),.D(s_output1[27:27]),.C(clk_i));
  FD desc3445(.Q(output_o[28:28]),.D(s_output1[28:28]),.C(clk_i));
  FD desc3446(.Q(output_o[1:1]),.D(N_14_i),.C(clk_i));
  FD desc3447(.Q(output_o[3:3]),.D(N_18_i),.C(clk_i));
  FD desc3448(.Q(output_o[4:4]),.D(N_20_i),.C(clk_i));
  FD desc3449(.Q(output_o[5:5]),.D(N_764_i),.C(clk_i));
  FD desc3450(.Q(output_o[7:7]),.D(N_766_i),.C(clk_i));
  FD desc3451(.Q(output_o[8:8]),.D(N_767_i),.C(clk_i));
  FD desc3452(.Q(output_o[9:9]),.D(N_768_i),.C(clk_i));
  FD desc3453(.Q(output_o[10:10]),.D(N_769_i),.C(clk_i));
  FD desc3454(.Q(output_o[11:11]),.D(N_770_i),.C(clk_i));
  FD desc3455(.Q(output_o[12:12]),.D(N_771_i),.C(clk_i));
  FD desc3456(.Q(output_o[13:13]),.D(N_772_i),.C(clk_i));
  FD zero_o_Z(.Q(zero_o),.D(\or_reduce.result_i_0_0 ),.C(clk_i));
  FD s_start_i_Z(.Q(s_start_i),.D(start_i),.C(clk_i));
  FD underflow_o_Z(.Q(underflow_o),.D(un3_s_underflow_o_0),.C(clk_i));
  FD snan_o_Z(.Q(snan_o),.D(un3_s_snan_o_0),.C(clk_i));
  FD s_ine_o_Z(.Q(s_ine_o),.D(s_ine_o_5),.C(clk_i));
  FD ine_o_Z(.Q(ine_o),.D(s_ine_o),.C(clk_i));
  FDR desc3457(.Q(s_output1[27:27]),.D(N_560),.C(clk_i),.R(N_2637_i));
  FDR desc3458(.Q(s_output1[28:28]),.D(N_561),.C(clk_i),.R(N_2637_i));
  FDR desc3459(.Q(s_output1[29:29]),.D(N_562),.C(clk_i),.R(N_2637_i));
  FDR desc3460(.Q(s_output1[30:30]),.D(N_563),.C(clk_i),.R(N_2637_i));
  FDR desc3461(.Q(s_output1[31:31]),.D(N_564),.C(clk_i),.R(N_2637_i));
  FDR desc3462(.Q(s_output1[12:12]),.D(N_545),.C(clk_i),.R(N_2637_i));
  FDR desc3463(.Q(s_output1[13:13]),.D(N_546),.C(clk_i),.R(N_2637_i));
  FDR desc3464(.Q(s_output1[14:14]),.D(N_547),.C(clk_i),.R(N_2637_i));
  FDR desc3465(.Q(s_output1[15:15]),.D(N_548),.C(clk_i),.R(N_2637_i));
  FDR desc3466(.Q(s_output1[16:16]),.D(N_549),.C(clk_i),.R(N_2637_i));
  FDR desc3467(.Q(s_output1[17:17]),.D(N_550),.C(clk_i),.R(N_2637_i));
  FDR desc3468(.Q(s_output1[18:18]),.D(N_551),.C(clk_i),.R(N_2637_i));
  FDR desc3469(.Q(s_output1[19:19]),.D(N_552),.C(clk_i),.R(N_2637_i));
  FDR desc3470(.Q(s_output1[20:20]),.D(N_553),.C(clk_i),.R(N_2637_i));
  FDR desc3471(.Q(s_output1[21:21]),.D(N_554),.C(clk_i),.R(N_2637_i));
  FDR desc3472(.Q(s_output1[22:22]),.D(N_555),.C(clk_i),.R(N_2637_i));
  FDR desc3473(.Q(s_output1[23:23]),.D(N_556),.C(clk_i),.R(N_2637_i));
  FDR desc3474(.Q(s_output1[24:24]),.D(N_557),.C(clk_i),.R(N_2637_i));
  FDR desc3475(.Q(s_output1[25:25]),.D(N_558),.C(clk_i),.R(N_2637_i));
  FDR desc3476(.Q(s_output1[26:26]),.D(N_559),.C(clk_i),.R(N_2637_i));
  FDR desc3477(.Q(s_output1[0:0]),.D(N_501_i),.C(clk_i),.R(N_2637_i));
  FDR desc3478(.Q(s_output1[1:1]),.D(N_502_i),.C(clk_i),.R(N_2637_i));
  FDR desc3479(.Q(s_output1[2:2]),.D(N_503_i),.C(clk_i),.R(N_2637_i));
  FDR desc3480(.Q(s_output1[3:3]),.D(N_536),.C(clk_i),.R(N_2637_i));
  FDR desc3481(.Q(s_output1[4:4]),.D(N_537),.C(clk_i),.R(N_2637_i));
  FDR desc3482(.Q(s_output1[5:5]),.D(N_538),.C(clk_i),.R(N_2637_i));
  FDR desc3483(.Q(s_output1[6:6]),.D(s_output1_6_2_i_m2[6:6]),.C(clk_i),.R(N_2637_i));
  FDR desc3484(.Q(s_output1[7:7]),.D(s_output1_6_2_i_m2[7:7]),.C(clk_i),.R(N_2637_i));
  FDR desc3485(.Q(s_output1[8:8]),.D(N_541),.C(clk_i),.R(N_2637_i));
  FDR desc3486(.Q(s_output1[9:9]),.D(N_542),.C(clk_i),.R(N_2637_i));
  FDR desc3487(.Q(s_output1[10:10]),.D(N_543),.C(clk_i),.R(N_2637_i));
  FDR desc3488(.Q(s_output1[11:11]),.D(N_544),.C(clk_i),.R(N_2637_i));
  FDR desc3489(.Q(s_count[31:31]),.D(un1_s_count_4_s_31),.C(clk_i),.R(s_start_i));
  FDR desc3490(.Q(s_count[16:16]),.D(un1_s_count_4_s_16),.C(clk_i),.R(s_start_i));
  FDR desc3491(.Q(s_count[17:17]),.D(un1_s_count_4_s_17),.C(clk_i),.R(s_start_i));
  FDR desc3492(.Q(s_count[18:18]),.D(un1_s_count_4_s_18),.C(clk_i),.R(s_start_i));
  FDR desc3493(.Q(s_count[19:19]),.D(un1_s_count_4_s_19),.C(clk_i),.R(s_start_i));
  FDR desc3494(.Q(s_count[20:20]),.D(un1_s_count_4_s_20),.C(clk_i),.R(s_start_i));
  FDR desc3495(.Q(s_count[21:21]),.D(un1_s_count_4_s_21),.C(clk_i),.R(s_start_i));
  FDR desc3496(.Q(s_count[22:22]),.D(un1_s_count_4_s_22),.C(clk_i),.R(s_start_i));
  FDR desc3497(.Q(s_count[23:23]),.D(un1_s_count_4_s_23),.C(clk_i),.R(s_start_i));
  FDR desc3498(.Q(s_count[24:24]),.D(un1_s_count_4_s_24),.C(clk_i),.R(s_start_i));
  FDR desc3499(.Q(s_count[25:25]),.D(un1_s_count_4_s_25),.C(clk_i),.R(s_start_i));
  FDR desc3500(.Q(s_count[26:26]),.D(un1_s_count_4_s_26),.C(clk_i),.R(s_start_i));
  FDR desc3501(.Q(s_count[27:27]),.D(un1_s_count_4_s_27),.C(clk_i),.R(s_start_i));
  FDR desc3502(.Q(s_count[28:28]),.D(un1_s_count_4_s_28),.C(clk_i),.R(s_start_i));
  FDR desc3503(.Q(s_count[29:29]),.D(un1_s_count_4_s_29),.C(clk_i),.R(s_start_i));
  FDR desc3504(.Q(s_count[30:30]),.D(un1_s_count_4_s_30),.C(clk_i),.R(s_start_i));
  FDR desc3505(.Q(s_count[4:4]),.D(un1_s_count_4_s_4),.C(clk_i),.R(s_start_i));
  FDR desc3506(.Q(s_count[6:6]),.D(un1_s_count_4_s_6),.C(clk_i),.R(s_start_i));
  FDR desc3507(.Q(s_count[7:7]),.D(un1_s_count_4_s_7),.C(clk_i),.R(s_start_i));
  FDR desc3508(.Q(s_count[8:8]),.D(un1_s_count_4_s_8),.C(clk_i),.R(s_start_i));
  FDR desc3509(.Q(s_count[9:9]),.D(un1_s_count_4_s_9),.C(clk_i),.R(s_start_i));
  FDR desc3510(.Q(s_count[10:10]),.D(un1_s_count_4_s_10),.C(clk_i),.R(s_start_i));
  FDR desc3511(.Q(s_count[11:11]),.D(un1_s_count_4_s_11),.C(clk_i),.R(s_start_i));
  FDR desc3512(.Q(s_count[12:12]),.D(un1_s_count_4_s_12),.C(clk_i),.R(s_start_i));
  FDR desc3513(.Q(s_count[13:13]),.D(un1_s_count_4_s_13),.C(clk_i),.R(s_start_i));
  FDR desc3514(.Q(s_count[14:14]),.D(un1_s_count_4_s_14),.C(clk_i),.R(s_start_i));
  FDR desc3515(.Q(s_count[15:15]),.D(un1_s_count_4_s_15),.C(clk_i),.R(s_start_i));
  MUXCY_L un1_s_count_4_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_s_count_4_cry_0_cy_RNO),.LO(un1_s_count_4_cry_0_cy));
  FD div_zero_o_Z(.Q(div_zero_o),.D(div_zero_o_0_0),.C(clk_i));
  LUT1_L desc3516(.I0(s_opa_i[29:29]),.LO(s_opa_i_i[29:29]));
defparam desc3516.INIT=2'h1;
  LUT1_L desc3517(.I0(s_opa_i[28:28]),.LO(s_opa_i_i[28:28]));
defparam desc3517.INIT=2'h1;
  LUT1_L un1_s_count_4_axb_31_cZ(.I0(s_count[31:31]),.LO(un1_s_count_4_axb_31));
defparam un1_s_count_4_axb_31_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_30_cZ(.I0(s_count[30:30]),.LO(un1_s_count_4_axb_30));
defparam un1_s_count_4_axb_30_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_29_cZ(.I0(s_count[29:29]),.LO(un1_s_count_4_axb_29));
defparam un1_s_count_4_axb_29_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_28_cZ(.I0(s_count[28:28]),.LO(un1_s_count_4_axb_28));
defparam un1_s_count_4_axb_28_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_27_cZ(.I0(s_count[27:27]),.LO(un1_s_count_4_axb_27));
defparam un1_s_count_4_axb_27_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_26_cZ(.I0(s_count[26:26]),.LO(un1_s_count_4_axb_26));
defparam un1_s_count_4_axb_26_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_25_cZ(.I0(s_count[25:25]),.LO(un1_s_count_4_axb_25));
defparam un1_s_count_4_axb_25_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_24_cZ(.I0(s_count[24:24]),.LO(un1_s_count_4_axb_24));
defparam un1_s_count_4_axb_24_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_23_cZ(.I0(s_count[23:23]),.LO(un1_s_count_4_axb_23));
defparam un1_s_count_4_axb_23_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_22_cZ(.I0(s_count[22:22]),.LO(un1_s_count_4_axb_22));
defparam un1_s_count_4_axb_22_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_21_cZ(.I0(s_count[21:21]),.LO(un1_s_count_4_axb_21));
defparam un1_s_count_4_axb_21_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_20_cZ(.I0(s_count[20:20]),.LO(un1_s_count_4_axb_20));
defparam un1_s_count_4_axb_20_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_19_cZ(.I0(s_count[19:19]),.LO(un1_s_count_4_axb_19));
defparam un1_s_count_4_axb_19_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_18_cZ(.I0(s_count[18:18]),.LO(un1_s_count_4_axb_18));
defparam un1_s_count_4_axb_18_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_17_cZ(.I0(s_count[17:17]),.LO(un1_s_count_4_axb_17));
defparam un1_s_count_4_axb_17_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_16_cZ(.I0(s_count[16:16]),.LO(un1_s_count_4_axb_16));
defparam un1_s_count_4_axb_16_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_15_cZ(.I0(s_count[15:15]),.LO(un1_s_count_4_axb_15));
defparam un1_s_count_4_axb_15_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_14_cZ(.I0(s_count[14:14]),.LO(un1_s_count_4_axb_14));
defparam un1_s_count_4_axb_14_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_13_cZ(.I0(s_count[13:13]),.LO(un1_s_count_4_axb_13));
defparam un1_s_count_4_axb_13_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_12_cZ(.I0(s_count[12:12]),.LO(un1_s_count_4_axb_12));
defparam un1_s_count_4_axb_12_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_11_cZ(.I0(s_count[11:11]),.LO(un1_s_count_4_axb_11));
defparam un1_s_count_4_axb_11_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_10_cZ(.I0(s_count[10:10]),.LO(un1_s_count_4_axb_10));
defparam un1_s_count_4_axb_10_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_9_cZ(.I0(s_count[9:9]),.LO(un1_s_count_4_axb_9));
defparam un1_s_count_4_axb_9_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_8_cZ(.I0(s_count[8:8]),.LO(un1_s_count_4_axb_8));
defparam un1_s_count_4_axb_8_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_7_cZ(.I0(s_count[7:7]),.LO(un1_s_count_4_axb_7));
defparam un1_s_count_4_axb_7_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_6_cZ(.I0(s_count[6:6]),.LO(un1_s_count_4_axb_6));
defparam un1_s_count_4_axb_6_cZ.INIT=2'h2;
  LUT1_L un1_s_count_4_axb_4_cZ(.I0(s_count[4:4]),.LO(un1_s_count_4_axb_4));
defparam un1_s_count_4_axb_4_cZ.INIT=2'h2;
  LUT4 desc3518(.I0(s_count[17:17]),.I1(s_count[18:18]),.I2(s_count[19:19]),.I3(s_count[20:20]),.O(m16_0_2_3));
defparam desc3518.INIT=16'h0001;
  LUT6 desc3519(.I0(s_count[4:4]),.I1(s_count[6:6]),.I2(s_count[7:7]),.I3(s_count[14:14]),.I4(s_count[15:15]),.I5(s_count[16:16]),.O(m16_0_3));
defparam desc3519.INIT=64'h0000000000000001;
  LUT6 desc3520(.I0(s_count[23:23]),.I1(s_count[24:24]),.I2(s_count[25:25]),.I3(s_count[26:26]),.I4(s_count[27:27]),.I5(s_count[28:28]),.O(m16_0_1));
defparam desc3520.INIT=64'h0000000000000001;
  LUT6 desc3521(.I0(s_count[8:8]),.I1(s_count[9:9]),.I2(s_count[10:10]),.I3(s_count[29:29]),.I4(s_count[30:30]),.I5(s_count[31:31]),.O(m16_0_0));
defparam desc3521.INIT=64'h0000000000000001;
  LUT5 desc3522(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(fpu_op_i[2:2]),.I3(s_count[0:0]),.I4(s_count[2:2]),.O(s_count_RNIME821));
defparam desc3522.INIT=32'h00001800;
  LUT6_L desc3523(.I0(fpu_op_i[0:0]),.I1(fpu_op_i[1:1]),.I2(fpu_op_i[2:2]),.I3(s_count[0:0]),.I4(s_count[2:2]),.I5(s_count[3:3]),.LO(s_count_RNIS5BE1));
defparam desc3523.INIT=64'h0000040000030000;
  LUT5_L desc3524(.I0(s_count[11:11]),.I1(s_count[12:12]),.I2(s_count[13:13]),.I3(m16_0_0),.I4(m16_0_1),.LO(m16_0_4));
defparam desc3524.INIT=32'h01000000;
  LUT5 desc3525(.I0(s_count[1:1]),.I1(s_count[5:5]),.I2(s_count[3:3]),.I3(s_count_RNIME821),.I4(s_count_RNIS5BE1),.O(i155_mux));
defparam desc3525.INIT=32'h26220400;
  LUT6 desc3526(.I0(s_count[21:21]),.I1(s_count[22:22]),.I2(m16_0_2_3),.I3(m16_0_3),.I4(i155_mux),.I5(m16_0_4),.O(s_count_RNIM79LF[21:21]));
defparam desc3526.INIT=64'h1000000000000000;
  XORCY un1_s_count_4_s_31_cZ(.LI(un1_s_count_4_axb_31),.CI(un1_s_count_4_cry_30),.O(un1_s_count_4_s_31));
  XORCY un1_s_count_4_s_30_cZ(.LI(un1_s_count_4_axb_30),.CI(un1_s_count_4_cry_29),.O(un1_s_count_4_s_30));
  MUXCY_L un1_s_count_4_cry_30_cZ(.DI(GND),.CI(un1_s_count_4_cry_29),.S(un1_s_count_4_axb_30),.LO(un1_s_count_4_cry_30));
  XORCY un1_s_count_4_s_29_cZ(.LI(un1_s_count_4_axb_29),.CI(un1_s_count_4_cry_28),.O(un1_s_count_4_s_29));
  MUXCY_L un1_s_count_4_cry_29_cZ(.DI(GND),.CI(un1_s_count_4_cry_28),.S(un1_s_count_4_axb_29),.LO(un1_s_count_4_cry_29));
  XORCY un1_s_count_4_s_28_cZ(.LI(un1_s_count_4_axb_28),.CI(un1_s_count_4_cry_27),.O(un1_s_count_4_s_28));
  MUXCY_L un1_s_count_4_cry_28_cZ(.DI(GND),.CI(un1_s_count_4_cry_27),.S(un1_s_count_4_axb_28),.LO(un1_s_count_4_cry_28));
  XORCY un1_s_count_4_s_27_cZ(.LI(un1_s_count_4_axb_27),.CI(un1_s_count_4_cry_26),.O(un1_s_count_4_s_27));
  MUXCY_L un1_s_count_4_cry_27_cZ(.DI(GND),.CI(un1_s_count_4_cry_26),.S(un1_s_count_4_axb_27),.LO(un1_s_count_4_cry_27));
  XORCY un1_s_count_4_s_26_cZ(.LI(un1_s_count_4_axb_26),.CI(un1_s_count_4_cry_25),.O(un1_s_count_4_s_26));
  MUXCY_L un1_s_count_4_cry_26_cZ(.DI(GND),.CI(un1_s_count_4_cry_25),.S(un1_s_count_4_axb_26),.LO(un1_s_count_4_cry_26));
  XORCY un1_s_count_4_s_25_cZ(.LI(un1_s_count_4_axb_25),.CI(un1_s_count_4_cry_24),.O(un1_s_count_4_s_25));
  MUXCY_L un1_s_count_4_cry_25_cZ(.DI(GND),.CI(un1_s_count_4_cry_24),.S(un1_s_count_4_axb_25),.LO(un1_s_count_4_cry_25));
  XORCY un1_s_count_4_s_24_cZ(.LI(un1_s_count_4_axb_24),.CI(un1_s_count_4_cry_23),.O(un1_s_count_4_s_24));
  MUXCY_L un1_s_count_4_cry_24_cZ(.DI(GND),.CI(un1_s_count_4_cry_23),.S(un1_s_count_4_axb_24),.LO(un1_s_count_4_cry_24));
  XORCY un1_s_count_4_s_23_cZ(.LI(un1_s_count_4_axb_23),.CI(un1_s_count_4_cry_22),.O(un1_s_count_4_s_23));
  MUXCY_L un1_s_count_4_cry_23_cZ(.DI(GND),.CI(un1_s_count_4_cry_22),.S(un1_s_count_4_axb_23),.LO(un1_s_count_4_cry_23));
  XORCY un1_s_count_4_s_22_cZ(.LI(un1_s_count_4_axb_22),.CI(un1_s_count_4_cry_21),.O(un1_s_count_4_s_22));
  MUXCY_L un1_s_count_4_cry_22_cZ(.DI(GND),.CI(un1_s_count_4_cry_21),.S(un1_s_count_4_axb_22),.LO(un1_s_count_4_cry_22));
  XORCY un1_s_count_4_s_21_cZ(.LI(un1_s_count_4_axb_21),.CI(un1_s_count_4_cry_20),.O(un1_s_count_4_s_21));
  MUXCY_L un1_s_count_4_cry_21_cZ(.DI(GND),.CI(un1_s_count_4_cry_20),.S(un1_s_count_4_axb_21),.LO(un1_s_count_4_cry_21));
  XORCY un1_s_count_4_s_20_cZ(.LI(un1_s_count_4_axb_20),.CI(un1_s_count_4_cry_19),.O(un1_s_count_4_s_20));
  MUXCY_L un1_s_count_4_cry_20_cZ(.DI(GND),.CI(un1_s_count_4_cry_19),.S(un1_s_count_4_axb_20),.LO(un1_s_count_4_cry_20));
  XORCY un1_s_count_4_s_19_cZ(.LI(un1_s_count_4_axb_19),.CI(un1_s_count_4_cry_18),.O(un1_s_count_4_s_19));
  MUXCY_L un1_s_count_4_cry_19_cZ(.DI(GND),.CI(un1_s_count_4_cry_18),.S(un1_s_count_4_axb_19),.LO(un1_s_count_4_cry_19));
  XORCY un1_s_count_4_s_18_cZ(.LI(un1_s_count_4_axb_18),.CI(un1_s_count_4_cry_17),.O(un1_s_count_4_s_18));
  MUXCY_L un1_s_count_4_cry_18_cZ(.DI(GND),.CI(un1_s_count_4_cry_17),.S(un1_s_count_4_axb_18),.LO(un1_s_count_4_cry_18));
  XORCY un1_s_count_4_s_17_cZ(.LI(un1_s_count_4_axb_17),.CI(un1_s_count_4_cry_16),.O(un1_s_count_4_s_17));
  MUXCY_L un1_s_count_4_cry_17_cZ(.DI(GND),.CI(un1_s_count_4_cry_16),.S(un1_s_count_4_axb_17),.LO(un1_s_count_4_cry_17));
  XORCY un1_s_count_4_s_16_cZ(.LI(un1_s_count_4_axb_16),.CI(un1_s_count_4_cry_15),.O(un1_s_count_4_s_16));
  MUXCY_L un1_s_count_4_cry_16_cZ(.DI(GND),.CI(un1_s_count_4_cry_15),.S(un1_s_count_4_axb_16),.LO(un1_s_count_4_cry_16));
  XORCY un1_s_count_4_s_15_cZ(.LI(un1_s_count_4_axb_15),.CI(un1_s_count_4_cry_14),.O(un1_s_count_4_s_15));
  MUXCY_L un1_s_count_4_cry_15_cZ(.DI(GND),.CI(un1_s_count_4_cry_14),.S(un1_s_count_4_axb_15),.LO(un1_s_count_4_cry_15));
  XORCY un1_s_count_4_s_14_cZ(.LI(un1_s_count_4_axb_14),.CI(un1_s_count_4_cry_13),.O(un1_s_count_4_s_14));
  MUXCY_L un1_s_count_4_cry_14_cZ(.DI(GND),.CI(un1_s_count_4_cry_13),.S(un1_s_count_4_axb_14),.LO(un1_s_count_4_cry_14));
  XORCY un1_s_count_4_s_13_cZ(.LI(un1_s_count_4_axb_13),.CI(un1_s_count_4_cry_12),.O(un1_s_count_4_s_13));
  MUXCY_L un1_s_count_4_cry_13_cZ(.DI(GND),.CI(un1_s_count_4_cry_12),.S(un1_s_count_4_axb_13),.LO(un1_s_count_4_cry_13));
  XORCY un1_s_count_4_s_12_cZ(.LI(un1_s_count_4_axb_12),.CI(un1_s_count_4_cry_11),.O(un1_s_count_4_s_12));
  MUXCY_L un1_s_count_4_cry_12_cZ(.DI(GND),.CI(un1_s_count_4_cry_11),.S(un1_s_count_4_axb_12),.LO(un1_s_count_4_cry_12));
  XORCY un1_s_count_4_s_11_cZ(.LI(un1_s_count_4_axb_11),.CI(un1_s_count_4_cry_10),.O(un1_s_count_4_s_11));
  MUXCY_L un1_s_count_4_cry_11_cZ(.DI(GND),.CI(un1_s_count_4_cry_10),.S(un1_s_count_4_axb_11),.LO(un1_s_count_4_cry_11));
  XORCY un1_s_count_4_s_10_cZ(.LI(un1_s_count_4_axb_10),.CI(un1_s_count_4_cry_9),.O(un1_s_count_4_s_10));
  MUXCY_L un1_s_count_4_cry_10_cZ(.DI(GND),.CI(un1_s_count_4_cry_9),.S(un1_s_count_4_axb_10),.LO(un1_s_count_4_cry_10));
  XORCY un1_s_count_4_s_9_cZ(.LI(un1_s_count_4_axb_9),.CI(un1_s_count_4_cry_8),.O(un1_s_count_4_s_9));
  MUXCY_L un1_s_count_4_cry_9_cZ(.DI(GND),.CI(un1_s_count_4_cry_8),.S(un1_s_count_4_axb_9),.LO(un1_s_count_4_cry_9));
  XORCY un1_s_count_4_s_8_cZ(.LI(un1_s_count_4_axb_8),.CI(un1_s_count_4_cry_7),.O(un1_s_count_4_s_8));
  MUXCY_L un1_s_count_4_cry_8_cZ(.DI(GND),.CI(un1_s_count_4_cry_7),.S(un1_s_count_4_axb_8),.LO(un1_s_count_4_cry_8));
  XORCY un1_s_count_4_s_7_cZ(.LI(un1_s_count_4_axb_7),.CI(un1_s_count_4_cry_6),.O(un1_s_count_4_s_7));
  MUXCY_L un1_s_count_4_cry_7_cZ(.DI(GND),.CI(un1_s_count_4_cry_6),.S(un1_s_count_4_axb_7),.LO(un1_s_count_4_cry_7));
  XORCY un1_s_count_4_s_6_cZ(.LI(un1_s_count_4_axb_6),.CI(un1_s_count_4_cry_5),.O(un1_s_count_4_s_6));
  MUXCY_L un1_s_count_4_cry_6_cZ(.DI(GND),.CI(un1_s_count_4_cry_5),.S(un1_s_count_4_axb_6),.LO(un1_s_count_4_cry_6));
  XORCY un1_s_count_4_s_5_cZ(.LI(un1_s_count_4_axb_5),.CI(un1_s_count_4_cry_4),.O(un1_s_count_4_s_5));
  MUXCY_L un1_s_count_4_cry_5_cZ(.DI(GND),.CI(un1_s_count_4_cry_4),.S(un1_s_count_4_axb_5),.LO(un1_s_count_4_cry_5));
  XORCY un1_s_count_4_s_4_cZ(.LI(un1_s_count_4_axb_4),.CI(un1_s_count_4_cry_3),.O(un1_s_count_4_s_4));
  MUXCY_L un1_s_count_4_cry_4_cZ(.DI(GND),.CI(un1_s_count_4_cry_3),.S(un1_s_count_4_axb_4),.LO(un1_s_count_4_cry_4));
  XORCY un1_s_count_4_s_3_cZ(.LI(un1_s_count_4_axb_3),.CI(un1_s_count_4_cry_2),.O(un1_s_count_4_s_3));
  MUXCY_L un1_s_count_4_cry_3_cZ(.DI(GND),.CI(un1_s_count_4_cry_2),.S(un1_s_count_4_axb_3),.LO(un1_s_count_4_cry_3));
  XORCY un1_s_count_4_s_2_cZ(.LI(un1_s_count_4_axb_2),.CI(un1_s_count_4_cry_1),.O(un1_s_count_4_s_2));
  MUXCY_L un1_s_count_4_cry_2_cZ(.DI(GND),.CI(un1_s_count_4_cry_1),.S(un1_s_count_4_axb_2),.LO(un1_s_count_4_cry_2));
  XORCY un1_s_count_4_s_1_cZ(.LI(un1_s_count_4_axb_1),.CI(un1_s_count_4_cry_0),.O(un1_s_count_4_s_1));
  MUXCY_L un1_s_count_4_cry_1_cZ(.DI(GND),.CI(un1_s_count_4_cry_0),.S(un1_s_count_4_axb_1),.LO(un1_s_count_4_cry_1));
  XORCY un1_s_count_4_s_0_cZ(.LI(un1_s_count_4_axb_0),.CI(un1_s_count_4_cry_0_cy),.O(un1_s_count_4_s_0));
  MUXCY_L un1_s_count_4_cry_0_cZ(.DI(GND),.CI(un1_s_count_4_cry_0_cy),.S(un1_s_count_4_axb_0),.LO(un1_s_count_4_cry_0));
  pre_norm_addsub_inj i_prenorm_addsub(.pre_norm_sqrt_fracta_o_0(pre_norm_sqrt_fracta_o[27:27]),.pre_norm_sqrt_fracta_o_18(pre_norm_sqrt_fracta_o[45:45]),.s_exp_10_o_0(\i_pre_norm_mul.s_exp_10_o_0 [0:0]),.s_exp_10_o(\i_pre_norm_mul.s_exp_10_o [0:0]),.prenorm_addsub_exp_o(prenorm_addsub_exp_o[7:0]),.v_count_56_0_2(\i_prenorm_addsub.v_count_56_0_2 [4:4]),.v_count_1_0_1(\i_pre_norm_div.v_count_1_0_1 ),.v_count_1_0_2(\i_pre_norm_div.v_count_1_0_2 ),.s_opa_i(s_opa_i[30:0]),.s_opb_i(s_opb_i[30:0]),.v_count(\i_pre_norm_sqrt.v_count [4:0]),.v_count_i(\i_pre_norm_sqrt.v_count_i ),.pre_norm_div_dvdnd_8(pre_norm_div_dvdnd[43:43]),.pre_norm_div_dvdnd_9(pre_norm_div_dvdnd[44:44]),.pre_norm_div_dvdnd_0(pre_norm_div_dvdnd[35:35]),.pre_norm_div_dvdnd_4(pre_norm_div_dvdnd[39:39]),.prenorm_addsub_fractb_28_o(prenorm_addsub_fractb_28_o[26:0]),.prenorm_addsub_fracta_28_o(prenorm_addsub_fracta_28_o[26:0]),.s_expa_lt_expb(\i_prenorm_addsub.s_expa_lt_expb ),.N_1084_i(N_1084_i),.N_41(\i_pre_norm_sqrt.s_fracta2_52_o.N_41 ),.N_43(\i_pre_norm_sqrt.s_fracta2_52_o.N_43 ),.N_1628(N_1628),.N_1630(N_1630),.N_1264(N_1264),.N_46(\i_pre_norm_sqrt.s_fracta2_52_o.N_46 ),.N_1236(N_1236),.N_70(\i_pre_norm_div.s_dvdnd_50_o.N_70 ),.N_1624(N_1624),.N_53(\i_pre_norm_sqrt.s_fracta2_52_o.N_53 ),.N_1242(N_1242),.N_1257_i(N_1257_i),.N_1077(N_1077),.N_1083(N_1083),.un2_s_snan_o_20(un2_s_snan_o_20),.N_1051(N_1051),.N_1050(N_1050),.N_987(N_987),.un4_s_expb_in_2_i_0_e(\i_pre_norm_div.un4_s_expb_in_2_i_0_e ),.N_378_i(N_378_i),.N_2103(N_2103),.m46_0_e(\i_prenorm_addsub.m46_0_e ),.clk_i(clk_i),.un4_s_expb_in_2_i_o2_2_lut6_2_O5(un4_s_expb_in_2_i_o2_2_lut6_2_O5),.N_1232_i(N_1232_i),.N_2220(N_2220),.un4_s_expb_in_2_i_o2_2(\i_pre_norm_div.un4_s_expb_in_2_i_o2_2 ),.un4_s_expb_in_2_i_o2_0(\i_pre_norm_div.un4_s_expb_in_2_i_o2_0 ),.un4_s_expb_in_2_i_o2_1(\i_pre_norm_div.un4_s_expb_in_2_i_o2_1 ),.result_1_i_o3(\or_reduce.result_1_i_o3 ),.result_i_o3_lut6_2_O6(\or_reduce.result_i_o3_lut6_2_O6 ),.N_2240(N_2240),.N_399(\i_pre_norm_div.N_399 ),.N_396(\i_pre_norm_div.N_396 ),.N_1227(N_1227),.N_48_0(N_48_0),.N_59(\i_pre_norm_div.s_dvdnd_50_o.N_59 ),.un1_s_infb(un1_s_infb),.result_2_10(\i_postnorm_addsub.or_reduce.result_2_10 ),.un2_s_snan_o_22(un2_s_snan_o_22),.un2_s_snan_o_8(un2_s_snan_o_8),.un4_s_infa_1(\i_prenorm_addsub.un4_s_infa_1 ),.un4_s_infa(un4_s_infa),.N_1041(N_1041),.N_1170(N_1170),.un3_s_snan_o_0(un3_s_snan_o_0),.N_1241(N_1241),.N_30_0(N_30_0),.N_38_0(N_38_0),.N_1617(N_1617),.N_1238(N_1238),.N_27_0(N_27_0),.N_1245(N_1245),.N_143_mux(N_143_mux),.N_1140(N_1140));
  addsub_28_inj i_addsub(.prenorm_addsub_fracta_28_o(prenorm_addsub_fracta_28_o[26:0]),.prenorm_addsub_fractb_28_o(prenorm_addsub_fractb_28_o[26:0]),.s_fpu_op_i(s_fpu_op_i[0:0]),.addsub_fract_o(addsub_fract_o[27:0]),.s_opb_i_26(s_opb_i[31:31]),.s_opb_i_1(s_opb_i[6:6]),.s_opb_i_0(s_opb_i[5:5]),.s_opb_i_2(s_opb_i[7:7]),.s_opa_i_27(s_opa_i[31:31]),.s_opa_i_0(s_opa_i[4:4]),.s_opa_i_1(s_opa_i[5:5]),.N_1941(N_1941),.N_1942_i(N_1942_i),.clk_i(clk_i),.result_2_2(\i_postnorm_addsub.or_reduce.result_2_2 ),.N_1055(N_1055),.un1_s_infb(un1_s_infb),.N_1979(N_1979),.addsub_sign_o(addsub_sign_o),.un2_s_snan_o_8(un2_s_snan_o_8),.N_1166(N_1166),.un4_s_infa(un4_s_infa),.result_3_0_0_i(\i_postnorm_addsub.or_reduce.result_3_0_0_i ),.N_36_0(N_36_0),.result_2(\i_postnorm_addsub.or_reduce.result_2 ),.N_1948(N_1948));
  post_norm_addsub_inj i_postnorm_addsub(.addsub_fract_o(addsub_fract_o[27:0]),.v_count_2_0(\i_pre_norm_div.v_count_2_0 [4:4]),.pre_norm_div_dvsor(pre_norm_div_dvsor[5:5]),.s_opa_i(s_opa_i[31:31]),.s_output_o_0_0(s_output_o_0[22:22]),.s_output_o_0_9(s_output_o_0[31:31]),.postnorm_addsub_output_o(postnorm_addsub_output_o[31:0]),.s_output1(s_output1[31:0]),.s_output_o_1(s_output_o[23:23]),.s_rmode_i(s_rmode_i[1:0]),.s_fpu_op_i(s_fpu_op_i[2:1]),.prenorm_addsub_exp_o(prenorm_addsub_exp_o[7:0]),.s_opb_i_15(s_opb_i[19:19]),.s_opb_i_14(s_opb_i[18:18]),.s_opb_i_2(s_opb_i[6:6]),.s_opb_i_1(s_opb_i[5:5]),.s_opb_i_3(s_opb_i[7:7]),.s_opb_i_17(s_opb_i[21:21]),.s_opb_i_0(s_opb_i[4:4]),.s_opb_i_16(s_opb_i[20:20]),.s_opb_i_18(s_opb_i[22:22]),.s_opb_i_27(s_opb_i[31:31]),.un4_s_infa(un4_s_infa),.un1_s_infb(un1_s_infb),.div_zero_o_0(div_zero_o_0),.un3_s_snan_o_0(un3_s_snan_o_0),.N_9_i_0_e(\i_postnorm_addsub.N_9_i_0_e ),.N_54(\i_pre_norm_div.s_dvsor_27_o.N_54 ),.result_2_10(\i_postnorm_addsub.or_reduce.result_2_10 ),.result_i_0_0(\or_reduce.result_i_0_0 ),.s_ine_o(s_ine_o),.un2_s_qnan_o_0_a2_0_e(\i_postnorm_addsub.un2_s_qnan_o_0_a2_0_e ),.N_6_i_0_e(\i_postnorm_addsub.N_6_i_0_e ),.clk_i(clk_i),.N_765_i_0_e(\i_postnorm_addsub.N_765_i_0_e ),.N_763_i_0_e(\i_postnorm_addsub.N_763_i_0_e ),.N_12_i_0_e(\i_postnorm_addsub.N_12_i_0_e ),.N_773_i_0_e(\i_postnorm_addsub.N_773_i_0_e ),.N_1941(N_1941),.un3_s_underflow_o_0(un3_s_underflow_o_0),.postnorm_addsub_ine_o(postnorm_addsub_ine_o),.result_2_2(\i_postnorm_addsub.or_reduce.result_2_2 ),.N_1055(N_1055),.result_2(\i_postnorm_addsub.or_reduce.result_2 ),.result_2_16(\i_postnorm_addsub.or_reduce.result_2_16 ),.N_1051(N_1051),.N_764_i(N_764_i),.N_766_i(N_766_i),.N_767_i(N_767_i),.N_768_i(N_768_i),.N_769_i(N_769_i),.N_770_i(N_770_i),.N_771_i(N_771_i),.N_772_i(N_772_i),.N_774_i(N_774_i),.N_775_i(N_775_i),.N_776_i(N_776_i),.N_777_i(N_777_i),.N_778_i(N_778_i),.N_779_i(N_779_i),.N_780_i(N_780_i),.N_14_i(N_14_i),.N_18_i(N_18_i),.N_20_i(N_20_i),.addsub_sign_o(addsub_sign_o),.N_1979(N_1979),.N_36_0(N_36_0),.N_1948(N_1948));
  pre_norm_mul_inj i_pre_norm_mul(.v_count(\i_pre_norm_sqrt.v_count [4:4]),.s_fracta_52_o_0_e(\i_pre_norm_sqrt.s_fracta_52_o_0_e [29:29]),.pre_norm_mul_exp_10(pre_norm_mul_exp_10[9:0]),.s_exp_10_o_1(\i_pre_norm_mul.s_exp_10_o [1:1]),.s_exp_10_o_0_d0(\i_pre_norm_mul.s_exp_10_o [0:0]),.s_exp_10_o_0_0(\i_pre_norm_mul.s_exp_10_o_0 [0:0]),.s_exp_10_o_0_1(\i_pre_norm_mul.s_exp_10_o_0 [1:1]),.s_opb_i(s_opb_i[30:23]),.s_opa_i(s_opa_i[30:23]),.un4_s_expb_in_2_i_o2_0(\i_pre_norm_div.un4_s_expb_in_2_i_o2_0 ),.N_48_0(N_48_0),.N_1245(N_1245),.clk_i(clk_i),.un4_s_expb_in_2_i_o2_1(\i_pre_norm_div.un4_s_expb_in_2_i_o2_1 ),.N_1077(N_1077),.result_i_o3_lut6_2_O6(\or_reduce.result_i_o3_lut6_2_O6 ),.N_1084_i(N_1084_i),.p_desc595_p_O_FD(p_desc595_p_O_FDpre_norm_mul_),.p_desc596_p_O_FD(p_desc596_p_O_FDpre_norm_mul_),.p_desc597_p_O_FD(p_desc597_p_O_FDpre_norm_mul_),.p_desc598_p_O_FD(p_desc598_p_O_FDpre_norm_mul_),.p_desc599_p_O_FD(p_desc599_p_O_FDpre_norm_mul_),.p_desc600_p_O_FD(p_desc600_p_O_FDpre_norm_mul_),.p_desc601_p_O_FD(p_desc601_p_O_FDpre_norm_mul_),.p_desc602_p_O_FD(p_desc602_p_O_FDpre_norm_mul_),.p_desc603_p_O_FD(p_desc603_p_O_FDpre_norm_mul_),.p_desc604_p_O_FD(p_desc604_p_O_FDpre_norm_mul_));
  mul_24_inj i_mul_24(.s_fractb_i_11(\i_mul_24.s_fractb_i [11:11]),.s_fractb_i_8(\i_mul_24.s_fractb_i [8:8]),.s_fractb_i_20(\i_mul_24.s_fractb_i [20:20]),.s_fractb_i_10(\i_mul_24.s_fractb_i [10:10]),.s_fractb_i_9(\i_mul_24.s_fractb_i [9:9]),.s_fractb_i_22(\i_mul_24.s_fractb_i [22:22]),.s_fractb_i_21(\i_mul_24.s_fractb_i [21:21]),.s_fractb_i_7(\i_mul_24.s_fractb_i [7:7]),.s_fractb_i_6(\i_mul_24.s_fractb_i [6:6]),.s_fractb_i_19(\i_mul_24.s_fractb_i [19:19]),.s_fractb_i_18(\i_mul_24.s_fractb_i [18:18]),.s_fractb_i_5(\i_mul_24.s_fractb_i [5:5]),.s_fractb_i_4(\i_mul_24.s_fractb_i [4:4]),.s_fractb_i_17(\i_mul_24.s_fractb_i [17:17]),.s_fractb_i_16(\i_mul_24.s_fractb_i [16:16]),.s_fractb_i_3(\i_mul_24.s_fractb_i [3:3]),.s_fractb_i_15(\i_mul_24.s_fractb_i [15:15]),.s_fractb_i_2(\i_mul_24.s_fractb_i [2:2]),.s_fractb_i_14(\i_mul_24.s_fractb_i [14:14]),.s_fractb_i_1(\i_mul_24.s_fractb_i [1:1]),.s_fractb_i_13(\i_mul_24.s_fractb_i [13:13]),.s_fractb_i_0(\i_mul_24.s_fractb_i [0:0]),.s_fractb_i_12(\i_mul_24.s_fractb_i [12:12]),.s_fracta_i(\i_mul_24.s_fracta_i [22:0]),.s_opb_i_31(s_opb_i[31:31]),.s_opb_i_11(s_opb_i[11:11]),.s_opb_i_10(s_opb_i[10:10]),.s_opb_i_22(s_opb_i[22:22]),.s_opb_i_9(s_opb_i[9:9]),.s_opb_i_21(s_opb_i[21:21]),.s_opb_i_8(s_opb_i[8:8]),.s_opb_i_20(s_opb_i[20:20]),.s_opb_i_7(s_opb_i[7:7]),.s_opb_i_19(s_opb_i[19:19]),.s_opb_i_6(s_opb_i[6:6]),.s_opb_i_18(s_opb_i[18:18]),.s_opb_i_5(s_opb_i[5:5]),.s_opb_i_17(s_opb_i[17:17]),.s_opb_i_4(s_opb_i[4:4]),.s_opb_i_16(s_opb_i[16:16]),.s_opb_i_3(s_opb_i[3:3]),.s_opb_i_15(s_opb_i[15:15]),.s_opb_i_2(s_opb_i[2:2]),.s_opb_i_14(s_opb_i[14:14]),.s_opb_i_1(s_opb_i[1:1]),.s_opb_i_13(s_opb_i[13:13]),.s_opb_i_0(s_opb_i[0:0]),.s_opb_i_12(s_opb_i[12:12]),.s_opa_i_31(s_opa_i[31:31]),.s_opa_i_11(s_opa_i[11:11]),.s_opa_i_10(s_opa_i[10:10]),.s_opa_i_22(s_opa_i[22:22]),.s_opa_i_9(s_opa_i[9:9]),.s_opa_i_21(s_opa_i[21:21]),.s_opa_i_8(s_opa_i[8:8]),.s_opa_i_20(s_opa_i[20:20]),.s_opa_i_7(s_opa_i[7:7]),.s_opa_i_19(s_opa_i[19:19]),.s_opa_i_6(s_opa_i[6:6]),.s_opa_i_18(s_opa_i[18:18]),.s_opa_i_5(s_opa_i[5:5]),.s_opa_i_17(s_opa_i[17:17]),.s_opa_i_4(s_opa_i[4:4]),.s_opa_i_16(s_opa_i[16:16]),.s_opa_i_3(s_opa_i[3:3]),.s_opa_i_15(s_opa_i[15:15]),.s_opa_i_2(s_opa_i[2:2]),.s_opa_i_14(s_opa_i[14:14]),.s_opa_i_1(s_opa_i[1:1]),.s_opa_i_13(s_opa_i[13:13]),.s_opa_i_0(s_opa_i[0:0]),.s_opa_i_12(s_opa_i[12:12]),.mul_24_fract_48(mul_24_fract_48[47:0]),.opa_i(opa_i[17:12]),.opb_i(opb_i[17:12]),.clk_i(clk_i),.s_start_i(s_start_i),.result_1_i_o3_0_e(\i_pre_norm_div.or_reduce.result_1_i_o3_0_e ),.s_signa_i(\i_mul_24.s_signa_i ),.s_signb_i(\i_mul_24.s_signb_i ),.result_i_o3_lut6_2_O6(\or_reduce.result_i_o3_lut6_2_O6 ));
  post_norm_mul_inj i_post_norm_mul(.pre_norm_mul_exp_10(pre_norm_mul_exp_10[9:0]),.mul_24_fract_48(mul_24_fract_48[47:0]),.s_fracta_i_20(\i_mul_24.s_fracta_i [20:20]),.s_fracta_i_21(\i_mul_24.s_fracta_i [21:21]),.s_fracta_i_0(\i_mul_24.s_fracta_i [0:0]),.s_fracta_i_1(\i_mul_24.s_fracta_i [1:1]),.s_fracta_i_2(\i_mul_24.s_fracta_i [2:2]),.s_fracta_i_3(\i_mul_24.s_fracta_i [3:3]),.s_fracta_i_4(\i_mul_24.s_fracta_i [4:4]),.s_fracta_i_5(\i_mul_24.s_fracta_i [5:5]),.s_fracta_i_6(\i_mul_24.s_fracta_i [6:6]),.s_fracta_i_7(\i_mul_24.s_fracta_i [7:7]),.s_fracta_i_8(\i_mul_24.s_fracta_i [8:8]),.s_fracta_i_9(\i_mul_24.s_fracta_i [9:9]),.s_fracta_i_10(\i_mul_24.s_fracta_i [10:10]),.s_fracta_i_11(\i_mul_24.s_fracta_i [11:11]),.s_fracta_i_12(\i_mul_24.s_fracta_i [12:12]),.s_fracta_i_13(\i_mul_24.s_fracta_i [13:13]),.s_fracta_i_14(\i_mul_24.s_fracta_i [14:14]),.s_fracta_i_15(\i_mul_24.s_fracta_i [15:15]),.s_rmode_i(\i_post_norm_mul.s_rmode_i [1:0]),.post_norm_mul_output(post_norm_mul_output[31:0]),.clk_i(clk_i),.N_6_i(N_6_i),.post_norm_mul_ine(post_norm_mul_ine),.s_infb(\i_post_norm_mul.s_infb ),.un1_s_infa(\i_post_norm_mul.un1_s_infa ),.result_5(\i_post_norm_mul.or_reduce.result_5 ),.un1_s_nan_b(\i_post_norm_mul.un1_s_nan_b ),.result_4(\i_post_norm_mul.or_reduce.result_4 ),.un1_s_nan_a(\i_post_norm_mul.un1_s_nan_a ),.un3_s_op_0(\i_post_norm_mul.un3_s_op_0 ),.result_11(\i_post_norm_sqrt.or_reduce.result_11 ),.result_3_21_1(\i_post_norm_mul.or_reduce.result_3_21_1 ),.result_3_21_3(\i_post_norm_mul.or_reduce.result_3_21_3 ),.p_desc1070_p_O_FD(p_desc1070_p_O_FDpost_norm_mul_),.p_desc1071_p_O_FD(p_desc1071_p_O_FDpost_norm_mul_),.p_desc1072_p_O_FD(p_desc1072_p_O_FDpost_norm_mul_),.p_desc1073_p_O_FD(p_desc1073_p_O_FDpost_norm_mul_),.p_desc1074_p_O_FD(p_desc1074_p_O_FDpost_norm_mul_),.p_desc1075_p_O_FD(p_desc1075_p_O_FDpost_norm_mul_),.p_desc1076_p_O_FD(p_desc1076_p_O_FDpost_norm_mul_),.p_desc1077_p_O_FD(p_desc1077_p_O_FDpost_norm_mul_),.p_desc1078_p_O_FD(p_desc1078_p_O_FDpost_norm_mul_),.p_desc1079_p_O_FD(p_desc1079_p_O_FDpost_norm_mul_),.p_desc1080_p_O_FD(p_desc1080_p_O_FDpost_norm_mul_),.p_desc1081_p_O_FD(p_desc1081_p_O_FDpost_norm_mul_),.p_desc1082_p_O_FD(p_desc1082_p_O_FDpost_norm_mul_),.p_desc1083_p_O_FD(p_desc1083_p_O_FDpost_norm_mul_),.p_desc1084_p_O_FD(p_desc1084_p_O_FDpost_norm_mul_),.p_desc1085_p_O_FD(p_desc1085_p_O_FDpost_norm_mul_),.p_desc1086_p_O_FD(p_desc1086_p_O_FDpost_norm_mul_),.p_desc1087_p_O_FD(p_desc1087_p_O_FDpost_norm_mul_),.p_desc1088_p_O_FD(p_desc1088_p_O_FDpost_norm_mul_),.p_desc1089_p_O_FD(p_desc1089_p_O_FDpost_norm_mul_),.p_desc1090_p_O_FD(p_desc1090_p_O_FDpost_norm_mul_),.p_desc1091_p_O_FD(p_desc1091_p_O_FDpost_norm_mul_),.p_desc1092_p_O_FD(p_desc1092_p_O_FDpost_norm_mul_),.p_desc1163_p_O_FD(p_desc1163_p_O_FDpost_norm_mul_),.p_desc1164_p_O_FD(p_desc1164_p_O_FDpost_norm_mul_),.p_desc1165_p_O_FD(p_desc1165_p_O_FDpost_norm_mul_),.p_desc1166_p_O_FD(p_desc1166_p_O_FDpost_norm_mul_),.p_desc1167_p_O_FD(p_desc1167_p_O_FDpost_norm_mul_),.p_desc1168_p_O_FD(p_desc1168_p_O_FDpost_norm_mul_),.p_desc1169_p_O_FD(p_desc1169_p_O_FDpost_norm_mul_),.p_desc1170_p_O_FD(p_desc1170_p_O_FDpost_norm_mul_),.p_desc1171_p_O_FD(p_desc1171_p_O_FDpost_norm_mul_),.p_desc1172_p_O_FD(p_desc1172_p_O_FDpost_norm_mul_),.p_desc1173_p_O_FD(p_desc1173_p_O_FDpost_norm_mul_),.p_desc1174_p_O_FD(p_desc1174_p_O_FDpost_norm_mul_),.p_desc1175_p_O_FD(p_desc1175_p_O_FDpost_norm_mul_),.p_desc1176_p_O_FD(p_desc1176_p_O_FDpost_norm_mul_),.p_desc1177_p_O_FD(p_desc1177_p_O_FDpost_norm_mul_),.p_desc1178_p_O_FD(p_desc1178_p_O_FDpost_norm_mul_),.p_desc1179_p_O_FD(p_desc1179_p_O_FDpost_norm_mul_),.p_desc1180_p_O_FD(p_desc1180_p_O_FDpost_norm_mul_),.p_desc1181_p_O_FD(p_desc1181_p_O_FDpost_norm_mul_),.p_desc1182_p_O_FD(p_desc1182_p_O_FDpost_norm_mul_),.p_desc1183_p_O_FD(p_desc1183_p_O_FDpost_norm_mul_),.p_desc1184_p_O_FD(p_desc1184_p_O_FDpost_norm_mul_),.p_desc1185_p_O_FD(p_desc1185_p_O_FDpost_norm_mul_),.p_desc1186_p_O_FD(p_desc1186_p_O_FDpost_norm_mul_),.p_desc1187_p_O_FD(p_desc1187_p_O_FDpost_norm_mul_),.p_desc1188_p_O_FD(p_desc1188_p_O_FDpost_norm_mul_),.p_desc1189_p_O_FD(p_desc1189_p_O_FDpost_norm_mul_),.p_desc1190_p_O_FD(p_desc1190_p_O_FDpost_norm_mul_),.p_desc1191_p_O_FD(p_desc1191_p_O_FDpost_norm_mul_),.p_desc1192_p_O_FD(p_desc1192_p_O_FDpost_norm_mul_),.p_desc1193_p_O_FD(p_desc1193_p_O_FDpost_norm_mul_),.p_desc1194_p_O_FD(p_desc1194_p_O_FDpost_norm_mul_),.p_desc1195_p_O_FD(p_desc1195_p_O_FDpost_norm_mul_),.p_desc1196_p_O_FD(p_desc1196_p_O_FDpost_norm_mul_),.p_desc1197_p_O_FD(p_desc1197_p_O_FDpost_norm_mul_),.p_desc1198_p_O_FD(p_desc1198_p_O_FDpost_norm_mul_),.p_desc1199_p_O_FD(p_desc1199_p_O_FDpost_norm_mul_),.p_desc1200_p_O_FD(p_desc1200_p_O_FDpost_norm_mul_),.p_desc1201_p_O_FD(p_desc1201_p_O_FDpost_norm_mul_),.p_desc1202_p_O_FD(p_desc1202_p_O_FDpost_norm_mul_),.p_desc1203_p_O_FD(p_desc1203_p_O_FDpost_norm_mul_),.p_desc1204_p_O_FD(p_desc1204_p_O_FDpost_norm_mul_),.p_desc1205_p_O_FD(p_desc1205_p_O_FDpost_norm_mul_),.p_desc1206_p_O_FD(p_desc1206_p_O_FDpost_norm_mul_),.p_desc1207_p_O_FD(p_desc1207_p_O_FDpost_norm_mul_),.p_desc1208_p_O_FD(p_desc1208_p_O_FDpost_norm_mul_),.p_desc1209_p_O_FD(p_desc1209_p_O_FDpost_norm_mul_),.p_desc1210_p_O_FD(p_desc1210_p_O_FDpost_norm_mul_),.p_desc1211_p_O_FD(p_desc1211_p_O_FDpost_norm_mul_),.p_desc1212_p_O_FD(p_desc1212_p_O_FDpost_norm_mul_),.p_desc1213_p_O_FD(p_desc1213_p_O_FDpost_norm_mul_),.p_desc1214_p_O_FD(p_desc1214_p_O_FDpost_norm_mul_),.p_desc1215_p_O_FD(p_desc1215_p_O_FDpost_norm_mul_),.p_desc1216_p_O_FD(p_desc1216_p_O_FDpost_norm_mul_),.p_desc1217_p_O_FD(p_desc1217_p_O_FDpost_norm_mul_),.p_desc1218_p_O_FD(p_desc1218_p_O_FDpost_norm_mul_),.p_desc1219_p_O_FD(p_desc1219_p_O_FDpost_norm_mul_),.p_desc1220_p_O_FD(p_desc1220_p_O_FDpost_norm_mul_),.p_desc1221_p_O_FD(p_desc1221_p_O_FDpost_norm_mul_),.p_s_sign_i_Z_p_O_FD(p_s_sign_i_Z_p_O_FDpost_norm_mul_),.p_ine_o_Z_p_O_FD(p_ine_o_Z_p_O_FDpost_norm_mul_),.p_desc1244_p_O_FD(p_desc1244_p_O_FDpost_norm_mul_),.p_desc1245_p_O_FD(p_desc1245_p_O_FDpost_norm_mul_),.p_desc1246_p_O_FD(p_desc1246_p_O_FDpost_norm_mul_),.p_desc1247_p_O_FD(p_desc1247_p_O_FDpost_norm_mul_),.p_desc1248_p_O_FD(p_desc1248_p_O_FDpost_norm_mul_),.p_desc1249_p_O_FD(p_desc1249_p_O_FDpost_norm_mul_),.p_desc1250_p_O_FD(p_desc1250_p_O_FDpost_norm_mul_),.p_desc1251_p_O_FD(p_desc1251_p_O_FDpost_norm_mul_),.p_desc1252_p_O_FD(p_desc1252_p_O_FDpost_norm_mul_),.p_desc1253_p_O_FD(p_desc1253_p_O_FDpost_norm_mul_),.p_desc1254_p_O_FD(p_desc1254_p_O_FDpost_norm_mul_),.p_desc1255_p_O_FD(p_desc1255_p_O_FDpost_norm_mul_),.p_desc1256_p_O_FD(p_desc1256_p_O_FDpost_norm_mul_),.p_desc1257_p_O_FD(p_desc1257_p_O_FDpost_norm_mul_),.p_desc1258_p_O_FD(p_desc1258_p_O_FDpost_norm_mul_),.p_desc1259_p_O_FD(p_desc1259_p_O_FDpost_norm_mul_),.p_desc1260_p_O_FD(p_desc1260_p_O_FDpost_norm_mul_),.p_desc1261_p_O_FD(p_desc1261_p_O_FDpost_norm_mul_),.p_desc1262_p_O_FD(p_desc1262_p_O_FDpost_norm_mul_),.p_desc1263_p_O_FD(p_desc1263_p_O_FDpost_norm_mul_),.p_desc1264_p_O_FD(p_desc1264_p_O_FDpost_norm_mul_),.p_desc1265_p_O_FD(p_desc1265_p_O_FDpost_norm_mul_),.p_desc1266_p_O_FD(p_desc1266_p_O_FDpost_norm_mul_),.p_desc1267_p_O_FD(p_desc1267_p_O_FDpost_norm_mul_),.p_desc1268_p_O_FD(p_desc1268_p_O_FDpost_norm_mul_),.p_desc1269_p_O_FD(p_desc1269_p_O_FDpost_norm_mul_),.p_desc1270_p_O_FD(p_desc1270_p_O_FDpost_norm_mul_),.p_desc1271_p_O_FD(p_desc1271_p_O_FDpost_norm_mul_),.p_desc1272_p_O_FD(p_desc1272_p_O_FDpost_norm_mul_),.p_desc1273_p_O_FD(p_desc1273_p_O_FDpost_norm_mul_),.p_desc1274_p_O_FD(p_desc1274_p_O_FDpost_norm_mul_),.p_desc1275_p_O_FD(p_desc1275_p_O_FDpost_norm_mul_),.p_desc1276_p_O_FD(p_desc1276_p_O_FDpost_norm_mul_),.p_desc1277_p_O_FD(p_desc1277_p_O_FDpost_norm_mul_),.p_desc1278_p_O_FD(p_desc1278_p_O_FDpost_norm_mul_),.p_desc1279_p_O_FD(p_desc1279_p_O_FDpost_norm_mul_),.p_desc1280_p_O_FD(p_desc1280_p_O_FDpost_norm_mul_),.p_desc1281_p_O_FD(p_desc1281_p_O_FDpost_norm_mul_),.p_desc1282_p_O_FD(p_desc1282_p_O_FDpost_norm_mul_),.p_desc1283_p_O_FD(p_desc1283_p_O_FDpost_norm_mul_),.p_desc1284_p_O_FD(p_desc1284_p_O_FDpost_norm_mul_),.p_desc1285_p_O_FD(p_desc1285_p_O_FDpost_norm_mul_),.p_desc1286_p_O_FD(p_desc1286_p_O_FDpost_norm_mul_),.p_desc1287_p_O_FD(p_desc1287_p_O_FDpost_norm_mul_),.p_desc1288_p_O_FD(p_desc1288_p_O_FDpost_norm_mul_),.p_desc1289_p_O_FD(p_desc1289_p_O_FDpost_norm_mul_),.p_desc1290_p_O_FD(p_desc1290_p_O_FDpost_norm_mul_),.p_desc1291_p_O_FD(p_desc1291_p_O_FDpost_norm_mul_));
  pre_norm_div_inj i_pre_norm_div(.v_count_3(\i_pre_norm_sqrt.v_count [3:3]),.v_count_2(\i_pre_norm_sqrt.v_count [2:2]),.v_count_1_0_0_a2_0(\i_pre_norm_div.v_count_1_0_0_a2_0 [1:1]),.v_count_2_0(\i_pre_norm_div.v_count_2_0 [4:4]),.s_exp_10_o_0(\i_pre_norm_mul.s_exp_10_o_0 [1:0]),.s_exp_10_o(\i_pre_norm_mul.s_exp_10_o [1:1]),.pre_norm_div_dvsor_0(pre_norm_div_dvsor_0[23:23]),.v_count_1_0_1(\i_pre_norm_div.v_count_1_0_1 ),.v_count_1_0_2(\i_pre_norm_div.v_count_1_0_2 ),.v_count_0_4(\i_pre_norm_sqrt.v_count [4:4]),.v_count_0_1(\i_pre_norm_sqrt.v_count [1:1]),.v_count_0_0(\i_pre_norm_sqrt.v_count [0:0]),.v_count_i(\i_pre_norm_sqrt.v_count_i ),.s_opb_i({\i_post_norm_mul.s_opb_i [30:29],s_opb_i[28:27],\i_post_norm_mul.s_opb_i [26:25],s_opb_i[24:0]}),.s_opb_i_0_0(\i_post_norm_mul.s_opb_i [24:24]),.s_opb_i_0_3(\i_post_norm_mul.s_opb_i [27:27]),.s_opb_i_0_4(\i_post_norm_mul.s_opb_i [28:28]),.s_opb_i_0_2(s_opb_i[26:26]),.s_opb_i_0_5(s_opb_i[29:29]),.s_opa_i_0({\i_post_norm_mul.s_opa_i [30:30],s_opa_i[29:28],\i_post_norm_mul.s_opa_i [27:26],s_opa_i[25:25],\i_post_norm_mul.s_opa_i [24:24]}),.s_opa_i({s_opa_i[30:30],\i_post_norm_mul.s_opa_i [29:28],s_opa_i[27:26],\i_post_norm_mul.s_opa_i [25:25],s_opa_i[24:0]}),.v_count_1_0_a2_7_i_0(\i_pre_norm_div.v_count_1_0_a2_7_i_0 ),.pre_norm_div_dvsor(pre_norm_div_dvsor[22:7]),.pre_norm_div_dvdnd_0(pre_norm_div_dvdnd[36:36]),.pre_norm_div_dvdnd_11(pre_norm_div_dvdnd[47:47]),.un11_s_exp_10_o_0(\i_pre_norm_div.un11_s_exp_10_o_0 [9:1]),.N_1083(N_1083),.N_143_mux(N_143_mux),.N_48_0(N_48_0),.N_59(\i_pre_norm_div.s_dvdnd_50_o.N_59 ),.N_54(\i_pre_norm_div.s_dvsor_27_o.N_54 ),.N_1630(N_1630),.N_55(\i_pre_norm_div.s_dvdnd_50_o.N_55 ),.N_63(\i_pre_norm_div.s_dvdnd_50_o.N_63 ),.N_1278_i(N_1278_i),.s_dvdnd_50_o_105_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_105_0_e ),.N_987(N_987),.s_expa_lt_expb(\i_prenorm_addsub.s_expa_lt_expb ),.N_2240(N_2240),.N_1232_i(N_1232_i),.un2_s_snan_o_22(un2_s_snan_o_22),.N_1174(N_1174),.result_i_o3_lut6_2_O6(\or_reduce.result_i_o3_lut6_2_O6 ),.result_3_0_0_i(\i_postnorm_addsub.or_reduce.result_3_0_0_i ),.N_1055(N_1055),.N_1077(N_1077),.N_399(\i_pre_norm_div.N_399 ),.un4_s_infa_1(\i_prenorm_addsub.un4_s_infa_1 ),.N_1140(N_1140),.N_1051(N_1051),.N_2220(N_2220),.N_1170(N_1170),.un4_s_expb_in_2_i_o2_2(\i_pre_norm_div.un4_s_expb_in_2_i_o2_2 ),.un4_s_expb_in_2_i_o2_2_lut6_2_O5(un4_s_expb_in_2_i_o2_2_lut6_2_O5),.N_1041(N_1041),.result_2_16(\i_postnorm_addsub.or_reduce.result_2_16 ),.s_dvdnd_50_o_104_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_104_0_e ),.un4_s_expb_in_2_i_0_e(\i_pre_norm_div.un4_s_expb_in_2_i_0_e ),.clk_i(clk_i),.s_dvdnd_50_o_103_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_103_0_e ),.s_dvdnd_50_o_102_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_102_0_e ),.s_dvdnd_50_o_106_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_106_0_e ),.s_dvdnd_50_o_108_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_108_0_e ),.N_1236(N_1236),.N_2103(N_2103),.s_dvdnd_50_o_107_0_e(\i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_107_0_e ),.un4_s_expb_in_2_i_o2_0(\i_pre_norm_div.un4_s_expb_in_2_i_o2_0 ),.un4_s_expb_in_2_i_o2_1(\i_pre_norm_div.un4_s_expb_in_2_i_o2_1 ),.result_1_i_o3_0_e(\i_pre_norm_div.or_reduce.result_1_i_o3_0_e ),.N_1227(N_1227),.N_378_i(N_378_i),.N_396(\i_pre_norm_div.N_396 ),.result_1_i_o3(\or_reduce.result_1_i_o3 ),.N_1084_i(N_1084_i),.un11_s_exp_10_o_axb_0_i(\i_pre_norm_div.un11_s_exp_10_o_axb_0_i ),.N_1050(N_1050),.N_1087(N_1087),.un2_s_snan_o_8(un2_s_snan_o_8),.result_2_10(\i_postnorm_addsub.or_reduce.result_2_10 ),.N_1617(N_1617),.N_41_0(\i_pre_norm_sqrt.s_fracta2_52_o.N_41 ),.N_43_0(\i_pre_norm_sqrt.s_fracta2_52_o.N_43 ),.N_44(\i_pre_norm_sqrt.s_fracta2_52_o.N_44 ),.N_45_0(\i_pre_norm_sqrt.s_fracta2_52_o.N_45 ),.N_1628(N_1628),.N_1624(N_1624),.N_1619(N_1619),.N_46(\i_pre_norm_sqrt.s_fracta2_52_o.N_46 ),.N_1620(N_1620),.N_95_0(\i_pre_norm_div.s_dvdnd_50_o.N_95 ),.N_70_0(\i_pre_norm_div.s_dvdnd_50_o.N_70 ),.N_27_0(N_27_0),.N_1238(N_1238));
  serial_div_inj i_serial_div(.fpu_op_i(fpu_op_i[2:0]),.s_state(\i_serial_div.s_state ),.pre_norm_div_dvdnd_0(pre_norm_div_dvdnd_0[49:49]),.pre_norm_div_dvdnd_8(pre_norm_div_dvdnd[42:42]),.pre_norm_div_dvdnd_9(pre_norm_div_dvdnd[43:43]),.pre_norm_div_dvdnd_10(pre_norm_div_dvdnd[44:44]),.pre_norm_div_dvdnd_11(pre_norm_div_dvdnd[45:45]),.pre_norm_div_dvdnd_12(pre_norm_div_dvdnd[46:46]),.pre_norm_div_dvdnd_13(pre_norm_div_dvdnd[47:47]),.pre_norm_div_dvdnd_14(pre_norm_div_dvdnd[48:48]),.pre_norm_div_dvdnd_0_d0(pre_norm_div_dvdnd[34:34]),.pre_norm_div_dvdnd_1(pre_norm_div_dvdnd[35:35]),.pre_norm_div_dvdnd_2(pre_norm_div_dvdnd[36:36]),.pre_norm_div_dvdnd_3(pre_norm_div_dvdnd[37:37]),.pre_norm_div_dvdnd_5(pre_norm_div_dvdnd[39:39]),.pre_norm_div_dvsor_0(pre_norm_div_dvsor_0[23:23]),.pre_norm_div_dvsor_5(pre_norm_div_dvsor[10:10]),.pre_norm_div_dvsor_6(pre_norm_div_dvsor[11:11]),.pre_norm_div_dvsor_7(pre_norm_div_dvsor[12:12]),.pre_norm_div_dvsor_8(pre_norm_div_dvsor[13:13]),.pre_norm_div_dvsor_9(pre_norm_div_dvsor[14:14]),.pre_norm_div_dvsor_10(pre_norm_div_dvsor[15:15]),.pre_norm_div_dvsor_11(pre_norm_div_dvsor[16:16]),.pre_norm_div_dvsor_12(pre_norm_div_dvsor[17:17]),.pre_norm_div_dvsor_13(pre_norm_div_dvsor[18:18]),.pre_norm_div_dvsor_14(pre_norm_div_dvsor[19:19]),.pre_norm_div_dvsor_15(pre_norm_div_dvsor[20:20]),.pre_norm_div_dvsor_16(pre_norm_div_dvsor[21:21]),.pre_norm_div_dvsor_17(pre_norm_div_dvsor[22:22]),.pre_norm_div_dvsor_0_d0(pre_norm_div_dvsor[5:5]),.pre_norm_div_dvsor_2(pre_norm_div_dvsor[7:7]),.pre_norm_div_dvsor_3(pre_norm_div_dvsor[8:8]),.pre_norm_div_dvsor_4(pre_norm_div_dvsor[9:9]),.post_norm_sqrt_output(post_norm_sqrt_output[31:0]),.postnorm_addsub_output_o(postnorm_addsub_output_o[31:0]),.s_output1_6_2_i_m2(s_output1_6_2_i_m2[7:6]),.post_norm_div_output(post_norm_div_output[31:0]),.post_norm_mul_output(post_norm_mul_output[31:0]),.serial_div_qutnt(serial_div_qutnt[26:0]),.serial_div_rmndr(serial_div_rmndr[26:0]),.N_2637_i(N_2637_i),.s_dvdnd_50_o_108_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_108_0_e ),.clk_i(clk_i),.s_dvdnd_50_o_104_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_104_0_e ),.s_dvdnd_50_o_106_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_106_0_e ),.s_dvdnd_50_o_107_0_e(\i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_107_0_e ),.s_dvdnd_50_o_108_0_e_0(\i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_108_0_e ),.s_dvdnd_50_o_106_0_e_0(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_106_0_e ),.m49_0_e(\i_prenorm_addsub.m49_0_e ),.s_dvdnd_50_o_105_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_105_0_e ),.s_dvdnd_50_o_102_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_102_0_e ),.m46_0_e(\i_prenorm_addsub.m46_0_e ),.s_dvdnd_50_o_105_0_e_0(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_105_0_e ),.s_dvdnd_50_o_109_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_109_0_e ),.s_dvdnd_50_o_102_0_e_0(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_102_0_e ),.s_dvdnd_50_o_103_0_e(\i_pre_norm_div.s_dvsor_27_o.s_dvdnd_50_o_103_0_e ),.s_start_i(\i_sqrt.s_start_i ),.div_zero_o_0_0(div_zero_o_0_0),.N_1257_i(N_1257_i),.N_1278_i(N_1278_i),.N_88(\i_pre_norm_sqrt.s_fracta2_52_o.N_88 ),.un12_s_state_0_a2_lut6_2_O5(un12_s_state_0_a2_lut6_2_O5),.post_norm_div_ine(post_norm_div_ine),.post_norm_mul_ine(post_norm_mul_ine),.N_564(N_564),.N_563(N_563),.N_562(N_562),.N_561(N_561),.N_560(N_560),.N_559(N_559),.N_558(N_558),.N_557(N_557),.N_556(N_556),.N_555(N_555),.N_554(N_554),.N_553(N_553),.N_552(N_552),.N_551(N_551),.N_550(N_550),.N_549(N_549),.N_548(N_548),.N_547(N_547),.N_546(N_546),.N_545(N_545),.N_544(N_544),.N_543(N_543),.N_542(N_542),.N_541(N_541),.N_538(N_538),.N_537(N_537),.N_536(N_536),.N_503_i(N_503_i),.N_502_i(N_502_i),.N_501_i(N_501_i),.post_norm_sqrt_ine_o(post_norm_sqrt_ine_o),.postnorm_addsub_ine_o(postnorm_addsub_ine_o),.s_ine_o_5(s_ine_o_5),.div_zero_o_0(div_zero_o_0));
  post_norm_div_inj i_post_norm_div(.un11_s_exp_10_o_0(\i_pre_norm_div.un11_s_exp_10_o_0 [9:1]),.s_opb_i_4(\i_post_norm_mul.s_opb_i [27:27]),.s_opb_i_5(\i_post_norm_mul.s_opb_i [28:28]),.s_opb_i_6(\i_post_norm_mul.s_opb_i [29:29]),.s_opb_i_7(\i_post_norm_mul.s_opb_i [30:30]),.s_opb_i_1(\i_post_norm_mul.s_opb_i [24:24]),.s_opb_i_2(\i_post_norm_mul.s_opb_i [25:25]),.s_opb_i_3(\i_post_norm_mul.s_opb_i [26:26]),.s_opb_i_0(s_opb_i[30:23]),.s_opa_i_1(\i_post_norm_mul.s_opa_i [24:24]),.s_opa_i_2(\i_post_norm_mul.s_opa_i [25:25]),.s_opa_i_3(\i_post_norm_mul.s_opa_i [26:26]),.s_opa_i_4(\i_post_norm_mul.s_opa_i [27:27]),.s_opa_i_5(\i_post_norm_mul.s_opa_i [28:28]),.s_opa_i_6(\i_post_norm_mul.s_opa_i [29:29]),.s_opa_i_7(\i_post_norm_mul.s_opa_i [30:30]),.s_opa_i_0(s_opa_i[30:23]),.serial_div_rmndr(serial_div_rmndr[26:0]),.serial_div_qutnt(serial_div_qutnt[26:0]),.s_rmode_i(\i_post_norm_mul.s_rmode_i [1:0]),.s_rmode_i_0(s_rmode_i[1:0]),.s_fractb_i(\i_mul_24.s_fractb_i [22:0]),.s_fracta_i(\i_mul_24.s_fracta_i [22:16]),.post_norm_div_output(post_norm_div_output[31:0]),.clk_i(clk_i),.un11_s_exp_10_o_axb_0_i(\i_pre_norm_div.un11_s_exp_10_o_axb_0_i ),.s_infb(\i_post_norm_mul.s_infb ),.un1_s_infa(\i_post_norm_mul.un1_s_infa ),.result_4(\i_post_norm_mul.or_reduce.result_4 ),.N_1942_i(N_1942_i),.post_norm_div_ine(post_norm_div_ine),.result_5(\i_post_norm_mul.or_reduce.result_5 ),.result_3_21_1(\i_post_norm_mul.or_reduce.result_3_21_1 ),.result_3_21_3(\i_post_norm_mul.or_reduce.result_3_21_3 ),.result_11(\i_post_norm_sqrt.or_reduce.result_11 ),.un1_s_nan_a(\i_post_norm_mul.un1_s_nan_a ),.un1_s_nan_b(\i_post_norm_mul.un1_s_nan_b ),.un3_s_op_0(\i_post_norm_mul.un3_s_op_0 ));
  pre_norm_sqrt_inj i_pre_norm_sqrt(.v_count(\i_pre_norm_sqrt.v_count [4:1]),.v_count_i(\i_pre_norm_sqrt.v_count_i ),.v_count_1_0_a2_7_i_0(\i_pre_norm_div.v_count_1_0_a2_7_i_0 ),.v_count_56_0_2(\i_prenorm_addsub.v_count_56_0_2 [4:4]),.pre_norm_sqrt_fracta_o_0(pre_norm_sqrt_fracta_o_0[51:51]),.s_fracta_52_o_0_e(\i_pre_norm_sqrt.s_fracta_52_o_0_e [33:30]),.pre_norm_div_dvdnd_0(pre_norm_div_dvdnd_0[49:49]),.pre_norm_sqrt_exp_o(pre_norm_sqrt_exp_o[7:0]),.v_count_1_0_0_a2_0(\i_pre_norm_div.v_count_1_0_0_a2_0 [1:1]),.v_count_1_0_1(\i_pre_norm_div.v_count_1_0_1 ),.v_count_1_0_2(\i_pre_norm_div.v_count_1_0_2 ),.pre_norm_div_dvdnd_17(pre_norm_div_dvdnd[43:43]),.pre_norm_div_dvdnd_16(pre_norm_div_dvdnd[42:42]),.pre_norm_div_dvdnd_9(pre_norm_div_dvdnd[35:35]),.pre_norm_div_dvdnd_10(pre_norm_div_dvdnd[36:36]),.pre_norm_div_dvdnd_11(pre_norm_div_dvdnd[37:37]),.pre_norm_div_dvdnd_8(pre_norm_div_dvdnd[34:34]),.pre_norm_div_dvdnd_21(pre_norm_div_dvdnd[47:47]),.pre_norm_div_dvdnd_22(pre_norm_div_dvdnd[48:48]),.pre_norm_div_dvdnd_18(pre_norm_div_dvdnd[44:44]),.pre_norm_div_dvdnd_20(pre_norm_div_dvdnd[46:46]),.pre_norm_div_dvdnd_19(pre_norm_div_dvdnd[45:45]),.s_opa_i_23(s_opa_i[23:23]),.s_opa_i_0(s_opa_i[0:0]),.s_opa_i_2(s_opa_i[2:2]),.s_opa_i_3(s_opa_i[3:3]),.s_opa_i_1(s_opa_i[1:1]),.s_opa_i_8(s_opa_i[8:8]),.s_opa_i_10(s_opa_i[10:10]),.s_opa_i_11(s_opa_i[11:11]),.s_opa_i_9(s_opa_i[9:9]),.s_opa_i_6(s_opa_i[6:6]),.s_opa_i_7(s_opa_i[7:7]),.s_opa_i_5(s_opa_i[5:5]),.s_opa_i_4(s_opa_i[4:4]),.s_opa_i_14(s_opa_i[14:14]),.s_opa_i_12(s_opa_i[12:12]),.s_opa_i_13(s_opa_i[13:13]),.s_opa_i_15(s_opa_i[15:15]),.s_opa_i_21(s_opa_i[21:21]),.s_opa_i_22(s_opa_i[22:22]),.s_opa_i_20(s_opa_i[20:20]),.s_opa_i_24(s_opa_i[24:24]),.s_opa_i_30(s_opa_i[30:30]),.s_opa_i_27(s_opa_i[27:27]),.s_opa_i_25(s_opa_i[25:25]),.s_opa_i_26(s_opa_i[26:26]),.pre_norm_sqrt_fracta_o_15(pre_norm_sqrt_fracta_o[43:43]),.pre_norm_sqrt_fracta_o_16(pre_norm_sqrt_fracta_o[44:44]),.pre_norm_sqrt_fracta_o_6(pre_norm_sqrt_fracta_o[34:34]),.pre_norm_sqrt_fracta_o_10(pre_norm_sqrt_fracta_o[38:38]),.pre_norm_sqrt_fracta_o_9(pre_norm_sqrt_fracta_o[37:37]),.pre_norm_sqrt_fracta_o_8(pre_norm_sqrt_fracta_o[36:36]),.pre_norm_sqrt_fracta_o_7(pre_norm_sqrt_fracta_o[35:35]),.pre_norm_sqrt_fracta_o_21(pre_norm_sqrt_fracta_o[49:49]),.pre_norm_sqrt_fracta_o_0_d0(pre_norm_sqrt_fracta_o[28:28]),.pre_norm_sqrt_fracta_o_18(pre_norm_sqrt_fracta_o[46:46]),.pre_norm_sqrt_fracta_o_19(pre_norm_sqrt_fracta_o[47:47]),.pre_norm_sqrt_fracta_o_22(pre_norm_sqrt_fracta_o[50:50]),.pre_norm_sqrt_fracta_o_11(pre_norm_sqrt_fracta_o[39:39]),.pre_norm_sqrt_fracta_o_12(pre_norm_sqrt_fracta_o[40:40]),.pre_norm_sqrt_fracta_o_13(pre_norm_sqrt_fracta_o[41:41]),.pre_norm_sqrt_fracta_o_14(pre_norm_sqrt_fracta_o[42:42]),.pre_norm_sqrt_fracta_o_20(pre_norm_sqrt_fracta_o[48:48]),.s_opa_i_i(s_opa_i_i[29:28]),.N_88(\i_pre_norm_sqrt.s_fracta2_52_o.N_88 ),.N_55(\i_pre_norm_div.s_dvdnd_50_o.N_55 ),.s_dvdnd_50_o_108_0_e(\i_pre_norm_div.s_dvdnd_50_o.s_dvdnd_50_o_108_0_e ),.N_38_0(N_38_0),.N_1620(N_1620),.s_dvdnd_50_o_105_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_105_0_e ),.N_45(\i_pre_norm_sqrt.s_fracta2_52_o.N_45 ),.N_1619(N_1619),.N_41(\i_pre_norm_sqrt.s_fracta2_52_o.N_41 ),.N_1624(N_1624),.N_1087(N_1087),.N_1166(N_1166),.N_1174(N_1174),.un2_s_snan_o_8(un2_s_snan_o_8),.N_95(\i_pre_norm_div.s_dvdnd_50_o.N_95 ),.N_1245(N_1245),.N_53(\i_pre_norm_sqrt.s_fracta2_52_o.N_53 ),.N_48_0(N_48_0),.s_dvdnd_50_o_106_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_106_0_e ),.m49_0_e(\i_prenorm_addsub.m49_0_e ),.s_dvdnd_50_o_102_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_102_0_e ),.s_dvdnd_50_o_109_0_e(\i_pre_norm_sqrt.s_fracta2_52_o.s_dvdnd_50_o_109_0_e ),.N_1238(N_1238),.N_1227(N_1227),.clk_i(clk_i),.un2_s_snan_o_20(un2_s_snan_o_20),.N_1077(N_1077),.N_399(\i_pre_norm_div.N_399 ),.N_396(\i_pre_norm_div.N_396 ),.N_44(\i_pre_norm_sqrt.s_fracta2_52_o.N_44 ),.N_1241(N_1241),.N_30_0(N_30_0),.un2_s_snan_o_22(un2_s_snan_o_22),.result_i_o3_lut6_2_O6(\or_reduce.result_i_o3_lut6_2_O6 ),.N_1242(N_1242),.N_27_0(N_27_0),.N_63(\i_pre_norm_div.s_dvdnd_50_o.N_63 ),.N_1264(N_1264));
  sqrt_inj i_sqrt(.s_state(\i_serial_div.s_state ),.s_fracta_52_o_0_e(\i_pre_norm_sqrt.s_fracta_52_o_0_e [33:29]),.sqrt_sqr_o(sqrt_sqr_o[24:0]),.pre_norm_sqrt_fracta_o_0(pre_norm_sqrt_fracta_o_0[51:51]),.pre_norm_sqrt_fracta_o_14(pre_norm_sqrt_fracta_o[41:41]),.pre_norm_sqrt_fracta_o_15(pre_norm_sqrt_fracta_o[42:42]),.pre_norm_sqrt_fracta_o_16(pre_norm_sqrt_fracta_o[43:43]),.pre_norm_sqrt_fracta_o_17(pre_norm_sqrt_fracta_o[44:44]),.pre_norm_sqrt_fracta_o_18(pre_norm_sqrt_fracta_o[45:45]),.pre_norm_sqrt_fracta_o_19(pre_norm_sqrt_fracta_o[46:46]),.pre_norm_sqrt_fracta_o_20(pre_norm_sqrt_fracta_o[47:47]),.pre_norm_sqrt_fracta_o_21(pre_norm_sqrt_fracta_o[48:48]),.pre_norm_sqrt_fracta_o_22(pre_norm_sqrt_fracta_o[49:49]),.pre_norm_sqrt_fracta_o_23(pre_norm_sqrt_fracta_o[50:50]),.pre_norm_sqrt_fracta_o_0_d0(pre_norm_sqrt_fracta_o[27:27]),.pre_norm_sqrt_fracta_o_1(pre_norm_sqrt_fracta_o[28:28]),.pre_norm_sqrt_fracta_o_7(pre_norm_sqrt_fracta_o[34:34]),.pre_norm_sqrt_fracta_o_8(pre_norm_sqrt_fracta_o[35:35]),.pre_norm_sqrt_fracta_o_9(pre_norm_sqrt_fracta_o[36:36]),.pre_norm_sqrt_fracta_o_10(pre_norm_sqrt_fracta_o[37:37]),.pre_norm_sqrt_fracta_o_11(pre_norm_sqrt_fracta_o[38:38]),.pre_norm_sqrt_fracta_o_12(pre_norm_sqrt_fracta_o[39:39]),.pre_norm_sqrt_fracta_o_13(pre_norm_sqrt_fracta_o[40:40]),.s_start_i(\i_sqrt.s_start_i ),.un12_s_state_0_a2_lut6_2_O5(un12_s_state_0_a2_lut6_2_O5),.clk_i(clk_i),.s_start_i_0(s_start_i),.sqrt_ine_o(sqrt_ine_o));
  post_norm_sqrt_inj i_post_norm_sqrt(.sqrt_sqr_o(sqrt_sqr_o[24:0]),.pre_norm_sqrt_exp_o(pre_norm_sqrt_exp_o[7:0]),.s_rmode_i(\i_post_norm_mul.s_rmode_i [1:0]),.post_norm_sqrt_output(post_norm_sqrt_output[31:0]),.s_signb_i(\i_mul_24.s_signb_i ),.s_signa_i(\i_mul_24.s_signa_i ),.un1_s_infa(\i_post_norm_mul.un1_s_infa ),.result_4(\i_post_norm_mul.or_reduce.result_4 ),.N_6_i(N_6_i),.un1_s_nan_a(\i_post_norm_mul.un1_s_nan_a ),.clk_i(clk_i),.sqrt_ine_o(sqrt_ine_o),.post_norm_sqrt_ine_o(post_norm_sqrt_ine_o));
  LUT2 un1_s_count_4_s_0_RNITDTBG_o6(.I0(s_count_RNIM79LF[21:21]),.I1(un1_s_count_4_s_3),.O(N_80_0_0));
defparam un1_s_count_4_s_0_RNITDTBG_o6.INIT=4'h4;
  LUT2 un1_s_count_4_s_0_RNITDTBG_o5(.I0(s_count_RNIM79LF[21:21]),.I1(un1_s_count_4_s_0),.O(N_2746_0));
defparam un1_s_count_4_s_0_RNITDTBG_o5.INIT=4'h4;
  LUT2 un1_s_count_4_s_2_RNI1ETBG_o6(.I0(s_count_RNIM79LF[21:21]),.I1(un1_s_count_4_s_5),.O(N_2745_0));
defparam un1_s_count_4_s_2_RNI1ETBG_o6.INIT=4'h4;
  LUT2 un1_s_count_4_s_2_RNI1ETBG_o5(.I0(s_count_RNIM79LF[21:21]),.I1(un1_s_count_4_s_2),.O(N_81_0_0));
defparam un1_s_count_4_s_2_RNI1ETBG_o5.INIT=4'h4;
  LUT4 ready_o_e_lut6_2_o6(.I0(ready_o),.I1(s_state),.I2(s_start_i),.I3(s_count_RNIM79LF[21:21]),.O(ready_o_0));
defparam ready_o_e_lut6_2_o6.INIT=16'hAFA8;
  LUT2 ready_o_e_lut6_2_o5(.I0(un1_s_count_4_s_1),.I1(s_count_RNIM79LF[21:21]),.O(N_2715_0));
defparam ready_o_e_lut6_2_o5.INIT=4'h2;
endmodule
