`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[110:0] testVector;
output[201:0] resultVector;
input[413:0] injectionVector;
qr_wrapper_wrapper_inj toplevel_instance (
.clk(clk),
.rst(rst),
.reduced_matrix(testVector[0]),
.start(testVector[1]),
.request_out(testVector[2]),
.valid_out(resultVector[0]),
.ready(resultVector[1]),
.in_A_r(testVector [50:3]),
.in_A_i(testVector [98:51]),
.sigma_in(testVector [110:99]),
.out_Q_r(resultVector [49:2]),
.out_Q_i(resultVector [97:50]),
.out_R_r(resultVector [145:98]),
.out_R_i(resultVector [193:146]),
.permut(resultVector [201:194]),
.p_output_reg_pipe_13_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[0]),
.p_output_reg_pipe_12_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[1]),
.p_output_reg_pipe_Z_p_O_FDshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[2]),
.p_desc951_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[3]),
.p_desc952_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[4]),
.p_desc953_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[5]),
.p_desc954_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[6]),
.p_desc955_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[7]),
.p_desc956_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[8]),
.p_desc957_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[9]),
.p_desc958_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[10]),
.p_desc959_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[11]),
.p_desc960_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[12]),
.p_desc961_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[13]),
.p_desc962_p_O_FDEinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[14]),
.p_desc48_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[15]),
.p_desc49_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[16]),
.p_desc50_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[17]),
.p_desc51_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[18]),
.p_desc52_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[19]),
.p_desc53_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[20]),
.p_desc54_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[21]),
.p_desc55_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[22]),
.p_desc56_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[23]),
.p_desc57_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[24]),
.p_desc58_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[25]),
.p_desc59_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[26]),
.p_desc60_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[27]),
.p_desc61_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[28]),
.p_desc62_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[29]),
.p_desc63_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[30]),
.p_desc64_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[31]),
.p_desc65_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[32]),
.p_desc66_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[33]),
.p_desc67_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[34]),
.p_desc68_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[35]),
.p_desc69_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[36]),
.p_desc70_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[37]),
.p_desc71_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[38]),
.p_desc72_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[39]),
.p_desc73_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[40]),
.p_desc74_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[41]),
.p_desc75_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[42]),
.p_desc76_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[43]),
.p_desc77_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[44]),
.p_desc78_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[45]),
.p_desc79_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[46]),
.p_desc80_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[47]),
.p_desc81_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[48]),
.p_desc82_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[49]),
.p_desc83_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[50]),
.p_desc84_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[51]),
.p_desc85_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[52]),
.p_desc86_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[53]),
.p_desc87_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[54]),
.p_desc88_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[55]),
.p_desc89_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[56]),
.p_desc90_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[57]),
.p_desc91_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[58]),
.p_desc92_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[59]),
.p_desc93_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[60]),
.p_desc94_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[61]),
.p_desc95_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[62]),
.p_desc96_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[63]),
.p_desc97_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[64]),
.p_desc98_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[65]),
.p_desc99_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[66]),
.p_desc100_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[67]),
.p_desc101_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[68]),
.p_desc102_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[69]),
.p_desc103_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[70]),
.p_desc104_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[71]),
.p_desc105_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[72]),
.p_desc106_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[73]),
.p_desc107_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[74]),
.p_desc108_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[75]),
.p_desc109_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[76]),
.p_desc110_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[77]),
.p_desc111_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[78]),
.p_desc112_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[79]),
.p_desc113_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[80]),
.p_desc114_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[81]),
.p_desc115_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[82]),
.p_desc116_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[83]),
.p_desc117_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[84]),
.p_desc118_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[85]),
.p_desc119_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[86]),
.p_desc120_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[87]),
.p_desc121_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[88]),
.p_desc122_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[89]),
.p_desc123_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[90]),
.p_desc124_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[91]),
.p_desc125_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[92]),
.p_desc126_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[93]),
.p_desc127_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[94]),
.p_desc128_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[95]),
.p_desc129_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[96]),
.p_desc130_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[97]),
.p_desc131_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[98]),
.p_desc132_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[99]),
.p_desc133_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[100]),
.p_desc134_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[101]),
.p_desc135_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[102]),
.p_desc136_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[103]),
.p_desc137_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[104]),
.p_desc138_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[105]),
.p_desc139_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[106]),
.p_desc140_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[107]),
.p_desc141_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[108]),
.p_desc142_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[109]),
.p_desc143_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[110]),
.p_desc144_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[111]),
.p_desc145_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[112]),
.p_desc146_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[113]),
.p_desc147_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[114]),
.p_desc148_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[115]),
.p_desc149_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[116]),
.p_desc150_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[117]),
.p_desc151_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[118]),
.p_desc152_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[119]),
.p_desc153_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[120]),
.p_desc154_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[121]),
.p_desc155_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[122]),
.p_desc156_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[123]),
.p_desc157_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[124]),
.p_desc158_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[125]),
.p_desc159_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[126]),
.p_desc160_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[127]),
.p_desc161_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[128]),
.p_desc162_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[129]),
.p_desc163_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[130]),
.p_desc164_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[131]),
.p_desc165_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[132]),
.p_desc166_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[133]),
.p_desc167_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[134]),
.p_desc168_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[135]),
.p_desc169_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[136]),
.p_desc170_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[137]),
.p_desc171_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[138]),
.p_desc172_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[139]),
.p_desc173_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[140]),
.p_desc174_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[141]),
.p_desc175_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[142]),
.p_desc176_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[143]),
.p_desc177_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[144]),
.p_desc178_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[145]),
.p_desc179_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[146]),
.p_desc180_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[147]),
.p_desc181_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[148]),
.p_desc182_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[149]),
.p_desc183_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[150]),
.p_desc184_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[151]),
.p_desc185_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[152]),
.p_desc186_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[153]),
.p_desc187_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[154]),
.p_desc188_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[155]),
.p_desc189_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[156]),
.p_desc190_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[157]),
.p_desc191_p_O_FDEr_mat_regs_qr_decomp_qr_wrapper_(injectionVector[158]),
.p_output_reg_pipe_1_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[159]),
.p_output_reg_pipe_4_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[160]),
.p_output_reg_pipe_5_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[161]),
.p_output_reg_pipe_6_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[162]),
.p_output_reg_pipe_9_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[163]),
.p_output_reg_pipe_10_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[164]),
.p_output_reg_pipe_11_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[165]),
.p_output_reg_pipe_14_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[166]),
.p_output_reg_pipe_15_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[167]),
.p_output_reg_pipe_16_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[168]),
.p_output_reg_pipe_19_Z_p_O_FDEshifterZ0_inv_sqrt_qr_decomp_qr_wrapper_(injectionVector[169]),
.p_desc739_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[170]),
.p_desc740_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[171]),
.p_desc741_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[172]),
.p_desc742_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[173]),
.p_desc743_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[174]),
.p_desc744_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[175]),
.p_desc745_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[176]),
.p_desc746_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[177]),
.p_desc747_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[178]),
.p_desc748_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[179]),
.p_desc749_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[180]),
.p_desc750_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[181]),
.p_desc751_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[182]),
.p_desc752_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[183]),
.p_desc753_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[184]),
.p_desc754_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[185]),
.p_desc755_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[186]),
.p_desc756_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[187]),
.p_desc757_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[188]),
.p_desc758_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[189]),
.p_desc759_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[190]),
.p_desc760_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[191]),
.p_desc761_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[192]),
.p_desc762_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[193]),
.p_desc763_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[194]),
.p_desc764_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[195]),
.p_desc765_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[196]),
.p_desc766_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[197]),
.p_desc767_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[198]),
.p_desc768_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[199]),
.p_desc769_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[200]),
.p_desc770_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[201]),
.p_desc771_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[202]),
.p_desc772_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[203]),
.p_desc773_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[204]),
.p_desc774_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[205]),
.p_desc775_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[206]),
.p_desc776_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[207]),
.p_desc777_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[208]),
.p_desc778_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[209]),
.p_desc779_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[210]),
.p_desc780_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[211]),
.p_desc781_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[212]),
.p_desc782_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[213]),
.p_desc783_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[214]),
.p_desc784_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[215]),
.p_desc785_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[216]),
.p_desc786_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[217]),
.p_desc787_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[218]),
.p_desc788_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[219]),
.p_desc789_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[220]),
.p_desc790_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[221]),
.p_desc791_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[222]),
.p_desc792_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[223]),
.p_desc793_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[224]),
.p_desc794_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[225]),
.p_desc795_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[226]),
.p_desc796_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[227]),
.p_desc797_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[228]),
.p_desc798_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[229]),
.p_desc799_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[230]),
.p_desc800_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[231]),
.p_desc801_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[232]),
.p_desc802_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[233]),
.p_desc803_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[234]),
.p_desc804_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[235]),
.p_desc805_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[236]),
.p_desc806_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[237]),
.p_desc807_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[238]),
.p_desc808_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[239]),
.p_desc809_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[240]),
.p_desc810_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[241]),
.p_desc811_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[242]),
.p_desc812_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[243]),
.p_desc813_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[244]),
.p_desc814_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[245]),
.p_desc815_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[246]),
.p_desc816_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[247]),
.p_desc817_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[248]),
.p_desc818_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[249]),
.p_desc819_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[250]),
.p_desc820_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[251]),
.p_desc821_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[252]),
.p_desc822_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[253]),
.p_desc823_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[254]),
.p_desc824_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[255]),
.p_desc825_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[256]),
.p_desc826_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[257]),
.p_desc827_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[258]),
.p_desc828_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[259]),
.p_desc829_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[260]),
.p_desc830_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[261]),
.p_desc831_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[262]),
.p_desc832_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[263]),
.p_desc833_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[264]),
.p_desc834_p_O_FDEvec_sub_qr_decomp_qr_wrapper_(injectionVector[265]),
.p_output_reg_pipe_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[266]),
.p_output_reg_pipe_3_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[267]),
.p_output_reg_pipe_6_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[268]),
.p_output_reg_pipe_9_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[269]),
.p_output_reg_pipe_12_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[270]),
.p_output_reg_pipe_15_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[271]),
.p_output_reg_pipe_16_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[272]),
.p_output_reg_pipe_17_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[273]),
.p_output_reg_pipe_18_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[274]),
.p_output_reg_pipe_21_Z_p_O_FDREinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[275]),
.p_desc318_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[276]),
.p_desc319_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[277]),
.p_desc320_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[278]),
.p_desc321_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[279]),
.p_desc322_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[280]),
.p_in_reg_enable_fsm_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[281]),
.p_done_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[282]),
.p_acc_enable_Z_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[283]),
.p_desc325_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[284]),
.p_desc326_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[285]),
.p_desc327_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[286]),
.p_desc328_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[287]),
.p_desc329_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[288]),
.p_desc330_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[289]),
.p_desc331_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[290]),
.p_desc332_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[291]),
.p_desc333_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[292]),
.p_desc334_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[293]),
.p_desc335_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[294]),
.p_desc336_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[295]),
.p_desc337_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[296]),
.p_desc338_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[297]),
.p_desc339_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[298]),
.p_desc340_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[299]),
.p_desc341_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[300]),
.p_desc342_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[301]),
.p_desc343_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[302]),
.p_desc344_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[303]),
.p_desc345_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[304]),
.p_desc346_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[305]),
.p_desc347_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[306]),
.p_desc348_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[307]),
.p_desc349_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[308]),
.p_desc350_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[309]),
.p_desc375_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[310]),
.p_desc376_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[311]),
.p_desc377_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[312]),
.p_desc378_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[313]),
.p_desc379_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[314]),
.p_desc380_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[315]),
.p_desc381_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[316]),
.p_desc382_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[317]),
.p_desc383_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[318]),
.p_desc384_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[319]),
.p_desc385_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[320]),
.p_desc386_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[321]),
.p_desc387_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[322]),
.p_desc388_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[323]),
.p_desc389_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[324]),
.p_desc390_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[325]),
.p_desc391_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[326]),
.p_desc392_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[327]),
.p_desc393_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[328]),
.p_desc394_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[329]),
.p_desc395_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[330]),
.p_desc396_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[331]),
.p_desc397_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[332]),
.p_desc398_p_O_FDCinner_prod_qr_decomp_qr_wrapper_(injectionVector[333]),
.p_done_Z_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[334]),
.p_desc946_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[335]),
.p_desc947_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[336]),
.p_desc948_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[337]),
.p_desc949_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[338]),
.p_desc950_p_O_FDCinv_sqrt_qr_decomp_qr_wrapper_(injectionVector[339]),
.p_desc1255_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[340]),
.p_desc1256_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[341]),
.p_desc1257_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[342]),
.p_desc1258_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[343]),
.p_start_inner_prod_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[344]),
.p_wr_en_AQ_int_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[345]),
.p_wr_en_R_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[346]),
.p_w_in_a_vec_sub_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[347]),
.p_start_inv_sqrt_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[348]),
.p_desc1274_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[349]),
.p_pre_red_mat_reg_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[350]),
.p_done_Z_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[351]),
.p_desc1275_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[352]),
.p_desc1276_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[353]),
.p_desc1277_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[354]),
.p_desc1278_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[355]),
.p_desc1279_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[356]),
.p_desc1281_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[357]),
.p_desc1282_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[358]),
.p_desc1283_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[359]),
.p_desc1284_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[360]),
.p_desc1285_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[361]),
.p_desc1286_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[362]),
.p_desc1287_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[363]),
.p_desc1288_p_O_FDCqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[364]),
.p_start_QR_Z_p_O_FDCqr_wrapper_(injectionVector[365]),
.p_wr_A_QR_Z_p_O_FDCqr_wrapper_(injectionVector[366]),
.p_valid_out_Z_p_O_FDCqr_wrapper_(injectionVector[367]),
.p_ready_Z_p_O_FDCqr_wrapper_(injectionVector[368]),
.p_red_mat_reg_Z_p_O_FDCqr_wrapper_(injectionVector[369]),
.p_desc1317_p_O_FDCqr_wrapper_(injectionVector[370]),
.p_desc1318_p_O_FDCqr_wrapper_(injectionVector[371]),
.p_desc1319_p_O_FDCqr_wrapper_(injectionVector[372]),
.p_desc1320_p_O_FDCqr_wrapper_(injectionVector[373]),
.p_desc1321_p_O_FDCqr_wrapper_(injectionVector[374]),
.p_desc1322_p_O_FDCqr_wrapper_(injectionVector[375]),
.p_acc_clear_Z_p_O_FDPinner_prod_qr_decomp_qr_wrapper_(injectionVector[376]),
.p_desc1265_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[377]),
.p_desc1268_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[378]),
.p_desc1280_p_O_FDPqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[379]),
.p_desc324_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[380]),
.p_desc351_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[381]),
.p_desc352_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[382]),
.p_desc353_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[383]),
.p_desc354_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[384]),
.p_desc355_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[385]),
.p_desc356_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[386]),
.p_desc357_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[387]),
.p_desc358_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[388]),
.p_desc359_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[389]),
.p_desc360_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[390]),
.p_desc361_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[391]),
.p_desc362_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[392]),
.p_desc363_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[393]),
.p_desc364_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[394]),
.p_desc365_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[395]),
.p_desc366_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[396]),
.p_desc367_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[397]),
.p_desc368_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[398]),
.p_desc369_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[399]),
.p_desc370_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[400]),
.p_desc371_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[401]),
.p_desc372_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[402]),
.p_desc373_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[403]),
.p_desc374_p_O_FDCEinner_prod_qr_decomp_qr_wrapper_(injectionVector[404]),
.p_desc1263_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[405]),
.p_desc1264_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[406]),
.p_desc1266_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[407]),
.p_desc1267_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[408]),
.p_desc1269_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[409]),
.p_desc1270_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[410]),
.p_desc1271_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[411]),
.p_desc1272_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[412]),
.p_desc1273_p_O_FDCEqr_decomp_ctl_qr_decomp_qr_wrapper_(injectionVector[413]));
endmodule