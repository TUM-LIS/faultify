`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[68:0] testVector;
output[4:0] resultVector;
input[281:0] injectionVector;
dec_viterbi_inj toplevel_instance (
.aclk(clk),
.aresetn(rst),
.s_axis_input_tvalid(testVector[0]),
.s_axis_input_tdata(testVector [32:1]),
.s_axis_input_tlast(testVector[33]),
.s_axis_input_tready(resultVector[0]),
.m_axis_output_tvalid(resultVector[1]),
.m_axis_output_tdata(resultVector[2]),
.m_axis_output_tlast(resultVector[3]),
.m_axis_output_tready(testVector[34]),
.s_axis_ctrl_tvalid(testVector[35]),
.s_axis_ctrl_tdata(testVector [67:36]),
.s_axis_ctrl_tlast(testVector[68]),
.s_axis_ctrl_tready(resultVector[4]),
.p_desc95_p_O_FDacsZ0_(injectionVector[0]),
.p_desc96_p_O_FDacsZ0_(injectionVector[1]),
.p_desc134_p_O_FDacsZ0_1_(injectionVector[2]),
.p_desc135_p_O_FDacsZ0_1_(injectionVector[3]),
.p_desc173_p_O_FDacsZ0_2_(injectionVector[4]),
.p_desc174_p_O_FDacsZ0_2_(injectionVector[5]),
.p_desc212_p_O_FDacsZ0_3_(injectionVector[6]),
.p_desc213_p_O_FDacsZ0_3_(injectionVector[7]),
.p_desc251_p_O_FDacsZ0_4_(injectionVector[8]),
.p_desc252_p_O_FDacsZ0_4_(injectionVector[9]),
.p_desc290_p_O_FDacsZ0_5_(injectionVector[10]),
.p_desc291_p_O_FDacsZ0_5_(injectionVector[11]),
.p_desc329_p_O_FDacsZ0_6_(injectionVector[12]),
.p_desc330_p_O_FDacsZ0_6_(injectionVector[13]),
.p_desc368_p_O_FDacsZ0_7_(injectionVector[14]),
.p_desc369_p_O_FDacsZ0_7_(injectionVector[15]),
.p_desc407_p_O_FDacsZ0_8_(injectionVector[16]),
.p_desc408_p_O_FDacsZ0_8_(injectionVector[17]),
.p_desc446_p_O_FDacsZ0_9_(injectionVector[18]),
.p_desc447_p_O_FDacsZ0_9_(injectionVector[19]),
.p_desc485_p_O_FDacsZ0_10_(injectionVector[20]),
.p_desc486_p_O_FDacsZ0_10_(injectionVector[21]),
.p_desc524_p_O_FDacsZ0_11_(injectionVector[22]),
.p_desc525_p_O_FDacsZ0_11_(injectionVector[23]),
.p_desc563_p_O_FDacsZ0_12_(injectionVector[24]),
.p_desc564_p_O_FDacsZ0_12_(injectionVector[25]),
.p_desc602_p_O_FDacsZ0_13_(injectionVector[26]),
.p_desc603_p_O_FDacsZ0_13_(injectionVector[27]),
.p_desc641_p_O_FDacsZ0_14_(injectionVector[28]),
.p_desc642_p_O_FDacsZ0_14_(injectionVector[29]),
.p_desc680_p_O_FDacsZ0_15_(injectionVector[30]),
.p_desc681_p_O_FDacsZ0_15_(injectionVector[31]),
.p_desc719_p_O_FDacsZ0_16_(injectionVector[32]),
.p_desc720_p_O_FDacsZ0_16_(injectionVector[33]),
.p_desc758_p_O_FDacsZ0_17_(injectionVector[34]),
.p_desc759_p_O_FDacsZ0_17_(injectionVector[35]),
.p_desc797_p_O_FDacsZ0_18_(injectionVector[36]),
.p_desc798_p_O_FDacsZ0_18_(injectionVector[37]),
.p_desc873_p_O_FDacsZ0_20_(injectionVector[38]),
.p_desc874_p_O_FDacsZ0_20_(injectionVector[39]),
.p_desc912_p_O_FDacsZ0_21_(injectionVector[40]),
.p_desc913_p_O_FDacsZ0_21_(injectionVector[41]),
.p_desc989_p_O_FDacsZ0_22_(injectionVector[42]),
.p_desc990_p_O_FDacsZ0_22_(injectionVector[43]),
.p_desc1028_p_O_FDacsZ0_23_(injectionVector[44]),
.p_desc1029_p_O_FDacsZ0_23_(injectionVector[45]),
.p_desc1067_p_O_FDacsZ0_24_(injectionVector[46]),
.p_desc1068_p_O_FDacsZ0_24_(injectionVector[47]),
.p_desc1106_p_O_FDacsZ0_25_(injectionVector[48]),
.p_desc1107_p_O_FDacsZ0_25_(injectionVector[49]),
.p_desc1145_p_O_FDacsZ0_26_(injectionVector[50]),
.p_desc1146_p_O_FDacsZ0_26_(injectionVector[51]),
.p_desc1184_p_O_FDacsZ0_27_(injectionVector[52]),
.p_desc1185_p_O_FDacsZ0_27_(injectionVector[53]),
.p_desc1223_p_O_FDacsZ0_28_(injectionVector[54]),
.p_desc1224_p_O_FDacsZ0_28_(injectionVector[55]),
.p_desc1262_p_O_FDacsZ0_29_(injectionVector[56]),
.p_desc1263_p_O_FDacsZ0_29_(injectionVector[57]),
.p_desc1301_p_O_FDacsZ0_30_(injectionVector[58]),
.p_desc1302_p_O_FDacsZ0_30_(injectionVector[59]),
.p_desc1340_p_O_FDacsZ0_31_(injectionVector[60]),
.p_desc1341_p_O_FDacsZ0_31_(injectionVector[61]),
.p_desc1379_p_O_FDacsZ0_32_(injectionVector[62]),
.p_desc1380_p_O_FDacsZ0_32_(injectionVector[63]),
.p_desc1418_p_O_FDacsZ0_33_(injectionVector[64]),
.p_desc1419_p_O_FDacsZ0_33_(injectionVector[65]),
.p_desc1457_p_O_FDacsZ0_34_(injectionVector[66]),
.p_desc1458_p_O_FDacsZ0_34_(injectionVector[67]),
.p_desc1496_p_O_FDacsZ0_35_(injectionVector[68]),
.p_desc1497_p_O_FDacsZ0_35_(injectionVector[69]),
.p_desc1535_p_O_FDacsZ0_36_(injectionVector[70]),
.p_desc1536_p_O_FDacsZ0_36_(injectionVector[71]),
.p_desc1574_p_O_FDacsZ0_37_(injectionVector[72]),
.p_desc1575_p_O_FDacsZ0_37_(injectionVector[73]),
.p_desc1613_p_O_FDacsZ0_38_(injectionVector[74]),
.p_desc1614_p_O_FDacsZ0_38_(injectionVector[75]),
.p_desc1652_p_O_FDacsZ0_39_(injectionVector[76]),
.p_desc1653_p_O_FDacsZ0_39_(injectionVector[77]),
.p_desc1691_p_O_FDacsZ0_40_(injectionVector[78]),
.p_desc1692_p_O_FDacsZ0_40_(injectionVector[79]),
.p_desc1730_p_O_FDacsZ0_41_(injectionVector[80]),
.p_desc1731_p_O_FDacsZ0_41_(injectionVector[81]),
.p_desc1769_p_O_FDacsZ0_42_(injectionVector[82]),
.p_desc1770_p_O_FDacsZ0_42_(injectionVector[83]),
.p_desc1808_p_O_FDacsZ0_43_(injectionVector[84]),
.p_desc1809_p_O_FDacsZ0_43_(injectionVector[85]),
.p_desc1847_p_O_FDacsZ0_44_(injectionVector[86]),
.p_desc1848_p_O_FDacsZ0_44_(injectionVector[87]),
.p_desc1886_p_O_FDacsZ0_45_(injectionVector[88]),
.p_desc1887_p_O_FDacsZ0_45_(injectionVector[89]),
.p_desc1925_p_O_FDacsZ0_46_(injectionVector[90]),
.p_desc1926_p_O_FDacsZ0_46_(injectionVector[91]),
.p_desc1964_p_O_FDacsZ0_47_(injectionVector[92]),
.p_desc1965_p_O_FDacsZ0_47_(injectionVector[93]),
.p_desc2003_p_O_FDacsZ0_48_(injectionVector[94]),
.p_desc2004_p_O_FDacsZ0_48_(injectionVector[95]),
.p_desc2042_p_O_FDacsZ0_49_(injectionVector[96]),
.p_desc2043_p_O_FDacsZ0_49_(injectionVector[97]),
.p_desc2081_p_O_FDacsZ0_50_(injectionVector[98]),
.p_desc2082_p_O_FDacsZ0_50_(injectionVector[99]),
.p_desc2120_p_O_FDacsZ0_51_(injectionVector[100]),
.p_desc2121_p_O_FDacsZ0_51_(injectionVector[101]),
.p_desc2159_p_O_FDacsZ0_52_(injectionVector[102]),
.p_desc2160_p_O_FDacsZ0_52_(injectionVector[103]),
.p_desc2198_p_O_FDacsZ0_53_(injectionVector[104]),
.p_desc2199_p_O_FDacsZ0_53_(injectionVector[105]),
.p_desc2237_p_O_FDacsZ0_54_(injectionVector[106]),
.p_desc2238_p_O_FDacsZ0_54_(injectionVector[107]),
.p_desc2276_p_O_FDacsZ0_55_(injectionVector[108]),
.p_desc2277_p_O_FDacsZ0_55_(injectionVector[109]),
.p_desc2315_p_O_FDacsZ0_56_(injectionVector[110]),
.p_desc2316_p_O_FDacsZ0_56_(injectionVector[111]),
.p_desc2354_p_O_FDacsZ0_57_(injectionVector[112]),
.p_desc2355_p_O_FDacsZ0_57_(injectionVector[113]),
.p_desc2393_p_O_FDacsZ0_58_(injectionVector[114]),
.p_desc2394_p_O_FDacsZ0_58_(injectionVector[115]),
.p_desc2432_p_O_FDacsZ0_59_(injectionVector[116]),
.p_desc2433_p_O_FDacsZ0_59_(injectionVector[117]),
.p_desc2471_p_O_FDacsZ0_60_(injectionVector[118]),
.p_desc2472_p_O_FDacsZ0_60_(injectionVector[119]),
.p_desc2510_p_O_FDacsZ0_61_(injectionVector[120]),
.p_desc2511_p_O_FDacsZ0_61_(injectionVector[121]),
.p_desc2549_p_O_FDacsZ0_62_(injectionVector[122]),
.p_desc2550_p_O_FDacsZ0_62_(injectionVector[123]),
.p_m_axis_output_tdata_0_rep2_Z_p_O_FDREbranch_distanceZ3_(injectionVector[124]),
.p_m_axis_output_tdata_0_rep1_Z_p_O_FDREbranch_distanceZ3_(injectionVector[125]),
.p_desc31_p_O_FDREbranch_distanceZ3_(injectionVector[126]),
.p_desc32_p_O_FDREbranch_distanceZ3_(injectionVector[127]),
.p_desc33_p_O_FDREbranch_distanceZ3_(injectionVector[128]),
.p_desc34_p_O_FDREbranch_distanceZ3_(injectionVector[129]),
.p_desc35_p_O_FDREbranch_distanceZ3_(injectionVector[130]),
.p_desc36_p_O_FDREbranch_distanceZ3_(injectionVector[131]),
.p_desc37_p_O_FDREbranch_distanceZ3_(injectionVector[132]),
.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ2_(injectionVector[133]),
.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ2_(injectionVector[134]),
.p_desc39_p_O_FDREbranch_distanceZ2_(injectionVector[135]),
.p_desc52_p_O_FDREbranch_distanceZ2_(injectionVector[136]),
.p_desc53_p_O_FDREbranch_distanceZ2_(injectionVector[137]),
.p_desc54_p_O_FDREbranch_distanceZ2_(injectionVector[138]),
.p_desc55_p_O_FDREbranch_distanceZ2_(injectionVector[139]),
.p_desc56_p_O_FDREbranch_distanceZ2_(injectionVector[140]),
.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ0_(injectionVector[141]),
.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ0_(injectionVector[142]),
.p_desc63_p_O_FDREbranch_distanceZ0_(injectionVector[143]),
.p_desc78_p_O_FDREbranch_distanceZ0_(injectionVector[144]),
.p_desc79_p_O_FDREbranch_distanceZ0_(injectionVector[145]),
.p_desc80_p_O_FDREbranch_distanceZ0_(injectionVector[146]),
.p_desc81_p_O_FDREbranch_distanceZ0_(injectionVector[147]),
.p_desc82_p_O_FDREbranch_distanceZ0_(injectionVector[148]),
.p_m_axis_output_tdata_1_0_rep2_Z_p_O_FDREbranch_distanceZ1_(injectionVector[149]),
.p_m_axis_output_tdata_1_0_rep1_Z_p_O_FDREbranch_distanceZ1_(injectionVector[150]),
.p_desc83_p_O_FDREbranch_distanceZ1_(injectionVector[151]),
.p_desc84_p_O_FDREbranch_distanceZ1_(injectionVector[152]),
.p_desc85_p_O_FDREbranch_distanceZ1_(injectionVector[153]),
.p_desc86_p_O_FDREbranch_distanceZ1_(injectionVector[154]),
.p_desc87_p_O_FDREbranch_distanceZ1_(injectionVector[155]),
.p_desc88_p_O_FDREbranch_distanceZ1_(injectionVector[156]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_(injectionVector[157]),
.p_desc125_p_O_FDREacsZ0_(injectionVector[158]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_1_(injectionVector[159]),
.p_desc164_p_O_FDREacsZ0_1_(injectionVector[160]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_2_(injectionVector[161]),
.p_desc203_p_O_FDREacsZ0_2_(injectionVector[162]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_3_(injectionVector[163]),
.p_desc242_p_O_FDREacsZ0_3_(injectionVector[164]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_4_(injectionVector[165]),
.p_desc281_p_O_FDREacsZ0_4_(injectionVector[166]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_5_(injectionVector[167]),
.p_desc320_p_O_FDREacsZ0_5_(injectionVector[168]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_6_(injectionVector[169]),
.p_desc359_p_O_FDREacsZ0_6_(injectionVector[170]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_7_(injectionVector[171]),
.p_desc398_p_O_FDREacsZ0_7_(injectionVector[172]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_8_(injectionVector[173]),
.p_desc437_p_O_FDREacsZ0_8_(injectionVector[174]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_9_(injectionVector[175]),
.p_desc476_p_O_FDREacsZ0_9_(injectionVector[176]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_10_(injectionVector[177]),
.p_desc515_p_O_FDREacsZ0_10_(injectionVector[178]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_11_(injectionVector[179]),
.p_desc554_p_O_FDREacsZ0_11_(injectionVector[180]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_12_(injectionVector[181]),
.p_desc593_p_O_FDREacsZ0_12_(injectionVector[182]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_13_(injectionVector[183]),
.p_desc632_p_O_FDREacsZ0_13_(injectionVector[184]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_14_(injectionVector[185]),
.p_desc671_p_O_FDREacsZ0_14_(injectionVector[186]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_15_(injectionVector[187]),
.p_desc710_p_O_FDREacsZ0_15_(injectionVector[188]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_16_(injectionVector[189]),
.p_desc749_p_O_FDREacsZ0_16_(injectionVector[190]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_17_(injectionVector[191]),
.p_desc788_p_O_FDREacsZ0_17_(injectionVector[192]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_18_(injectionVector[193]),
.p_desc827_p_O_FDREacsZ0_18_(injectionVector[194]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_19_(injectionVector[195]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_20_(injectionVector[196]),
.p_desc903_p_O_FDREacsZ0_20_(injectionVector[197]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_21_(injectionVector[198]),
.p_desc942_p_O_FDREacsZ0_21_(injectionVector[199]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_22_(injectionVector[200]),
.p_desc1019_p_O_FDREacsZ0_22_(injectionVector[201]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_23_(injectionVector[202]),
.p_desc1058_p_O_FDREacsZ0_23_(injectionVector[203]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_24_(injectionVector[204]),
.p_desc1097_p_O_FDREacsZ0_24_(injectionVector[205]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_25_(injectionVector[206]),
.p_desc1136_p_O_FDREacsZ0_25_(injectionVector[207]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_26_(injectionVector[208]),
.p_desc1175_p_O_FDREacsZ0_26_(injectionVector[209]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_27_(injectionVector[210]),
.p_desc1214_p_O_FDREacsZ0_27_(injectionVector[211]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_28_(injectionVector[212]),
.p_desc1253_p_O_FDREacsZ0_28_(injectionVector[213]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_29_(injectionVector[214]),
.p_desc1292_p_O_FDREacsZ0_29_(injectionVector[215]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_30_(injectionVector[216]),
.p_desc1331_p_O_FDREacsZ0_30_(injectionVector[217]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_31_(injectionVector[218]),
.p_desc1370_p_O_FDREacsZ0_31_(injectionVector[219]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_32_(injectionVector[220]),
.p_desc1409_p_O_FDREacsZ0_32_(injectionVector[221]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_33_(injectionVector[222]),
.p_desc1448_p_O_FDREacsZ0_33_(injectionVector[223]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_34_(injectionVector[224]),
.p_desc1487_p_O_FDREacsZ0_34_(injectionVector[225]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_35_(injectionVector[226]),
.p_desc1526_p_O_FDREacsZ0_35_(injectionVector[227]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_36_(injectionVector[228]),
.p_desc1565_p_O_FDREacsZ0_36_(injectionVector[229]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_37_(injectionVector[230]),
.p_desc1604_p_O_FDREacsZ0_37_(injectionVector[231]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_38_(injectionVector[232]),
.p_desc1643_p_O_FDREacsZ0_38_(injectionVector[233]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_39_(injectionVector[234]),
.p_desc1682_p_O_FDREacsZ0_39_(injectionVector[235]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_40_(injectionVector[236]),
.p_desc1721_p_O_FDREacsZ0_40_(injectionVector[237]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_41_(injectionVector[238]),
.p_desc1760_p_O_FDREacsZ0_41_(injectionVector[239]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_42_(injectionVector[240]),
.p_desc1799_p_O_FDREacsZ0_42_(injectionVector[241]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_43_(injectionVector[242]),
.p_desc1838_p_O_FDREacsZ0_43_(injectionVector[243]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_44_(injectionVector[244]),
.p_desc1877_p_O_FDREacsZ0_44_(injectionVector[245]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_45_(injectionVector[246]),
.p_desc1916_p_O_FDREacsZ0_45_(injectionVector[247]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_46_(injectionVector[248]),
.p_desc1955_p_O_FDREacsZ0_46_(injectionVector[249]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_47_(injectionVector[250]),
.p_desc1994_p_O_FDREacsZ0_47_(injectionVector[251]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_48_(injectionVector[252]),
.p_desc2033_p_O_FDREacsZ0_48_(injectionVector[253]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_49_(injectionVector[254]),
.p_desc2072_p_O_FDREacsZ0_49_(injectionVector[255]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_50_(injectionVector[256]),
.p_desc2111_p_O_FDREacsZ0_50_(injectionVector[257]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_51_(injectionVector[258]),
.p_desc2150_p_O_FDREacsZ0_51_(injectionVector[259]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_52_(injectionVector[260]),
.p_desc2189_p_O_FDREacsZ0_52_(injectionVector[261]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_53_(injectionVector[262]),
.p_desc2228_p_O_FDREacsZ0_53_(injectionVector[263]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_54_(injectionVector[264]),
.p_desc2267_p_O_FDREacsZ0_54_(injectionVector[265]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_55_(injectionVector[266]),
.p_desc2306_p_O_FDREacsZ0_55_(injectionVector[267]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_56_(injectionVector[268]),
.p_desc2345_p_O_FDREacsZ0_56_(injectionVector[269]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_57_(injectionVector[270]),
.p_desc2384_p_O_FDREacsZ0_57_(injectionVector[271]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_58_(injectionVector[272]),
.p_desc2423_p_O_FDREacsZ0_58_(injectionVector[273]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_59_(injectionVector[274]),
.p_desc2462_p_O_FDREacsZ0_59_(injectionVector[275]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_60_(injectionVector[276]),
.p_desc2501_p_O_FDREacsZ0_60_(injectionVector[277]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_61_(injectionVector[278]),
.p_desc2540_p_O_FDREacsZ0_61_(injectionVector[279]),
.p_m_axis_outdec_tdata_Z_p_O_FDREacsZ0_62_(injectionVector[280]),
.p_desc2579_p_O_FDREacsZ0_62_(injectionVector[281]));
endmodule