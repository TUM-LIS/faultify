

(* blackbox *)
module DFFX1 (input CLK, D, output Q, QN, input VDD, VSS);
endmodule

(* blackbox *)
module DFFX2 (input CLK, D, output Q, QN, input VDD, VSS);
endmodule


(* blackbox *)
module DFFARX1 (input CLK, D, output Q, QN, input RSTB, VDD, VSS);
endmodule

(* blackbox *)
module DFFSSRX1 (input CLK, D, output Q, QN, input RSTB, SETB, VDD, VSS);
endmodule

(* blackbox *)
module INVX0 (input INP, input VDD, input VSS, output ZN);
endmodule

(* blackbox *)
module AO21X1 (input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AO22X1 (input IN1, IN2, IN3, IN4, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AO22X2 (input IN1, IN2, IN3, IN4, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module OR2X1 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module OR4X1 ( input IN1, IN2, IN3, IN4, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XOR2X1 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XOR2X2 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XOR3X1 ( input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XOR3X2 ( input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module NAND2X0 (input IN1, IN2, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NOR2X0 (input IN1, IN2, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OR3X1 (input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module NOR3X0 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NOR3X1 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NOR4X0 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NOR4X1 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NAND2X1 (input IN1, IN2, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NAND3X0 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NAND3X1 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NAND3X4 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module NAND4X0 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module AND2X1 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AND2X2 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AND2X4 ( input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AND3X1 ( input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AND4X1 ( input IN1, IN2, IN3, IN4, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XNOR2X1 (input IN1, IN2, output Q, input VDD, VSS);
endmodule


(* blackbox *)
module XNOR2X2 (input IN1, IN2, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module XNOR3X1 (input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module OAI22X1 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OAI22X2 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OA22X1 (input IN1, IN2, IN3, IN4, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AOI22X1 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule


(* blackbox *)
module AOI22X2 (input IN1, IN2, IN3, IN4, output QN, input VDD, VSS);
endmodule


(* blackbox *)
module OAI21X1 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OAI21X2 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OA221X1 (input IN1, IN2, IN3, IN4, IN5, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AOI21X1 (input IN1, IN2, IN3, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module AO221X1 (input IN1, input IN2, input IN3, input IN4, input IN5, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AO221X2 (input IN1, input IN2, input IN3, input IN4, input IN5, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AO222X1 (input IN1, IN2, IN3, IN4, IN5, IN6, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module AOI221X1 (input IN1, IN2, IN3, IN4, IN5, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module AOI221X2 (input IN1, IN2, IN3, IN4, IN5, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module AOI222X1 (input IN1, IN2, IN3, IN4, IN5, IN6, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module AOI222X2 (input IN1, IN2, IN3, IN4, IN5, IN6, output QN, input VDD, VSS);
endmodule


(* blackbox *)
module OA222X1 (input IN1, IN2, IN3, IN4, IN5, IN6, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module OA222X2 (input IN1, IN2, IN3, IN4, IN5, IN6, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module OAI221X1 (input IN1, IN2, IN3, IN4, IN5, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OAI222X1 (input IN1, IN2, IN3, IN4, IN5, IN6, output QN, input VDD, VSS);
endmodule

(* blackbox *)
module OA21X1 (input IN1, IN2, IN3, output Q, input VDD, VSS);
endmodule

(* blackbox *)
module FADDX1 (input A, B, CI, output CO, S, input VDD, VSS);
endmodule

(* blackbox *)
module FADDX2 (input A, B, CI, output CO, S, input VDD, VSS);
endmodule

(* blackbox *)
module HADDX1 (input A0, B0, output C1, S0, input VDD, VSS);
endmodule

(* blackbox *)
module HADDX2 (input A0, B0, output C1, S0, input VDD, VSS);
endmodule

(* blackbox *)
module NBUFFX2 (input INP, VDD, VSS, output Z);
endmodule

(* blackbox *)
module NBUFFX4 (input INP, VDD, VSS, output Z);
endmodule

(* blackbox *)
module NBUFFX8 (input INP, VDD, VSS, output Z);
endmodule

(* blackbox *)
module NBUFFX16 (input INP, VDD, VSS, output Z);
endmodule

(* blackbox *)
module MUX21X1 (input IN1, IN2, output Q, input S, VDD, VSS);
endmodule

(* blackbox *)
module MUX21X2 (input IN1, IN2, output Q, input S, VDD, VSS);
endmodule

(* blackbox *)
module MUX41X1 (input IN1, IN2, IN3, IN4, output Q, input S0, S1, VDD, VSS);
endmodule

(* blackbox *)
module MUX41X2 (input IN1, IN2, IN3, IN4, output Q, input S0, S1, VDD, VSS);
endmodule


(* blackbox *)
module DELLN1X2 (input INP, VDD, VSS, output Z);
endmodule

(* blackbox *)
module DELLN2X2 (input INP, VDD, VSS, output Z);
endmodule


