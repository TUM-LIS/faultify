`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[267:0] injectionVector;
fpu_inj toplevel_instance (
.clk_i(clk),
.opa_i(testVector [31:0]),
.opb_i(testVector [63:32]),
.fpu_op_i(testVector [66:64]),
.rmode_i(testVector [68:67]),
.output_o(resultVector [31:0]),
.start_i(testVector[69]),
.ready_o(resultVector[32]),
.ine_o(resultVector[33]),
.overflow_o(resultVector[34]),
.underflow_o(resultVector[35]),
.div_zero_o(resultVector[36]),
.inf_o(resultVector[37]),
.zero_o(resultVector[38]),
.qnan_o(resultVector[39]),
.snan_o(resultVector[40]),
.p_desc1797_p_O_FDpre_norm_div_(injectionVector[0]),
.p_desc1806_p_O_FDpre_norm_div_(injectionVector[1]),
.p_desc1930_p_O_FDserial_div_(injectionVector[2]),
.p_desc1931_p_O_FDserial_div_(injectionVector[3]),
.p_desc1932_p_O_FDserial_div_(injectionVector[4]),
.p_desc1933_p_O_FDserial_div_(injectionVector[5]),
.p_desc1934_p_O_FDserial_div_(injectionVector[6]),
.p_desc1935_p_O_FDserial_div_(injectionVector[7]),
.p_desc1936_p_O_FDserial_div_(injectionVector[8]),
.p_desc1937_p_O_FDserial_div_(injectionVector[9]),
.p_desc1938_p_O_FDserial_div_(injectionVector[10]),
.p_desc1939_p_O_FDserial_div_(injectionVector[11]),
.p_desc1940_p_O_FDserial_div_(injectionVector[12]),
.p_desc1941_p_O_FDserial_div_(injectionVector[13]),
.p_desc1942_p_O_FDserial_div_(injectionVector[14]),
.p_desc1943_p_O_FDserial_div_(injectionVector[15]),
.p_desc1984_p_O_FDserial_div_(injectionVector[16]),
.p_desc1985_p_O_FDserial_div_(injectionVector[17]),
.p_desc1986_p_O_FDserial_div_(injectionVector[18]),
.p_desc1987_p_O_FDserial_div_(injectionVector[19]),
.p_desc1988_p_O_FDserial_div_(injectionVector[20]),
.p_desc1989_p_O_FDserial_div_(injectionVector[21]),
.p_desc1990_p_O_FDserial_div_(injectionVector[22]),
.p_desc1991_p_O_FDserial_div_(injectionVector[23]),
.p_desc1992_p_O_FDserial_div_(injectionVector[24]),
.p_desc1993_p_O_FDserial_div_(injectionVector[25]),
.p_desc1994_p_O_FDserial_div_(injectionVector[26]),
.p_desc1995_p_O_FDserial_div_(injectionVector[27]),
.p_desc1996_p_O_FDserial_div_(injectionVector[28]),
.p_desc1997_p_O_FDserial_div_(injectionVector[29]),
.p_desc1998_p_O_FDserial_div_(injectionVector[30]),
.p_desc1999_p_O_FDserial_div_(injectionVector[31]),
.p_desc2000_p_O_FDserial_div_(injectionVector[32]),
.p_desc2001_p_O_FDserial_div_(injectionVector[33]),
.p_desc2002_p_O_FDserial_div_(injectionVector[34]),
.p_desc2003_p_O_FDserial_div_(injectionVector[35]),
.p_desc2004_p_O_FDserial_div_(injectionVector[36]),
.p_desc2005_p_O_FDserial_div_(injectionVector[37]),
.p_desc2006_p_O_FDserial_div_(injectionVector[38]),
.p_desc2007_p_O_FDserial_div_(injectionVector[39]),
.p_desc2008_p_O_FDserial_div_(injectionVector[40]),
.p_desc2009_p_O_FDserial_div_(injectionVector[41]),
.p_desc2010_p_O_FDserial_div_(injectionVector[42]),
.p_desc2011_p_O_FDserial_div_(injectionVector[43]),
.p_desc2012_p_O_FDserial_div_(injectionVector[44]),
.p_desc2013_p_O_FDserial_div_(injectionVector[45]),
.p_desc2014_p_O_FDserial_div_(injectionVector[46]),
.p_desc2015_p_O_FDserial_div_(injectionVector[47]),
.p_desc2016_p_O_FDserial_div_(injectionVector[48]),
.p_desc2017_p_O_FDserial_div_(injectionVector[49]),
.p_desc2261_p_O_FDpost_norm_div_(injectionVector[50]),
.p_desc2262_p_O_FDpost_norm_div_(injectionVector[51]),
.p_desc2263_p_O_FDpost_norm_div_(injectionVector[52]),
.p_desc2264_p_O_FDpost_norm_div_(injectionVector[53]),
.p_desc2265_p_O_FDpost_norm_div_(injectionVector[54]),
.p_desc2266_p_O_FDpost_norm_div_(injectionVector[55]),
.p_desc2267_p_O_FDpost_norm_div_(injectionVector[56]),
.p_desc2268_p_O_FDpost_norm_div_(injectionVector[57]),
.p_desc2269_p_O_FDpost_norm_div_(injectionVector[58]),
.p_desc2270_p_O_FDpost_norm_div_(injectionVector[59]),
.p_desc2271_p_O_FDpost_norm_div_(injectionVector[60]),
.p_desc2272_p_O_FDpost_norm_div_(injectionVector[61]),
.p_desc2273_p_O_FDpost_norm_div_(injectionVector[62]),
.p_desc2274_p_O_FDpost_norm_div_(injectionVector[63]),
.p_desc2275_p_O_FDpost_norm_div_(injectionVector[64]),
.p_desc2276_p_O_FDpost_norm_div_(injectionVector[65]),
.p_desc2277_p_O_FDpost_norm_div_(injectionVector[66]),
.p_desc2278_p_O_FDpost_norm_div_(injectionVector[67]),
.p_desc2279_p_O_FDpost_norm_div_(injectionVector[68]),
.p_desc2280_p_O_FDpost_norm_div_(injectionVector[69]),
.p_desc2281_p_O_FDpost_norm_div_(injectionVector[70]),
.p_desc2282_p_O_FDpost_norm_div_(injectionVector[71]),
.p_desc2283_p_O_FDpost_norm_div_(injectionVector[72]),
.p_desc2284_p_O_FDpost_norm_div_(injectionVector[73]),
.p_desc2285_p_O_FDpost_norm_div_(injectionVector[74]),
.p_desc2286_p_O_FDpost_norm_div_(injectionVector[75]),
.p_desc2287_p_O_FDpost_norm_div_(injectionVector[76]),
.p_desc2288_p_O_FDpost_norm_div_(injectionVector[77]),
.p_desc2289_p_O_FDpost_norm_div_(injectionVector[78]),
.p_desc2290_p_O_FDpost_norm_div_(injectionVector[79]),
.p_desc2291_p_O_FDpost_norm_div_(injectionVector[80]),
.p_desc2292_p_O_FDpost_norm_div_(injectionVector[81]),
.p_desc2293_p_O_FDpost_norm_div_(injectionVector[82]),
.p_desc2294_p_O_FDpost_norm_div_(injectionVector[83]),
.p_desc2295_p_O_FDpost_norm_div_(injectionVector[84]),
.p_desc2296_p_O_FDpost_norm_div_(injectionVector[85]),
.p_desc2297_p_O_FDpost_norm_div_(injectionVector[86]),
.p_desc2298_p_O_FDpost_norm_div_(injectionVector[87]),
.p_desc2299_p_O_FDpost_norm_div_(injectionVector[88]),
.p_desc2300_p_O_FDpost_norm_div_(injectionVector[89]),
.p_desc2301_p_O_FDpost_norm_div_(injectionVector[90]),
.p_desc2302_p_O_FDpost_norm_div_(injectionVector[91]),
.p_desc2303_p_O_FDpost_norm_div_(injectionVector[92]),
.p_desc2304_p_O_FDpost_norm_div_(injectionVector[93]),
.p_desc2305_p_O_FDpost_norm_div_(injectionVector[94]),
.p_desc2306_p_O_FDpost_norm_div_(injectionVector[95]),
.p_desc2307_p_O_FDpost_norm_div_(injectionVector[96]),
.p_desc2308_p_O_FDpost_norm_div_(injectionVector[97]),
.p_desc2309_p_O_FDpost_norm_div_(injectionVector[98]),
.p_desc2310_p_O_FDpost_norm_div_(injectionVector[99]),
.p_desc2311_p_O_FDpost_norm_div_(injectionVector[100]),
.p_desc2312_p_O_FDpost_norm_div_(injectionVector[101]),
.p_desc2313_p_O_FDpost_norm_div_(injectionVector[102]),
.p_desc2314_p_O_FDpost_norm_div_(injectionVector[103]),
.p_desc2315_p_O_FDpost_norm_div_(injectionVector[104]),
.p_desc2316_p_O_FDpost_norm_div_(injectionVector[105]),
.p_desc2317_p_O_FDpost_norm_div_(injectionVector[106]),
.p_desc2318_p_O_FDpost_norm_div_(injectionVector[107]),
.p_desc2319_p_O_FDpost_norm_div_(injectionVector[108]),
.p_desc2320_p_O_FDpost_norm_div_(injectionVector[109]),
.p_desc2321_p_O_FDpost_norm_div_(injectionVector[110]),
.p_desc2322_p_O_FDpost_norm_div_(injectionVector[111]),
.p_desc2323_p_O_FDpost_norm_div_(injectionVector[112]),
.p_desc2324_p_O_FDpost_norm_div_(injectionVector[113]),
.p_desc2325_p_O_FDpost_norm_div_(injectionVector[114]),
.p_desc2326_p_O_FDpost_norm_div_(injectionVector[115]),
.p_desc2327_p_O_FDpost_norm_div_(injectionVector[116]),
.p_desc2328_p_O_FDpost_norm_div_(injectionVector[117]),
.p_desc2329_p_O_FDpost_norm_div_(injectionVector[118]),
.p_desc2330_p_O_FDpost_norm_div_(injectionVector[119]),
.p_desc2331_p_O_FDpost_norm_div_(injectionVector[120]),
.p_desc2332_p_O_FDpost_norm_div_(injectionVector[121]),
.p_desc2333_p_O_FDpost_norm_div_(injectionVector[122]),
.p_desc2334_p_O_FDpost_norm_div_(injectionVector[123]),
.p_desc2335_p_O_FDpost_norm_div_(injectionVector[124]),
.p_desc2336_p_O_FDpost_norm_div_(injectionVector[125]),
.p_desc2337_p_O_FDpost_norm_div_(injectionVector[126]),
.p_desc2338_p_O_FDpost_norm_div_(injectionVector[127]),
.p_desc2339_p_O_FDpost_norm_div_(injectionVector[128]),
.p_desc2340_p_O_FDpost_norm_div_(injectionVector[129]),
.p_desc2341_p_O_FDpost_norm_div_(injectionVector[130]),
.p_desc2342_p_O_FDpost_norm_div_(injectionVector[131]),
.p_desc2343_p_O_FDpost_norm_div_(injectionVector[132]),
.p_desc2344_p_O_FDpost_norm_div_(injectionVector[133]),
.p_desc2345_p_O_FDpost_norm_div_(injectionVector[134]),
.p_desc2346_p_O_FDpost_norm_div_(injectionVector[135]),
.p_desc2347_p_O_FDpost_norm_div_(injectionVector[136]),
.p_desc2348_p_O_FDpost_norm_div_(injectionVector[137]),
.p_desc2349_p_O_FDpost_norm_div_(injectionVector[138]),
.p_desc2350_p_O_FDpost_norm_div_(injectionVector[139]),
.p_desc2351_p_O_FDpost_norm_div_(injectionVector[140]),
.p_desc2352_p_O_FDpost_norm_div_(injectionVector[141]),
.p_desc2353_p_O_FDpost_norm_div_(injectionVector[142]),
.p_desc2354_p_O_FDpost_norm_div_(injectionVector[143]),
.p_desc2355_p_O_FDpost_norm_div_(injectionVector[144]),
.p_desc2356_p_O_FDpost_norm_div_(injectionVector[145]),
.p_desc2357_p_O_FDpost_norm_div_(injectionVector[146]),
.p_desc2358_p_O_FDpost_norm_div_(injectionVector[147]),
.p_desc2359_p_O_FDpost_norm_div_(injectionVector[148]),
.p_desc2360_p_O_FDpost_norm_div_(injectionVector[149]),
.p_desc2361_p_O_FDpost_norm_div_(injectionVector[150]),
.p_desc2362_p_O_FDpost_norm_div_(injectionVector[151]),
.p_desc2363_p_O_FDpost_norm_div_(injectionVector[152]),
.p_desc2364_p_O_FDpost_norm_div_(injectionVector[153]),
.p_desc2365_p_O_FDpost_norm_div_(injectionVector[154]),
.p_desc2366_p_O_FDpost_norm_div_(injectionVector[155]),
.p_desc2367_p_O_FDpost_norm_div_(injectionVector[156]),
.p_desc2368_p_O_FDpost_norm_div_(injectionVector[157]),
.p_desc2369_p_O_FDpost_norm_div_(injectionVector[158]),
.p_desc2370_p_O_FDpost_norm_div_(injectionVector[159]),
.p_desc2371_p_O_FDpost_norm_div_(injectionVector[160]),
.p_desc2372_p_O_FDpost_norm_div_(injectionVector[161]),
.p_desc2373_p_O_FDpost_norm_div_(injectionVector[162]),
.p_desc2374_p_O_FDpost_norm_div_(injectionVector[163]),
.p_desc2375_p_O_FDpost_norm_div_(injectionVector[164]),
.p_desc2376_p_O_FDpost_norm_div_(injectionVector[165]),
.p_desc2377_p_O_FDpost_norm_div_(injectionVector[166]),
.p_desc2378_p_O_FDpost_norm_div_(injectionVector[167]),
.p_desc2379_p_O_FDpost_norm_div_(injectionVector[168]),
.p_desc2380_p_O_FDpost_norm_div_(injectionVector[169]),
.p_desc2381_p_O_FDpost_norm_div_(injectionVector[170]),
.p_desc2382_p_O_FDpost_norm_div_(injectionVector[171]),
.p_desc2383_p_O_FDpost_norm_div_(injectionVector[172]),
.p_desc2384_p_O_FDpost_norm_div_(injectionVector[173]),
.p_desc2385_p_O_FDpost_norm_div_(injectionVector[174]),
.p_desc2386_p_O_FDpost_norm_div_(injectionVector[175]),
.p_desc2387_p_O_FDpost_norm_div_(injectionVector[176]),
.p_desc2388_p_O_FDpost_norm_div_(injectionVector[177]),
.p_desc2389_p_O_FDpost_norm_div_(injectionVector[178]),
.p_desc2390_p_O_FDpost_norm_div_(injectionVector[179]),
.p_desc2391_p_O_FDpost_norm_div_(injectionVector[180]),
.p_desc2392_p_O_FDpost_norm_div_(injectionVector[181]),
.p_desc2393_p_O_FDpost_norm_div_(injectionVector[182]),
.p_s_sign_i_Z_p_O_FDpost_norm_div_(injectionVector[183]),
.p_ine_o_Z_p_O_FDpost_norm_div_(injectionVector[184]),
.p_desc2423_p_O_FDpost_norm_div_(injectionVector[185]),
.p_desc2424_p_O_FDpost_norm_div_(injectionVector[186]),
.p_desc2425_p_O_FDpost_norm_div_(injectionVector[187]),
.p_desc2426_p_O_FDpost_norm_div_(injectionVector[188]),
.p_desc2427_p_O_FDpost_norm_div_(injectionVector[189]),
.p_desc2428_p_O_FDpost_norm_div_(injectionVector[190]),
.p_desc2429_p_O_FDpost_norm_div_(injectionVector[191]),
.p_desc2430_p_O_FDpost_norm_div_(injectionVector[192]),
.p_desc2431_p_O_FDpost_norm_div_(injectionVector[193]),
.p_desc2432_p_O_FDpost_norm_div_(injectionVector[194]),
.p_desc2464_p_O_FDpost_norm_div_(injectionVector[195]),
.p_desc2018_p_O_FDEserial_div_(injectionVector[196]),
.p_desc2019_p_O_FDEserial_div_(injectionVector[197]),
.p_desc2020_p_O_FDEserial_div_(injectionVector[198]),
.p_desc2021_p_O_FDEserial_div_(injectionVector[199]),
.p_desc2022_p_O_FDEserial_div_(injectionVector[200]),
.p_desc2023_p_O_FDEserial_div_(injectionVector[201]),
.p_desc2024_p_O_FDEserial_div_(injectionVector[202]),
.p_desc2025_p_O_FDEserial_div_(injectionVector[203]),
.p_desc2026_p_O_FDEserial_div_(injectionVector[204]),
.p_desc2027_p_O_FDEserial_div_(injectionVector[205]),
.p_desc2028_p_O_FDEserial_div_(injectionVector[206]),
.p_desc2029_p_O_FDEserial_div_(injectionVector[207]),
.p_desc2030_p_O_FDEserial_div_(injectionVector[208]),
.p_desc2031_p_O_FDEserial_div_(injectionVector[209]),
.p_desc2032_p_O_FDEserial_div_(injectionVector[210]),
.p_desc2033_p_O_FDEserial_div_(injectionVector[211]),
.p_desc2034_p_O_FDEserial_div_(injectionVector[212]),
.p_desc2035_p_O_FDEserial_div_(injectionVector[213]),
.p_desc2036_p_O_FDEserial_div_(injectionVector[214]),
.p_desc2037_p_O_FDEserial_div_(injectionVector[215]),
.p_desc2038_p_O_FDEserial_div_(injectionVector[216]),
.p_desc2039_p_O_FDEserial_div_(injectionVector[217]),
.p_desc2040_p_O_FDEserial_div_(injectionVector[218]),
.p_desc2041_p_O_FDEserial_div_(injectionVector[219]),
.p_desc2042_p_O_FDEserial_div_(injectionVector[220]),
.p_desc2043_p_O_FDEserial_div_(injectionVector[221]),
.p_desc1944_p_O_FDREserial_div_(injectionVector[222]),
.p_desc1947_p_O_FDREserial_div_(injectionVector[223]),
.p_desc2142_p_O_FDREserial_div_(injectionVector[224]),
.p_desc2143_p_O_FDREserial_div_(injectionVector[225]),
.p_desc2144_p_O_FDREserial_div_(injectionVector[226]),
.p_desc2145_p_O_FDREserial_div_(injectionVector[227]),
.p_desc2146_p_O_FDREserial_div_(injectionVector[228]),
.p_desc2147_p_O_FDREserial_div_(injectionVector[229]),
.p_desc2148_p_O_FDREserial_div_(injectionVector[230]),
.p_desc2149_p_O_FDREserial_div_(injectionVector[231]),
.p_desc2150_p_O_FDREserial_div_(injectionVector[232]),
.p_desc2151_p_O_FDREserial_div_(injectionVector[233]),
.p_desc2152_p_O_FDREserial_div_(injectionVector[234]),
.p_desc2153_p_O_FDREserial_div_(injectionVector[235]),
.p_desc2154_p_O_FDREserial_div_(injectionVector[236]),
.p_desc2155_p_O_FDREserial_div_(injectionVector[237]),
.p_desc2156_p_O_FDREserial_div_(injectionVector[238]),
.p_desc2157_p_O_FDREserial_div_(injectionVector[239]),
.p_desc2158_p_O_FDREserial_div_(injectionVector[240]),
.p_desc2159_p_O_FDREserial_div_(injectionVector[241]),
.p_desc2160_p_O_FDREserial_div_(injectionVector[242]),
.p_desc2161_p_O_FDREserial_div_(injectionVector[243]),
.p_desc2162_p_O_FDREserial_div_(injectionVector[244]),
.p_desc2163_p_O_FDREserial_div_(injectionVector[245]),
.p_desc2164_p_O_FDREserial_div_(injectionVector[246]),
.p_desc2165_p_O_FDREserial_div_(injectionVector[247]),
.p_desc2166_p_O_FDREserial_div_(injectionVector[248]),
.p_desc2167_p_O_FDREserial_div_(injectionVector[249]),
.p_desc2168_p_O_FDREserial_div_(injectionVector[250]),
.p_desc2182_p_O_FDREserial_div_(injectionVector[251]),
.p_desc2183_p_O_FDREserial_div_(injectionVector[252]),
.p_desc2184_p_O_FDREserial_div_(injectionVector[253]),
.p_desc2185_p_O_FDREserial_div_(injectionVector[254]),
.p_desc2186_p_O_FDREserial_div_(injectionVector[255]),
.p_desc2187_p_O_FDREserial_div_(injectionVector[256]),
.p_desc2188_p_O_FDREserial_div_(injectionVector[257]),
.p_desc2189_p_O_FDREserial_div_(injectionVector[258]),
.p_desc2190_p_O_FDREserial_div_(injectionVector[259]),
.p_desc2191_p_O_FDREserial_div_(injectionVector[260]),
.p_desc2192_p_O_FDREserial_div_(injectionVector[261]),
.p_desc2193_p_O_FDREserial_div_(injectionVector[262]),
.p_desc2194_p_O_FDREserial_div_(injectionVector[263]),
.p_desc2195_p_O_FDREserial_div_(injectionVector[264]),
.p_desc2196_p_O_FDREserial_div_(injectionVector[265]),
.p_desc2197_p_O_FDREserial_div_(injectionVector[266]),
.p_desc2198_p_O_FDREserial_div_(injectionVector[267]));
endmodule