
module mat_regs_WORD_WIDTH12_N4_LOG2_N2 ( .vector_in_r({\vector_in_r[0][11] , 
        \vector_in_r[0][10] , \vector_in_r[0][9] , \vector_in_r[0][8] , 
        \vector_in_r[0][7] , \vector_in_r[0][6] , \vector_in_r[0][5] , 
        \vector_in_r[0][4] , \vector_in_r[0][3] , \vector_in_r[0][2] , 
        \vector_in_r[0][1] , \vector_in_r[0][0] , \vector_in_r[1][11] , 
        \vector_in_r[1][10] , \vector_in_r[1][9] , \vector_in_r[1][8] , 
        \vector_in_r[1][7] , \vector_in_r[1][6] , \vector_in_r[1][5] , 
        \vector_in_r[1][4] , \vector_in_r[1][3] , \vector_in_r[1][2] , 
        \vector_in_r[1][1] , \vector_in_r[1][0] , \vector_in_r[2][11] , 
        \vector_in_r[2][10] , \vector_in_r[2][9] , \vector_in_r[2][8] , 
        \vector_in_r[2][7] , \vector_in_r[2][6] , \vector_in_r[2][5] , 
        \vector_in_r[2][4] , \vector_in_r[2][3] , \vector_in_r[2][2] , 
        \vector_in_r[2][1] , \vector_in_r[2][0] , \vector_in_r[3][11] , 
        \vector_in_r[3][10] , \vector_in_r[3][9] , \vector_in_r[3][8] , 
        \vector_in_r[3][7] , \vector_in_r[3][6] , \vector_in_r[3][5] , 
        \vector_in_r[3][4] , \vector_in_r[3][3] , \vector_in_r[3][2] , 
        \vector_in_r[3][1] , \vector_in_r[3][0] }), .vector_in_i({
        \vector_in_i[0][11] , \vector_in_i[0][10] , \vector_in_i[0][9] , 
        \vector_in_i[0][8] , \vector_in_i[0][7] , \vector_in_i[0][6] , 
        \vector_in_i[0][5] , \vector_in_i[0][4] , \vector_in_i[0][3] , 
        \vector_in_i[0][2] , \vector_in_i[0][1] , \vector_in_i[0][0] , 
        \vector_in_i[1][11] , \vector_in_i[1][10] , \vector_in_i[1][9] , 
        \vector_in_i[1][8] , \vector_in_i[1][7] , \vector_in_i[1][6] , 
        \vector_in_i[1][5] , \vector_in_i[1][4] , \vector_in_i[1][3] , 
        \vector_in_i[1][2] , \vector_in_i[1][1] , \vector_in_i[1][0] , 
        \vector_in_i[2][11] , \vector_in_i[2][10] , \vector_in_i[2][9] , 
        \vector_in_i[2][8] , \vector_in_i[2][7] , \vector_in_i[2][6] , 
        \vector_in_i[2][5] , \vector_in_i[2][4] , \vector_in_i[2][3] , 
        \vector_in_i[2][2] , \vector_in_i[2][1] , \vector_in_i[2][0] , 
        \vector_in_i[3][11] , \vector_in_i[3][10] , \vector_in_i[3][9] , 
        \vector_in_i[3][8] , \vector_in_i[3][7] , \vector_in_i[3][6] , 
        \vector_in_i[3][5] , \vector_in_i[3][4] , \vector_in_i[3][3] , 
        \vector_in_i[3][2] , \vector_in_i[3][1] , \vector_in_i[3][0] }), 
        w_col_sel, .vector_out_r({\vector_out_r[0][11] , \vector_out_r[0][10] , 
        \vector_out_r[0][9] , \vector_out_r[0][8] , \vector_out_r[0][7] , 
        \vector_out_r[0][6] , \vector_out_r[0][5] , \vector_out_r[0][4] , 
        \vector_out_r[0][3] , \vector_out_r[0][2] , \vector_out_r[0][1] , 
        \vector_out_r[0][0] , \vector_out_r[1][11] , \vector_out_r[1][10] , 
        \vector_out_r[1][9] , \vector_out_r[1][8] , \vector_out_r[1][7] , 
        \vector_out_r[1][6] , \vector_out_r[1][5] , \vector_out_r[1][4] , 
        \vector_out_r[1][3] , \vector_out_r[1][2] , \vector_out_r[1][1] , 
        \vector_out_r[1][0] , \vector_out_r[2][11] , \vector_out_r[2][10] , 
        \vector_out_r[2][9] , \vector_out_r[2][8] , \vector_out_r[2][7] , 
        \vector_out_r[2][6] , \vector_out_r[2][5] , \vector_out_r[2][4] , 
        \vector_out_r[2][3] , \vector_out_r[2][2] , \vector_out_r[2][1] , 
        \vector_out_r[2][0] , \vector_out_r[3][11] , \vector_out_r[3][10] , 
        \vector_out_r[3][9] , \vector_out_r[3][8] , \vector_out_r[3][7] , 
        \vector_out_r[3][6] , \vector_out_r[3][5] , \vector_out_r[3][4] , 
        \vector_out_r[3][3] , \vector_out_r[3][2] , \vector_out_r[3][1] , 
        \vector_out_r[3][0] }), .vector_out_i({\vector_out_i[0][11] , 
        \vector_out_i[0][10] , \vector_out_i[0][9] , \vector_out_i[0][8] , 
        \vector_out_i[0][7] , \vector_out_i[0][6] , \vector_out_i[0][5] , 
        \vector_out_i[0][4] , \vector_out_i[0][3] , \vector_out_i[0][2] , 
        \vector_out_i[0][1] , \vector_out_i[0][0] , \vector_out_i[1][11] , 
        \vector_out_i[1][10] , \vector_out_i[1][9] , \vector_out_i[1][8] , 
        \vector_out_i[1][7] , \vector_out_i[1][6] , \vector_out_i[1][5] , 
        \vector_out_i[1][4] , \vector_out_i[1][3] , \vector_out_i[1][2] , 
        \vector_out_i[1][1] , \vector_out_i[1][0] , \vector_out_i[2][11] , 
        \vector_out_i[2][10] , \vector_out_i[2][9] , \vector_out_i[2][8] , 
        \vector_out_i[2][7] , \vector_out_i[2][6] , \vector_out_i[2][5] , 
        \vector_out_i[2][4] , \vector_out_i[2][3] , \vector_out_i[2][2] , 
        \vector_out_i[2][1] , \vector_out_i[2][0] , \vector_out_i[3][11] , 
        \vector_out_i[3][10] , \vector_out_i[3][9] , \vector_out_i[3][8] , 
        \vector_out_i[3][7] , \vector_out_i[3][6] , \vector_out_i[3][5] , 
        \vector_out_i[3][4] , \vector_out_i[3][3] , \vector_out_i[3][2] , 
        \vector_out_i[3][1] , \vector_out_i[3][0] }), single_out_r, 
        single_out_i, col_sel, row_sel, .vector_out_r2({\vector_out_r2[0][11] , 
        \vector_out_r2[0][10] , \vector_out_r2[0][9] , \vector_out_r2[0][8] , 
        \vector_out_r2[0][7] , \vector_out_r2[0][6] , \vector_out_r2[0][5] , 
        \vector_out_r2[0][4] , \vector_out_r2[0][3] , \vector_out_r2[0][2] , 
        \vector_out_r2[0][1] , \vector_out_r2[0][0] , \vector_out_r2[1][11] , 
        \vector_out_r2[1][10] , \vector_out_r2[1][9] , \vector_out_r2[1][8] , 
        \vector_out_r2[1][7] , \vector_out_r2[1][6] , \vector_out_r2[1][5] , 
        \vector_out_r2[1][4] , \vector_out_r2[1][3] , \vector_out_r2[1][2] , 
        \vector_out_r2[1][1] , \vector_out_r2[1][0] , \vector_out_r2[2][11] , 
        \vector_out_r2[2][10] , \vector_out_r2[2][9] , \vector_out_r2[2][8] , 
        \vector_out_r2[2][7] , \vector_out_r2[2][6] , \vector_out_r2[2][5] , 
        \vector_out_r2[2][4] , \vector_out_r2[2][3] , \vector_out_r2[2][2] , 
        \vector_out_r2[2][1] , \vector_out_r2[2][0] , \vector_out_r2[3][11] , 
        \vector_out_r2[3][10] , \vector_out_r2[3][9] , \vector_out_r2[3][8] , 
        \vector_out_r2[3][7] , \vector_out_r2[3][6] , \vector_out_r2[3][5] , 
        \vector_out_r2[3][4] , \vector_out_r2[3][3] , \vector_out_r2[3][2] , 
        \vector_out_r2[3][1] , \vector_out_r2[3][0] }), .vector_out_i2({
        \vector_out_i2[0][11] , \vector_out_i2[0][10] , \vector_out_i2[0][9] , 
        \vector_out_i2[0][8] , \vector_out_i2[0][7] , \vector_out_i2[0][6] , 
        \vector_out_i2[0][5] , \vector_out_i2[0][4] , \vector_out_i2[0][3] , 
        \vector_out_i2[0][2] , \vector_out_i2[0][1] , \vector_out_i2[0][0] , 
        \vector_out_i2[1][11] , \vector_out_i2[1][10] , \vector_out_i2[1][9] , 
        \vector_out_i2[1][8] , \vector_out_i2[1][7] , \vector_out_i2[1][6] , 
        \vector_out_i2[1][5] , \vector_out_i2[1][4] , \vector_out_i2[1][3] , 
        \vector_out_i2[1][2] , \vector_out_i2[1][1] , \vector_out_i2[1][0] , 
        \vector_out_i2[2][11] , \vector_out_i2[2][10] , \vector_out_i2[2][9] , 
        \vector_out_i2[2][8] , \vector_out_i2[2][7] , \vector_out_i2[2][6] , 
        \vector_out_i2[2][5] , \vector_out_i2[2][4] , \vector_out_i2[2][3] , 
        \vector_out_i2[2][2] , \vector_out_i2[2][1] , \vector_out_i2[2][0] , 
        \vector_out_i2[3][11] , \vector_out_i2[3][10] , \vector_out_i2[3][9] , 
        \vector_out_i2[3][8] , \vector_out_i2[3][7] , \vector_out_i2[3][6] , 
        \vector_out_i2[3][5] , \vector_out_i2[3][4] , \vector_out_i2[3][3] , 
        \vector_out_i2[3][2] , \vector_out_i2[3][1] , \vector_out_i2[3][0] }), 
        single_out_r2, single_out_i2, col_sel2, row_sel2, clk, wr_enable );
  input [1:0] w_col_sel;
  output [11:0] single_out_r;
  output [11:0] single_out_i;
  input [1:0] col_sel;
  input [1:0] row_sel;
  output [11:0] single_out_r2;
  output [11:0] single_out_i2;
  input [1:0] col_sel2;
  input [1:0] row_sel2;
  input \vector_in_r[0][11] , \vector_in_r[0][10] , \vector_in_r[0][9] ,
         \vector_in_r[0][8] , \vector_in_r[0][7] , \vector_in_r[0][6] ,
         \vector_in_r[0][5] , \vector_in_r[0][4] , \vector_in_r[0][3] ,
         \vector_in_r[0][2] , \vector_in_r[0][1] , \vector_in_r[0][0] ,
         \vector_in_r[1][11] , \vector_in_r[1][10] , \vector_in_r[1][9] ,
         \vector_in_r[1][8] , \vector_in_r[1][7] , \vector_in_r[1][6] ,
         \vector_in_r[1][5] , \vector_in_r[1][4] , \vector_in_r[1][3] ,
         \vector_in_r[1][2] , \vector_in_r[1][1] , \vector_in_r[1][0] ,
         \vector_in_r[2][11] , \vector_in_r[2][10] , \vector_in_r[2][9] ,
         \vector_in_r[2][8] , \vector_in_r[2][7] , \vector_in_r[2][6] ,
         \vector_in_r[2][5] , \vector_in_r[2][4] , \vector_in_r[2][3] ,
         \vector_in_r[2][2] , \vector_in_r[2][1] , \vector_in_r[2][0] ,
         \vector_in_r[3][11] , \vector_in_r[3][10] , \vector_in_r[3][9] ,
         \vector_in_r[3][8] , \vector_in_r[3][7] , \vector_in_r[3][6] ,
         \vector_in_r[3][5] , \vector_in_r[3][4] , \vector_in_r[3][3] ,
         \vector_in_r[3][2] , \vector_in_r[3][1] , \vector_in_r[3][0] ,
         \vector_in_i[0][11] , \vector_in_i[0][10] , \vector_in_i[0][9] ,
         \vector_in_i[0][8] , \vector_in_i[0][7] , \vector_in_i[0][6] ,
         \vector_in_i[0][5] , \vector_in_i[0][4] , \vector_in_i[0][3] ,
         \vector_in_i[0][2] , \vector_in_i[0][1] , \vector_in_i[0][0] ,
         \vector_in_i[1][11] , \vector_in_i[1][10] , \vector_in_i[1][9] ,
         \vector_in_i[1][8] , \vector_in_i[1][7] , \vector_in_i[1][6] ,
         \vector_in_i[1][5] , \vector_in_i[1][4] , \vector_in_i[1][3] ,
         \vector_in_i[1][2] , \vector_in_i[1][1] , \vector_in_i[1][0] ,
         \vector_in_i[2][11] , \vector_in_i[2][10] , \vector_in_i[2][9] ,
         \vector_in_i[2][8] , \vector_in_i[2][7] , \vector_in_i[2][6] ,
         \vector_in_i[2][5] , \vector_in_i[2][4] , \vector_in_i[2][3] ,
         \vector_in_i[2][2] , \vector_in_i[2][1] , \vector_in_i[2][0] ,
         \vector_in_i[3][11] , \vector_in_i[3][10] , \vector_in_i[3][9] ,
         \vector_in_i[3][8] , \vector_in_i[3][7] , \vector_in_i[3][6] ,
         \vector_in_i[3][5] , \vector_in_i[3][4] , \vector_in_i[3][3] ,
         \vector_in_i[3][2] , \vector_in_i[3][1] , \vector_in_i[3][0] , clk,
         wr_enable;
  output \vector_out_r[0][11] , \vector_out_r[0][10] , \vector_out_r[0][9] ,
         \vector_out_r[0][8] , \vector_out_r[0][7] , \vector_out_r[0][6] ,
         \vector_out_r[0][5] , \vector_out_r[0][4] , \vector_out_r[0][3] ,
         \vector_out_r[0][2] , \vector_out_r[0][1] , \vector_out_r[0][0] ,
         \vector_out_r[1][11] , \vector_out_r[1][10] , \vector_out_r[1][9] ,
         \vector_out_r[1][8] , \vector_out_r[1][7] , \vector_out_r[1][6] ,
         \vector_out_r[1][5] , \vector_out_r[1][4] , \vector_out_r[1][3] ,
         \vector_out_r[1][2] , \vector_out_r[1][1] , \vector_out_r[1][0] ,
         \vector_out_r[2][11] , \vector_out_r[2][10] , \vector_out_r[2][9] ,
         \vector_out_r[2][8] , \vector_out_r[2][7] , \vector_out_r[2][6] ,
         \vector_out_r[2][5] , \vector_out_r[2][4] , \vector_out_r[2][3] ,
         \vector_out_r[2][2] , \vector_out_r[2][1] , \vector_out_r[2][0] ,
         \vector_out_r[3][11] , \vector_out_r[3][10] , \vector_out_r[3][9] ,
         \vector_out_r[3][8] , \vector_out_r[3][7] , \vector_out_r[3][6] ,
         \vector_out_r[3][5] , \vector_out_r[3][4] , \vector_out_r[3][3] ,
         \vector_out_r[3][2] , \vector_out_r[3][1] , \vector_out_r[3][0] ,
         \vector_out_i[0][11] , \vector_out_i[0][10] , \vector_out_i[0][9] ,
         \vector_out_i[0][8] , \vector_out_i[0][7] , \vector_out_i[0][6] ,
         \vector_out_i[0][5] , \vector_out_i[0][4] , \vector_out_i[0][3] ,
         \vector_out_i[0][2] , \vector_out_i[0][1] , \vector_out_i[0][0] ,
         \vector_out_i[1][11] , \vector_out_i[1][10] , \vector_out_i[1][9] ,
         \vector_out_i[1][8] , \vector_out_i[1][7] , \vector_out_i[1][6] ,
         \vector_out_i[1][5] , \vector_out_i[1][4] , \vector_out_i[1][3] ,
         \vector_out_i[1][2] , \vector_out_i[1][1] , \vector_out_i[1][0] ,
         \vector_out_i[2][11] , \vector_out_i[2][10] , \vector_out_i[2][9] ,
         \vector_out_i[2][8] , \vector_out_i[2][7] , \vector_out_i[2][6] ,
         \vector_out_i[2][5] , \vector_out_i[2][4] , \vector_out_i[2][3] ,
         \vector_out_i[2][2] , \vector_out_i[2][1] , \vector_out_i[2][0] ,
         \vector_out_i[3][11] , \vector_out_i[3][10] , \vector_out_i[3][9] ,
         \vector_out_i[3][8] , \vector_out_i[3][7] , \vector_out_i[3][6] ,
         \vector_out_i[3][5] , \vector_out_i[3][4] , \vector_out_i[3][3] ,
         \vector_out_i[3][2] , \vector_out_i[3][1] , \vector_out_i[3][0] ,
         \vector_out_r2[0][11] , \vector_out_r2[0][10] , \vector_out_r2[0][9] ,
         \vector_out_r2[0][8] , \vector_out_r2[0][7] , \vector_out_r2[0][6] ,
         \vector_out_r2[0][5] , \vector_out_r2[0][4] , \vector_out_r2[0][3] ,
         \vector_out_r2[0][2] , \vector_out_r2[0][1] , \vector_out_r2[0][0] ,
         \vector_out_r2[1][11] , \vector_out_r2[1][10] , \vector_out_r2[1][9] ,
         \vector_out_r2[1][8] , \vector_out_r2[1][7] , \vector_out_r2[1][6] ,
         \vector_out_r2[1][5] , \vector_out_r2[1][4] , \vector_out_r2[1][3] ,
         \vector_out_r2[1][2] , \vector_out_r2[1][1] , \vector_out_r2[1][0] ,
         \vector_out_r2[2][11] , \vector_out_r2[2][10] , \vector_out_r2[2][9] ,
         \vector_out_r2[2][8] , \vector_out_r2[2][7] , \vector_out_r2[2][6] ,
         \vector_out_r2[2][5] , \vector_out_r2[2][4] , \vector_out_r2[2][3] ,
         \vector_out_r2[2][2] , \vector_out_r2[2][1] , \vector_out_r2[2][0] ,
         \vector_out_r2[3][11] , \vector_out_r2[3][10] , \vector_out_r2[3][9] ,
         \vector_out_r2[3][8] , \vector_out_r2[3][7] , \vector_out_r2[3][6] ,
         \vector_out_r2[3][5] , \vector_out_r2[3][4] , \vector_out_r2[3][3] ,
         \vector_out_r2[3][2] , \vector_out_r2[3][1] , \vector_out_r2[3][0] ,
         \vector_out_i2[0][11] , \vector_out_i2[0][10] , \vector_out_i2[0][9] ,
         \vector_out_i2[0][8] , \vector_out_i2[0][7] , \vector_out_i2[0][6] ,
         \vector_out_i2[0][5] , \vector_out_i2[0][4] , \vector_out_i2[0][3] ,
         \vector_out_i2[0][2] , \vector_out_i2[0][1] , \vector_out_i2[0][0] ,
         \vector_out_i2[1][11] , \vector_out_i2[1][10] , \vector_out_i2[1][9] ,
         \vector_out_i2[1][8] , \vector_out_i2[1][7] , \vector_out_i2[1][6] ,
         \vector_out_i2[1][5] , \vector_out_i2[1][4] , \vector_out_i2[1][3] ,
         \vector_out_i2[1][2] , \vector_out_i2[1][1] , \vector_out_i2[1][0] ,
         \vector_out_i2[2][11] , \vector_out_i2[2][10] , \vector_out_i2[2][9] ,
         \vector_out_i2[2][8] , \vector_out_i2[2][7] , \vector_out_i2[2][6] ,
         \vector_out_i2[2][5] , \vector_out_i2[2][4] , \vector_out_i2[2][3] ,
         \vector_out_i2[2][2] , \vector_out_i2[2][1] , \vector_out_i2[2][0] ,
         \vector_out_i2[3][11] , \vector_out_i2[3][10] , \vector_out_i2[3][9] ,
         \vector_out_i2[3][8] , \vector_out_i2[3][7] , \vector_out_i2[3][6] ,
         \vector_out_i2[3][5] , \vector_out_i2[3][4] , \vector_out_i2[3][3] ,
         \vector_out_i2[3][2] , \vector_out_i2[3][1] , \vector_out_i2[3][0] ;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, \mat_r[0][0][11] ,
         \mat_r[0][0][10] , \mat_r[0][0][9] , \mat_r[0][0][8] ,
         \mat_r[0][0][7] , \mat_r[0][0][6] , \mat_r[0][0][5] ,
         \mat_r[0][0][4] , \mat_r[0][0][3] , \mat_r[0][0][2] ,
         \mat_r[0][0][1] , \mat_r[0][0][0] , \mat_r[0][1][11] ,
         \mat_r[0][1][10] , \mat_r[0][1][9] , \mat_r[0][1][8] ,
         \mat_r[0][1][7] , \mat_r[0][1][6] , \mat_r[0][1][5] ,
         \mat_r[0][1][4] , \mat_r[0][1][3] , \mat_r[0][1][2] ,
         \mat_r[0][1][1] , \mat_r[0][1][0] , \mat_r[0][2][11] ,
         \mat_r[0][2][10] , \mat_r[0][2][9] , \mat_r[0][2][8] ,
         \mat_r[0][2][7] , \mat_r[0][2][6] , \mat_r[0][2][5] ,
         \mat_r[0][2][4] , \mat_r[0][2][3] , \mat_r[0][2][2] ,
         \mat_r[0][2][1] , \mat_r[0][2][0] , \mat_r[0][3][11] ,
         \mat_r[0][3][10] , \mat_r[0][3][9] , \mat_r[0][3][8] ,
         \mat_r[0][3][7] , \mat_r[0][3][6] , \mat_r[0][3][5] ,
         \mat_r[0][3][4] , \mat_r[0][3][3] , \mat_r[0][3][2] ,
         \mat_r[0][3][1] , \mat_r[0][3][0] , \mat_r[1][0][11] ,
         \mat_r[1][0][10] , \mat_r[1][0][9] , \mat_r[1][0][8] ,
         \mat_r[1][0][7] , \mat_r[1][0][6] , \mat_r[1][0][5] ,
         \mat_r[1][0][4] , \mat_r[1][0][3] , \mat_r[1][0][2] ,
         \mat_r[1][0][1] , \mat_r[1][0][0] , \mat_r[1][1][11] ,
         \mat_r[1][1][10] , \mat_r[1][1][9] , \mat_r[1][1][8] ,
         \mat_r[1][1][7] , \mat_r[1][1][6] , \mat_r[1][1][5] ,
         \mat_r[1][1][4] , \mat_r[1][1][3] , \mat_r[1][1][2] ,
         \mat_r[1][1][1] , \mat_r[1][1][0] , \mat_r[1][2][11] ,
         \mat_r[1][2][10] , \mat_r[1][2][9] , \mat_r[1][2][8] ,
         \mat_r[1][2][7] , \mat_r[1][2][6] , \mat_r[1][2][5] ,
         \mat_r[1][2][4] , \mat_r[1][2][3] , \mat_r[1][2][2] ,
         \mat_r[1][2][1] , \mat_r[1][2][0] , \mat_r[1][3][11] ,
         \mat_r[1][3][10] , \mat_r[1][3][9] , \mat_r[1][3][8] ,
         \mat_r[1][3][7] , \mat_r[1][3][6] , \mat_r[1][3][5] ,
         \mat_r[1][3][4] , \mat_r[1][3][3] , \mat_r[1][3][2] ,
         \mat_r[1][3][1] , \mat_r[1][3][0] , \mat_r[2][0][11] ,
         \mat_r[2][0][10] , \mat_r[2][0][9] , \mat_r[2][0][8] ,
         \mat_r[2][0][7] , \mat_r[2][0][6] , \mat_r[2][0][5] ,
         \mat_r[2][0][4] , \mat_r[2][0][3] , \mat_r[2][0][2] ,
         \mat_r[2][0][1] , \mat_r[2][0][0] , \mat_r[2][1][11] ,
         \mat_r[2][1][10] , \mat_r[2][1][9] , \mat_r[2][1][8] ,
         \mat_r[2][1][7] , \mat_r[2][1][6] , \mat_r[2][1][5] ,
         \mat_r[2][1][4] , \mat_r[2][1][3] , \mat_r[2][1][2] ,
         \mat_r[2][1][1] , \mat_r[2][1][0] , \mat_r[2][2][11] ,
         \mat_r[2][2][10] , \mat_r[2][2][9] , \mat_r[2][2][8] ,
         \mat_r[2][2][7] , \mat_r[2][2][6] , \mat_r[2][2][5] ,
         \mat_r[2][2][4] , \mat_r[2][2][3] , \mat_r[2][2][2] ,
         \mat_r[2][2][1] , \mat_r[2][2][0] , \mat_r[2][3][11] ,
         \mat_r[2][3][10] , \mat_r[2][3][9] , \mat_r[2][3][8] ,
         \mat_r[2][3][7] , \mat_r[2][3][6] , \mat_r[2][3][5] ,
         \mat_r[2][3][4] , \mat_r[2][3][3] , \mat_r[2][3][2] ,
         \mat_r[2][3][1] , \mat_r[2][3][0] , \mat_r[3][0][11] ,
         \mat_r[3][0][10] , \mat_r[3][0][9] , \mat_r[3][0][8] ,
         \mat_r[3][0][7] , \mat_r[3][0][6] , \mat_r[3][0][5] ,
         \mat_r[3][0][4] , \mat_r[3][0][3] , \mat_r[3][0][2] ,
         \mat_r[3][0][1] , \mat_r[3][0][0] , \mat_r[3][1][11] ,
         \mat_r[3][1][10] , \mat_r[3][1][9] , \mat_r[3][1][8] ,
         \mat_r[3][1][7] , \mat_r[3][1][6] , \mat_r[3][1][5] ,
         \mat_r[3][1][4] , \mat_r[3][1][3] , \mat_r[3][1][2] ,
         \mat_r[3][1][1] , \mat_r[3][1][0] , \mat_r[3][2][11] ,
         \mat_r[3][2][10] , \mat_r[3][2][9] , \mat_r[3][2][8] ,
         \mat_r[3][2][7] , \mat_r[3][2][6] , \mat_r[3][2][5] ,
         \mat_r[3][2][4] , \mat_r[3][2][3] , \mat_r[3][2][2] ,
         \mat_r[3][2][1] , \mat_r[3][2][0] , \mat_r[3][3][11] ,
         \mat_r[3][3][10] , \mat_r[3][3][9] , \mat_r[3][3][8] ,
         \mat_r[3][3][7] , \mat_r[3][3][6] , \mat_r[3][3][5] ,
         \mat_r[3][3][4] , \mat_r[3][3][3] , \mat_r[3][3][2] ,
         \mat_r[3][3][1] , \mat_r[3][3][0] , \mat_i[0][0][11] ,
         \mat_i[0][0][10] , \mat_i[0][0][9] , \mat_i[0][0][8] ,
         \mat_i[0][0][7] , \mat_i[0][0][6] , \mat_i[0][0][5] ,
         \mat_i[0][0][4] , \mat_i[0][0][3] , \mat_i[0][0][2] ,
         \mat_i[0][0][1] , \mat_i[0][0][0] , \mat_i[0][1][11] ,
         \mat_i[0][1][10] , \mat_i[0][1][9] , \mat_i[0][1][8] ,
         \mat_i[0][1][7] , \mat_i[0][1][6] , \mat_i[0][1][5] ,
         \mat_i[0][1][4] , \mat_i[0][1][3] , \mat_i[0][1][2] ,
         \mat_i[0][1][1] , \mat_i[0][1][0] , \mat_i[0][2][11] ,
         \mat_i[0][2][10] , \mat_i[0][2][9] , \mat_i[0][2][8] ,
         \mat_i[0][2][7] , \mat_i[0][2][6] , \mat_i[0][2][5] ,
         \mat_i[0][2][4] , \mat_i[0][2][3] , \mat_i[0][2][2] ,
         \mat_i[0][2][1] , \mat_i[0][2][0] , \mat_i[0][3][11] ,
         \mat_i[0][3][10] , \mat_i[0][3][9] , \mat_i[0][3][8] ,
         \mat_i[0][3][7] , \mat_i[0][3][6] , \mat_i[0][3][5] ,
         \mat_i[0][3][4] , \mat_i[0][3][3] , \mat_i[0][3][2] ,
         \mat_i[0][3][1] , \mat_i[0][3][0] , \mat_i[1][0][11] ,
         \mat_i[1][0][10] , \mat_i[1][0][9] , \mat_i[1][0][8] ,
         \mat_i[1][0][7] , \mat_i[1][0][6] , \mat_i[1][0][5] ,
         \mat_i[1][0][4] , \mat_i[1][0][3] , \mat_i[1][0][2] ,
         \mat_i[1][0][1] , \mat_i[1][0][0] , \mat_i[1][1][11] ,
         \mat_i[1][1][10] , \mat_i[1][1][9] , \mat_i[1][1][8] ,
         \mat_i[1][1][7] , \mat_i[1][1][6] , \mat_i[1][1][5] ,
         \mat_i[1][1][4] , \mat_i[1][1][3] , \mat_i[1][1][2] ,
         \mat_i[1][1][1] , \mat_i[1][1][0] , \mat_i[1][2][11] ,
         \mat_i[1][2][10] , \mat_i[1][2][9] , \mat_i[1][2][8] ,
         \mat_i[1][2][7] , \mat_i[1][2][6] , \mat_i[1][2][5] ,
         \mat_i[1][2][4] , \mat_i[1][2][3] , \mat_i[1][2][2] ,
         \mat_i[1][2][1] , \mat_i[1][2][0] , \mat_i[1][3][11] ,
         \mat_i[1][3][10] , \mat_i[1][3][9] , \mat_i[1][3][8] ,
         \mat_i[1][3][7] , \mat_i[1][3][6] , \mat_i[1][3][5] ,
         \mat_i[1][3][4] , \mat_i[1][3][3] , \mat_i[1][3][2] ,
         \mat_i[1][3][1] , \mat_i[1][3][0] , \mat_i[2][0][11] ,
         \mat_i[2][0][10] , \mat_i[2][0][9] , \mat_i[2][0][8] ,
         \mat_i[2][0][7] , \mat_i[2][0][6] , \mat_i[2][0][5] ,
         \mat_i[2][0][4] , \mat_i[2][0][3] , \mat_i[2][0][2] ,
         \mat_i[2][0][1] , \mat_i[2][0][0] , \mat_i[2][1][11] ,
         \mat_i[2][1][10] , \mat_i[2][1][9] , \mat_i[2][1][8] ,
         \mat_i[2][1][7] , \mat_i[2][1][6] , \mat_i[2][1][5] ,
         \mat_i[2][1][4] , \mat_i[2][1][3] , \mat_i[2][1][2] ,
         \mat_i[2][1][1] , \mat_i[2][1][0] , \mat_i[2][2][11] ,
         \mat_i[2][2][10] , \mat_i[2][2][9] , \mat_i[2][2][8] ,
         \mat_i[2][2][7] , \mat_i[2][2][6] , \mat_i[2][2][5] ,
         \mat_i[2][2][4] , \mat_i[2][2][3] , \mat_i[2][2][2] ,
         \mat_i[2][2][1] , \mat_i[2][2][0] , \mat_i[2][3][11] ,
         \mat_i[2][3][10] , \mat_i[2][3][9] , \mat_i[2][3][8] ,
         \mat_i[2][3][7] , \mat_i[2][3][6] , \mat_i[2][3][5] ,
         \mat_i[2][3][4] , \mat_i[2][3][3] , \mat_i[2][3][2] ,
         \mat_i[2][3][1] , \mat_i[2][3][0] , \mat_i[3][0][11] ,
         \mat_i[3][0][10] , \mat_i[3][0][9] , \mat_i[3][0][8] ,
         \mat_i[3][0][7] , \mat_i[3][0][6] , \mat_i[3][0][5] ,
         \mat_i[3][0][4] , \mat_i[3][0][3] , \mat_i[3][0][2] ,
         \mat_i[3][0][1] , \mat_i[3][0][0] , \mat_i[3][1][11] ,
         \mat_i[3][1][10] , \mat_i[3][1][9] , \mat_i[3][1][8] ,
         \mat_i[3][1][7] , \mat_i[3][1][6] , \mat_i[3][1][5] ,
         \mat_i[3][1][4] , \mat_i[3][1][3] , \mat_i[3][1][2] ,
         \mat_i[3][1][1] , \mat_i[3][1][0] , \mat_i[3][2][11] ,
         \mat_i[3][2][10] , \mat_i[3][2][9] , \mat_i[3][2][8] ,
         \mat_i[3][2][7] , \mat_i[3][2][6] , \mat_i[3][2][5] ,
         \mat_i[3][2][4] , \mat_i[3][2][3] , \mat_i[3][2][2] ,
         \mat_i[3][2][1] , \mat_i[3][2][0] , \mat_i[3][3][11] ,
         \mat_i[3][3][10] , \mat_i[3][3][9] , \mat_i[3][3][8] ,
         \mat_i[3][3][7] , \mat_i[3][3][6] , \mat_i[3][3][5] ,
         \mat_i[3][3][4] , \mat_i[3][3][3] , \mat_i[3][3][2] ,
         \mat_i[3][3][1] , \mat_i[3][3][0] , n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462;
  assign N6 = col_sel[0];
  assign N7 = col_sel[1];
  assign N8 = col_sel2[0];
  assign N9 = col_sel2[1];
  assign N10 = row_sel[0];
  assign N11 = row_sel[1];
  assign N12 = row_sel2[0];
  assign N13 = row_sel2[1];

  DFFX1 \mat_i_reg[0][0][11]  ( .D(n394), .CLK(clk), .Q(\mat_i[0][0][11] ) );
  DFFX1 \mat_i_reg[0][0][10]  ( .D(n393), .CLK(clk), .Q(\mat_i[0][0][10] ) );
  DFFX1 \mat_i_reg[0][0][9]  ( .D(n392), .CLK(clk), .Q(\mat_i[0][0][9] ) );
  DFFX1 \mat_i_reg[0][0][8]  ( .D(n391), .CLK(clk), .Q(\mat_i[0][0][8] ) );
  DFFX1 \mat_i_reg[0][0][7]  ( .D(n390), .CLK(clk), .Q(\mat_i[0][0][7] ) );
  DFFX1 \mat_i_reg[0][0][6]  ( .D(n389), .CLK(clk), .Q(\mat_i[0][0][6] ) );
  DFFX1 \mat_i_reg[0][0][5]  ( .D(n388), .CLK(clk), .Q(\mat_i[0][0][5] ) );
  DFFX1 \mat_i_reg[0][0][4]  ( .D(n387), .CLK(clk), .Q(\mat_i[0][0][4] ) );
  DFFX1 \mat_i_reg[0][0][3]  ( .D(n386), .CLK(clk), .Q(\mat_i[0][0][3] ) );
  DFFX1 \mat_i_reg[0][0][2]  ( .D(n385), .CLK(clk), .Q(\mat_i[0][0][2] ) );
  DFFX1 \mat_i_reg[0][0][1]  ( .D(n384), .CLK(clk), .Q(\mat_i[0][0][1] ) );
  DFFX1 \mat_i_reg[0][0][0]  ( .D(n383), .CLK(clk), .Q(\mat_i[0][0][0] ) );
  DFFX1 \mat_i_reg[0][1][11]  ( .D(n382), .CLK(clk), .Q(\mat_i[0][1][11] ) );
  DFFX1 \mat_i_reg[0][1][10]  ( .D(n381), .CLK(clk), .Q(\mat_i[0][1][10] ) );
  DFFX1 \mat_i_reg[0][1][9]  ( .D(n380), .CLK(clk), .Q(\mat_i[0][1][9] ) );
  DFFX1 \mat_i_reg[0][1][8]  ( .D(n379), .CLK(clk), .Q(\mat_i[0][1][8] ) );
  DFFX1 \mat_i_reg[0][1][7]  ( .D(n378), .CLK(clk), .Q(\mat_i[0][1][7] ) );
  DFFX1 \mat_i_reg[0][1][6]  ( .D(n377), .CLK(clk), .Q(\mat_i[0][1][6] ) );
  DFFX1 \mat_i_reg[0][1][5]  ( .D(n376), .CLK(clk), .Q(\mat_i[0][1][5] ) );
  DFFX1 \mat_i_reg[0][1][4]  ( .D(n375), .CLK(clk), .Q(\mat_i[0][1][4] ) );
  DFFX1 \mat_i_reg[0][1][3]  ( .D(n374), .CLK(clk), .Q(\mat_i[0][1][3] ) );
  DFFX1 \mat_i_reg[0][1][2]  ( .D(n373), .CLK(clk), .Q(\mat_i[0][1][2] ) );
  DFFX1 \mat_i_reg[0][1][1]  ( .D(n372), .CLK(clk), .Q(\mat_i[0][1][1] ) );
  DFFX1 \mat_i_reg[0][1][0]  ( .D(n371), .CLK(clk), .Q(\mat_i[0][1][0] ) );
  DFFX1 \mat_i_reg[0][2][11]  ( .D(n370), .CLK(clk), .Q(\mat_i[0][2][11] ) );
  DFFX1 \mat_i_reg[0][2][10]  ( .D(n369), .CLK(clk), .Q(\mat_i[0][2][10] ) );
  DFFX1 \mat_i_reg[0][2][9]  ( .D(n368), .CLK(clk), .Q(\mat_i[0][2][9] ) );
  DFFX1 \mat_i_reg[0][2][8]  ( .D(n367), .CLK(clk), .Q(\mat_i[0][2][8] ) );
  DFFX1 \mat_i_reg[0][2][7]  ( .D(n366), .CLK(clk), .Q(\mat_i[0][2][7] ) );
  DFFX1 \mat_i_reg[0][2][6]  ( .D(n365), .CLK(clk), .Q(\mat_i[0][2][6] ) );
  DFFX1 \mat_i_reg[0][2][5]  ( .D(n364), .CLK(clk), .Q(\mat_i[0][2][5] ) );
  DFFX1 \mat_i_reg[0][2][4]  ( .D(n363), .CLK(clk), .Q(\mat_i[0][2][4] ) );
  DFFX1 \mat_i_reg[0][2][3]  ( .D(n362), .CLK(clk), .Q(\mat_i[0][2][3] ) );
  DFFX1 \mat_i_reg[0][2][2]  ( .D(n361), .CLK(clk), .Q(\mat_i[0][2][2] ) );
  DFFX1 \mat_i_reg[0][2][1]  ( .D(n360), .CLK(clk), .Q(\mat_i[0][2][1] ) );
  DFFX1 \mat_i_reg[0][2][0]  ( .D(n359), .CLK(clk), .Q(\mat_i[0][2][0] ) );
  DFFX1 \mat_i_reg[0][3][11]  ( .D(n358), .CLK(clk), .Q(\mat_i[0][3][11] ) );
  DFFX1 \mat_i_reg[0][3][10]  ( .D(n357), .CLK(clk), .Q(\mat_i[0][3][10] ) );
  DFFX1 \mat_i_reg[0][3][9]  ( .D(n356), .CLK(clk), .Q(\mat_i[0][3][9] ) );
  DFFX1 \mat_i_reg[0][3][8]  ( .D(n355), .CLK(clk), .Q(\mat_i[0][3][8] ) );
  DFFX1 \mat_i_reg[0][3][7]  ( .D(n354), .CLK(clk), .Q(\mat_i[0][3][7] ) );
  DFFX1 \mat_i_reg[0][3][6]  ( .D(n353), .CLK(clk), .Q(\mat_i[0][3][6] ) );
  DFFX1 \mat_i_reg[0][3][5]  ( .D(n352), .CLK(clk), .Q(\mat_i[0][3][5] ) );
  DFFX1 \mat_i_reg[0][3][4]  ( .D(n351), .CLK(clk), .Q(\mat_i[0][3][4] ) );
  DFFX1 \mat_i_reg[0][3][3]  ( .D(n350), .CLK(clk), .Q(\mat_i[0][3][3] ) );
  DFFX1 \mat_i_reg[0][3][2]  ( .D(n349), .CLK(clk), .Q(\mat_i[0][3][2] ) );
  DFFX1 \mat_i_reg[0][3][1]  ( .D(n348), .CLK(clk), .Q(\mat_i[0][3][1] ) );
  DFFX1 \mat_i_reg[0][3][0]  ( .D(n347), .CLK(clk), .Q(\mat_i[0][3][0] ) );
  DFFX1 \mat_i_reg[1][0][11]  ( .D(n346), .CLK(clk), .Q(\mat_i[1][0][11] ) );
  DFFX1 \mat_i_reg[1][0][10]  ( .D(n345), .CLK(clk), .Q(\mat_i[1][0][10] ) );
  DFFX1 \mat_i_reg[1][0][9]  ( .D(n344), .CLK(clk), .Q(\mat_i[1][0][9] ) );
  DFFX1 \mat_i_reg[1][0][8]  ( .D(n343), .CLK(clk), .Q(\mat_i[1][0][8] ) );
  DFFX1 \mat_i_reg[1][0][7]  ( .D(n342), .CLK(clk), .Q(\mat_i[1][0][7] ) );
  DFFX1 \mat_i_reg[1][0][6]  ( .D(n341), .CLK(clk), .Q(\mat_i[1][0][6] ) );
  DFFX1 \mat_i_reg[1][0][5]  ( .D(n340), .CLK(clk), .Q(\mat_i[1][0][5] ) );
  DFFX1 \mat_i_reg[1][0][4]  ( .D(n339), .CLK(clk), .Q(\mat_i[1][0][4] ) );
  DFFX1 \mat_i_reg[1][0][3]  ( .D(n338), .CLK(clk), .Q(\mat_i[1][0][3] ) );
  DFFX1 \mat_i_reg[1][0][2]  ( .D(n337), .CLK(clk), .Q(\mat_i[1][0][2] ) );
  DFFX1 \mat_i_reg[1][0][1]  ( .D(n336), .CLK(clk), .Q(\mat_i[1][0][1] ) );
  DFFX1 \mat_i_reg[1][0][0]  ( .D(n335), .CLK(clk), .Q(\mat_i[1][0][0] ) );
  DFFX1 \mat_i_reg[1][1][11]  ( .D(n334), .CLK(clk), .Q(\mat_i[1][1][11] ) );
  DFFX1 \mat_i_reg[1][1][10]  ( .D(n333), .CLK(clk), .Q(\mat_i[1][1][10] ) );
  DFFX1 \mat_i_reg[1][1][9]  ( .D(n332), .CLK(clk), .Q(\mat_i[1][1][9] ) );
  DFFX1 \mat_i_reg[1][1][8]  ( .D(n331), .CLK(clk), .Q(\mat_i[1][1][8] ) );
  DFFX1 \mat_i_reg[1][1][7]  ( .D(n330), .CLK(clk), .Q(\mat_i[1][1][7] ) );
  DFFX1 \mat_i_reg[1][1][6]  ( .D(n329), .CLK(clk), .Q(\mat_i[1][1][6] ) );
  DFFX1 \mat_i_reg[1][1][5]  ( .D(n328), .CLK(clk), .Q(\mat_i[1][1][5] ) );
  DFFX1 \mat_i_reg[1][1][4]  ( .D(n327), .CLK(clk), .Q(\mat_i[1][1][4] ) );
  DFFX1 \mat_i_reg[1][1][3]  ( .D(n326), .CLK(clk), .Q(\mat_i[1][1][3] ) );
  DFFX1 \mat_i_reg[1][1][2]  ( .D(n325), .CLK(clk), .Q(\mat_i[1][1][2] ) );
  DFFX1 \mat_i_reg[1][1][1]  ( .D(n324), .CLK(clk), .Q(\mat_i[1][1][1] ) );
  DFFX1 \mat_i_reg[1][1][0]  ( .D(n323), .CLK(clk), .Q(\mat_i[1][1][0] ) );
  DFFX1 \mat_i_reg[1][2][11]  ( .D(n322), .CLK(clk), .Q(\mat_i[1][2][11] ) );
  DFFX1 \mat_i_reg[1][2][10]  ( .D(n321), .CLK(clk), .Q(\mat_i[1][2][10] ) );
  DFFX1 \mat_i_reg[1][2][9]  ( .D(n320), .CLK(clk), .Q(\mat_i[1][2][9] ) );
  DFFX1 \mat_i_reg[1][2][8]  ( .D(n319), .CLK(clk), .Q(\mat_i[1][2][8] ) );
  DFFX1 \mat_i_reg[1][2][7]  ( .D(n318), .CLK(clk), .Q(\mat_i[1][2][7] ) );
  DFFX1 \mat_i_reg[1][2][6]  ( .D(n317), .CLK(clk), .Q(\mat_i[1][2][6] ) );
  DFFX1 \mat_i_reg[1][2][5]  ( .D(n316), .CLK(clk), .Q(\mat_i[1][2][5] ) );
  DFFX1 \mat_i_reg[1][2][4]  ( .D(n315), .CLK(clk), .Q(\mat_i[1][2][4] ) );
  DFFX1 \mat_i_reg[1][2][3]  ( .D(n314), .CLK(clk), .Q(\mat_i[1][2][3] ) );
  DFFX1 \mat_i_reg[1][2][2]  ( .D(n313), .CLK(clk), .Q(\mat_i[1][2][2] ) );
  DFFX1 \mat_i_reg[1][2][1]  ( .D(n312), .CLK(clk), .Q(\mat_i[1][2][1] ) );
  DFFX1 \mat_i_reg[1][2][0]  ( .D(n311), .CLK(clk), .Q(\mat_i[1][2][0] ) );
  DFFX1 \mat_i_reg[1][3][11]  ( .D(n310), .CLK(clk), .Q(\mat_i[1][3][11] ) );
  DFFX1 \mat_i_reg[1][3][10]  ( .D(n309), .CLK(clk), .Q(\mat_i[1][3][10] ) );
  DFFX1 \mat_i_reg[1][3][9]  ( .D(n308), .CLK(clk), .Q(\mat_i[1][3][9] ) );
  DFFX1 \mat_i_reg[1][3][8]  ( .D(n307), .CLK(clk), .Q(\mat_i[1][3][8] ) );
  DFFX1 \mat_i_reg[1][3][7]  ( .D(n306), .CLK(clk), .Q(\mat_i[1][3][7] ) );
  DFFX1 \mat_i_reg[1][3][6]  ( .D(n305), .CLK(clk), .Q(\mat_i[1][3][6] ) );
  DFFX1 \mat_i_reg[1][3][5]  ( .D(n304), .CLK(clk), .Q(\mat_i[1][3][5] ) );
  DFFX1 \mat_i_reg[1][3][4]  ( .D(n303), .CLK(clk), .Q(\mat_i[1][3][4] ) );
  DFFX1 \mat_i_reg[1][3][3]  ( .D(n302), .CLK(clk), .Q(\mat_i[1][3][3] ) );
  DFFX1 \mat_i_reg[1][3][2]  ( .D(n301), .CLK(clk), .Q(\mat_i[1][3][2] ) );
  DFFX1 \mat_i_reg[1][3][1]  ( .D(n300), .CLK(clk), .Q(\mat_i[1][3][1] ) );
  DFFX1 \mat_i_reg[1][3][0]  ( .D(n299), .CLK(clk), .Q(\mat_i[1][3][0] ) );
  DFFX1 \mat_i_reg[2][0][11]  ( .D(n298), .CLK(clk), .Q(\mat_i[2][0][11] ) );
  DFFX1 \mat_i_reg[2][0][10]  ( .D(n297), .CLK(clk), .Q(\mat_i[2][0][10] ) );
  DFFX1 \mat_i_reg[2][0][9]  ( .D(n296), .CLK(clk), .Q(\mat_i[2][0][9] ) );
  DFFX1 \mat_i_reg[2][0][8]  ( .D(n295), .CLK(clk), .Q(\mat_i[2][0][8] ) );
  DFFX1 \mat_i_reg[2][0][7]  ( .D(n294), .CLK(clk), .Q(\mat_i[2][0][7] ) );
  DFFX1 \mat_i_reg[2][0][6]  ( .D(n293), .CLK(clk), .Q(\mat_i[2][0][6] ) );
  DFFX1 \mat_i_reg[2][0][5]  ( .D(n292), .CLK(clk), .Q(\mat_i[2][0][5] ) );
  DFFX1 \mat_i_reg[2][0][4]  ( .D(n291), .CLK(clk), .Q(\mat_i[2][0][4] ) );
  DFFX1 \mat_i_reg[2][0][3]  ( .D(n290), .CLK(clk), .Q(\mat_i[2][0][3] ) );
  DFFX1 \mat_i_reg[2][0][2]  ( .D(n289), .CLK(clk), .Q(\mat_i[2][0][2] ) );
  DFFX1 \mat_i_reg[2][0][1]  ( .D(n288), .CLK(clk), .Q(\mat_i[2][0][1] ) );
  DFFX1 \mat_i_reg[2][0][0]  ( .D(n287), .CLK(clk), .Q(\mat_i[2][0][0] ) );
  DFFX1 \mat_i_reg[2][1][11]  ( .D(n286), .CLK(clk), .Q(\mat_i[2][1][11] ) );
  DFFX1 \mat_i_reg[2][1][10]  ( .D(n285), .CLK(clk), .Q(\mat_i[2][1][10] ) );
  DFFX1 \mat_i_reg[2][1][9]  ( .D(n284), .CLK(clk), .Q(\mat_i[2][1][9] ) );
  DFFX1 \mat_i_reg[2][1][8]  ( .D(n283), .CLK(clk), .Q(\mat_i[2][1][8] ) );
  DFFX1 \mat_i_reg[2][1][7]  ( .D(n282), .CLK(clk), .Q(\mat_i[2][1][7] ) );
  DFFX1 \mat_i_reg[2][1][6]  ( .D(n281), .CLK(clk), .Q(\mat_i[2][1][6] ) );
  DFFX1 \mat_i_reg[2][1][5]  ( .D(n280), .CLK(clk), .Q(\mat_i[2][1][5] ) );
  DFFX1 \mat_i_reg[2][1][4]  ( .D(n279), .CLK(clk), .Q(\mat_i[2][1][4] ) );
  DFFX1 \mat_i_reg[2][1][3]  ( .D(n278), .CLK(clk), .Q(\mat_i[2][1][3] ) );
  DFFX1 \mat_i_reg[2][1][2]  ( .D(n277), .CLK(clk), .Q(\mat_i[2][1][2] ) );
  DFFX1 \mat_i_reg[2][1][1]  ( .D(n276), .CLK(clk), .Q(\mat_i[2][1][1] ) );
  DFFX1 \mat_i_reg[2][1][0]  ( .D(n275), .CLK(clk), .Q(\mat_i[2][1][0] ) );
  DFFX1 \mat_i_reg[2][2][11]  ( .D(n274), .CLK(clk), .Q(\mat_i[2][2][11] ) );
  DFFX1 \mat_i_reg[2][2][10]  ( .D(n273), .CLK(clk), .Q(\mat_i[2][2][10] ) );
  DFFX1 \mat_i_reg[2][2][9]  ( .D(n272), .CLK(clk), .Q(\mat_i[2][2][9] ) );
  DFFX1 \mat_i_reg[2][2][8]  ( .D(n271), .CLK(clk), .Q(\mat_i[2][2][8] ) );
  DFFX1 \mat_i_reg[2][2][7]  ( .D(n270), .CLK(clk), .Q(\mat_i[2][2][7] ) );
  DFFX1 \mat_i_reg[2][2][6]  ( .D(n269), .CLK(clk), .Q(\mat_i[2][2][6] ) );
  DFFX1 \mat_i_reg[2][2][5]  ( .D(n268), .CLK(clk), .Q(\mat_i[2][2][5] ) );
  DFFX1 \mat_i_reg[2][2][4]  ( .D(n267), .CLK(clk), .Q(\mat_i[2][2][4] ) );
  DFFX1 \mat_i_reg[2][2][3]  ( .D(n266), .CLK(clk), .Q(\mat_i[2][2][3] ) );
  DFFX1 \mat_i_reg[2][2][2]  ( .D(n265), .CLK(clk), .Q(\mat_i[2][2][2] ) );
  DFFX1 \mat_i_reg[2][2][1]  ( .D(n264), .CLK(clk), .Q(\mat_i[2][2][1] ) );
  DFFX1 \mat_i_reg[2][2][0]  ( .D(n263), .CLK(clk), .Q(\mat_i[2][2][0] ) );
  DFFX1 \mat_i_reg[2][3][11]  ( .D(n262), .CLK(clk), .Q(\mat_i[2][3][11] ) );
  DFFX1 \mat_i_reg[2][3][10]  ( .D(n261), .CLK(clk), .Q(\mat_i[2][3][10] ) );
  DFFX1 \mat_i_reg[2][3][9]  ( .D(n260), .CLK(clk), .Q(\mat_i[2][3][9] ) );
  DFFX1 \mat_i_reg[2][3][8]  ( .D(n259), .CLK(clk), .Q(\mat_i[2][3][8] ) );
  DFFX1 \mat_i_reg[2][3][7]  ( .D(n258), .CLK(clk), .Q(\mat_i[2][3][7] ) );
  DFFX1 \mat_i_reg[2][3][6]  ( .D(n257), .CLK(clk), .Q(\mat_i[2][3][6] ) );
  DFFX1 \mat_i_reg[2][3][5]  ( .D(n256), .CLK(clk), .Q(\mat_i[2][3][5] ) );
  DFFX1 \mat_i_reg[2][3][4]  ( .D(n255), .CLK(clk), .Q(\mat_i[2][3][4] ) );
  DFFX1 \mat_i_reg[2][3][3]  ( .D(n254), .CLK(clk), .Q(\mat_i[2][3][3] ) );
  DFFX1 \mat_i_reg[2][3][2]  ( .D(n253), .CLK(clk), .Q(\mat_i[2][3][2] ) );
  DFFX1 \mat_i_reg[2][3][1]  ( .D(n252), .CLK(clk), .Q(\mat_i[2][3][1] ) );
  DFFX1 \mat_i_reg[2][3][0]  ( .D(n251), .CLK(clk), .Q(\mat_i[2][3][0] ) );
  DFFX1 \mat_i_reg[3][0][11]  ( .D(n250), .CLK(clk), .Q(\mat_i[3][0][11] ) );
  DFFX1 \mat_i_reg[3][0][10]  ( .D(n249), .CLK(clk), .Q(\mat_i[3][0][10] ) );
  DFFX1 \mat_i_reg[3][0][9]  ( .D(n248), .CLK(clk), .Q(\mat_i[3][0][9] ) );
  DFFX1 \mat_i_reg[3][0][8]  ( .D(n247), .CLK(clk), .Q(\mat_i[3][0][8] ) );
  DFFX1 \mat_i_reg[3][0][7]  ( .D(n246), .CLK(clk), .Q(\mat_i[3][0][7] ) );
  DFFX1 \mat_i_reg[3][0][6]  ( .D(n245), .CLK(clk), .Q(\mat_i[3][0][6] ) );
  DFFX1 \mat_i_reg[3][0][5]  ( .D(n244), .CLK(clk), .Q(\mat_i[3][0][5] ) );
  DFFX1 \mat_i_reg[3][0][4]  ( .D(n243), .CLK(clk), .Q(\mat_i[3][0][4] ) );
  DFFX1 \mat_i_reg[3][0][3]  ( .D(n242), .CLK(clk), .Q(\mat_i[3][0][3] ) );
  DFFX1 \mat_i_reg[3][0][2]  ( .D(n241), .CLK(clk), .Q(\mat_i[3][0][2] ) );
  DFFX1 \mat_i_reg[3][0][1]  ( .D(n240), .CLK(clk), .Q(\mat_i[3][0][1] ) );
  DFFX1 \mat_i_reg[3][0][0]  ( .D(n239), .CLK(clk), .Q(\mat_i[3][0][0] ) );
  DFFX1 \mat_i_reg[3][1][11]  ( .D(n238), .CLK(clk), .Q(\mat_i[3][1][11] ) );
  DFFX1 \mat_i_reg[3][1][10]  ( .D(n237), .CLK(clk), .Q(\mat_i[3][1][10] ) );
  DFFX1 \mat_i_reg[3][1][9]  ( .D(n236), .CLK(clk), .Q(\mat_i[3][1][9] ) );
  DFFX1 \mat_i_reg[3][1][8]  ( .D(n235), .CLK(clk), .Q(\mat_i[3][1][8] ) );
  DFFX1 \mat_i_reg[3][1][7]  ( .D(n234), .CLK(clk), .Q(\mat_i[3][1][7] ) );
  DFFX1 \mat_i_reg[3][1][6]  ( .D(n233), .CLK(clk), .Q(\mat_i[3][1][6] ) );
  DFFX1 \mat_i_reg[3][1][5]  ( .D(n232), .CLK(clk), .Q(\mat_i[3][1][5] ) );
  DFFX1 \mat_i_reg[3][1][4]  ( .D(n231), .CLK(clk), .Q(\mat_i[3][1][4] ) );
  DFFX1 \mat_i_reg[3][1][3]  ( .D(n230), .CLK(clk), .Q(\mat_i[3][1][3] ) );
  DFFX1 \mat_i_reg[3][1][2]  ( .D(n229), .CLK(clk), .Q(\mat_i[3][1][2] ) );
  DFFX1 \mat_i_reg[3][1][1]  ( .D(n228), .CLK(clk), .Q(\mat_i[3][1][1] ) );
  DFFX1 \mat_i_reg[3][1][0]  ( .D(n227), .CLK(clk), .Q(\mat_i[3][1][0] ) );
  DFFX1 \mat_i_reg[3][2][11]  ( .D(n226), .CLK(clk), .Q(\mat_i[3][2][11] ) );
  DFFX1 \mat_i_reg[3][2][10]  ( .D(n225), .CLK(clk), .Q(\mat_i[3][2][10] ) );
  DFFX1 \mat_i_reg[3][2][9]  ( .D(n224), .CLK(clk), .Q(\mat_i[3][2][9] ) );
  DFFX1 \mat_i_reg[3][2][8]  ( .D(n223), .CLK(clk), .Q(\mat_i[3][2][8] ) );
  DFFX1 \mat_i_reg[3][2][7]  ( .D(n222), .CLK(clk), .Q(\mat_i[3][2][7] ) );
  DFFX1 \mat_i_reg[3][2][6]  ( .D(n221), .CLK(clk), .Q(\mat_i[3][2][6] ) );
  DFFX1 \mat_i_reg[3][2][5]  ( .D(n220), .CLK(clk), .Q(\mat_i[3][2][5] ) );
  DFFX1 \mat_i_reg[3][2][4]  ( .D(n219), .CLK(clk), .Q(\mat_i[3][2][4] ) );
  DFFX1 \mat_i_reg[3][2][3]  ( .D(n218), .CLK(clk), .Q(\mat_i[3][2][3] ) );
  DFFX1 \mat_i_reg[3][2][2]  ( .D(n217), .CLK(clk), .Q(\mat_i[3][2][2] ) );
  DFFX1 \mat_i_reg[3][2][1]  ( .D(n216), .CLK(clk), .Q(\mat_i[3][2][1] ) );
  DFFX1 \mat_i_reg[3][2][0]  ( .D(n215), .CLK(clk), .Q(\mat_i[3][2][0] ) );
  DFFX1 \mat_i_reg[3][3][11]  ( .D(n214), .CLK(clk), .Q(\mat_i[3][3][11] ) );
  DFFX1 \mat_i_reg[3][3][10]  ( .D(n213), .CLK(clk), .Q(\mat_i[3][3][10] ) );
  DFFX1 \mat_i_reg[3][3][9]  ( .D(n212), .CLK(clk), .Q(\mat_i[3][3][9] ) );
  DFFX1 \mat_i_reg[3][3][8]  ( .D(n211), .CLK(clk), .Q(\mat_i[3][3][8] ) );
  DFFX1 \mat_i_reg[3][3][7]  ( .D(n210), .CLK(clk), .Q(\mat_i[3][3][7] ) );
  DFFX1 \mat_i_reg[3][3][6]  ( .D(n209), .CLK(clk), .Q(\mat_i[3][3][6] ) );
  DFFX1 \mat_i_reg[3][3][5]  ( .D(n208), .CLK(clk), .Q(\mat_i[3][3][5] ) );
  DFFX1 \mat_i_reg[3][3][4]  ( .D(n207), .CLK(clk), .Q(\mat_i[3][3][4] ) );
  DFFX1 \mat_i_reg[3][3][3]  ( .D(n206), .CLK(clk), .Q(\mat_i[3][3][3] ) );
  DFFX1 \mat_i_reg[3][3][2]  ( .D(n205), .CLK(clk), .Q(\mat_i[3][3][2] ) );
  DFFX1 \mat_i_reg[3][3][1]  ( .D(n204), .CLK(clk), .Q(\mat_i[3][3][1] ) );
  DFFX1 \mat_i_reg[3][3][0]  ( .D(n203), .CLK(clk), .Q(\mat_i[3][3][0] ) );
  DFFX1 \mat_r_reg[0][0][11]  ( .D(n202), .CLK(clk), .Q(\mat_r[0][0][11] ) );
  DFFX1 \mat_r_reg[0][0][10]  ( .D(n201), .CLK(clk), .Q(\mat_r[0][0][10] ) );
  DFFX1 \mat_r_reg[0][0][9]  ( .D(n200), .CLK(clk), .Q(\mat_r[0][0][9] ) );
  DFFX1 \mat_r_reg[0][0][8]  ( .D(n199), .CLK(clk), .Q(\mat_r[0][0][8] ) );
  DFFX1 \mat_r_reg[0][0][7]  ( .D(n198), .CLK(clk), .Q(\mat_r[0][0][7] ) );
  DFFX1 \mat_r_reg[0][0][6]  ( .D(n197), .CLK(clk), .Q(\mat_r[0][0][6] ) );
  DFFX1 \mat_r_reg[0][0][5]  ( .D(n196), .CLK(clk), .Q(\mat_r[0][0][5] ) );
  DFFX1 \mat_r_reg[0][0][4]  ( .D(n195), .CLK(clk), .Q(\mat_r[0][0][4] ) );
  DFFX1 \mat_r_reg[0][0][3]  ( .D(n194), .CLK(clk), .Q(\mat_r[0][0][3] ) );
  DFFX1 \mat_r_reg[0][0][2]  ( .D(n193), .CLK(clk), .Q(\mat_r[0][0][2] ) );
  DFFX1 \mat_r_reg[0][0][1]  ( .D(n192), .CLK(clk), .Q(\mat_r[0][0][1] ) );
  DFFX1 \mat_r_reg[0][0][0]  ( .D(n191), .CLK(clk), .Q(\mat_r[0][0][0] ) );
  DFFX1 \mat_r_reg[0][1][11]  ( .D(n190), .CLK(clk), .Q(\mat_r[0][1][11] ) );
  DFFX1 \mat_r_reg[0][1][10]  ( .D(n189), .CLK(clk), .Q(\mat_r[0][1][10] ) );
  DFFX1 \mat_r_reg[0][1][9]  ( .D(n188), .CLK(clk), .Q(\mat_r[0][1][9] ) );
  DFFX1 \mat_r_reg[0][1][8]  ( .D(n187), .CLK(clk), .Q(\mat_r[0][1][8] ) );
  DFFX1 \mat_r_reg[0][1][7]  ( .D(n186), .CLK(clk), .Q(\mat_r[0][1][7] ) );
  DFFX1 \mat_r_reg[0][1][6]  ( .D(n185), .CLK(clk), .Q(\mat_r[0][1][6] ) );
  DFFX1 \mat_r_reg[0][1][5]  ( .D(n184), .CLK(clk), .Q(\mat_r[0][1][5] ) );
  DFFX1 \mat_r_reg[0][1][4]  ( .D(n183), .CLK(clk), .Q(\mat_r[0][1][4] ) );
  DFFX1 \mat_r_reg[0][1][3]  ( .D(n182), .CLK(clk), .Q(\mat_r[0][1][3] ) );
  DFFX1 \mat_r_reg[0][1][2]  ( .D(n181), .CLK(clk), .Q(\mat_r[0][1][2] ) );
  DFFX1 \mat_r_reg[0][1][1]  ( .D(n180), .CLK(clk), .Q(\mat_r[0][1][1] ) );
  DFFX1 \mat_r_reg[0][1][0]  ( .D(n179), .CLK(clk), .Q(\mat_r[0][1][0] ) );
  DFFX1 \mat_r_reg[0][2][11]  ( .D(n178), .CLK(clk), .Q(\mat_r[0][2][11] ) );
  DFFX1 \mat_r_reg[0][2][10]  ( .D(n177), .CLK(clk), .Q(\mat_r[0][2][10] ) );
  DFFX1 \mat_r_reg[0][2][9]  ( .D(n176), .CLK(clk), .Q(\mat_r[0][2][9] ) );
  DFFX1 \mat_r_reg[0][2][8]  ( .D(n175), .CLK(clk), .Q(\mat_r[0][2][8] ) );
  DFFX1 \mat_r_reg[0][2][7]  ( .D(n174), .CLK(clk), .Q(\mat_r[0][2][7] ) );
  DFFX1 \mat_r_reg[0][2][6]  ( .D(n173), .CLK(clk), .Q(\mat_r[0][2][6] ) );
  DFFX1 \mat_r_reg[0][2][5]  ( .D(n172), .CLK(clk), .Q(\mat_r[0][2][5] ) );
  DFFX1 \mat_r_reg[0][2][4]  ( .D(n171), .CLK(clk), .Q(\mat_r[0][2][4] ) );
  DFFX1 \mat_r_reg[0][2][3]  ( .D(n170), .CLK(clk), .Q(\mat_r[0][2][3] ) );
  DFFX1 \mat_r_reg[0][2][2]  ( .D(n169), .CLK(clk), .Q(\mat_r[0][2][2] ) );
  DFFX1 \mat_r_reg[0][2][1]  ( .D(n168), .CLK(clk), .Q(\mat_r[0][2][1] ) );
  DFFX1 \mat_r_reg[0][2][0]  ( .D(n167), .CLK(clk), .Q(\mat_r[0][2][0] ) );
  DFFX1 \mat_r_reg[0][3][11]  ( .D(n166), .CLK(clk), .Q(\mat_r[0][3][11] ) );
  DFFX1 \mat_r_reg[0][3][10]  ( .D(n165), .CLK(clk), .Q(\mat_r[0][3][10] ) );
  DFFX1 \mat_r_reg[0][3][9]  ( .D(n164), .CLK(clk), .Q(\mat_r[0][3][9] ) );
  DFFX1 \mat_r_reg[0][3][8]  ( .D(n163), .CLK(clk), .Q(\mat_r[0][3][8] ) );
  DFFX1 \mat_r_reg[0][3][7]  ( .D(n162), .CLK(clk), .Q(\mat_r[0][3][7] ) );
  DFFX1 \mat_r_reg[0][3][6]  ( .D(n161), .CLK(clk), .Q(\mat_r[0][3][6] ) );
  DFFX1 \mat_r_reg[0][3][5]  ( .D(n160), .CLK(clk), .Q(\mat_r[0][3][5] ) );
  DFFX1 \mat_r_reg[0][3][4]  ( .D(n159), .CLK(clk), .Q(\mat_r[0][3][4] ) );
  DFFX1 \mat_r_reg[0][3][3]  ( .D(n158), .CLK(clk), .Q(\mat_r[0][3][3] ) );
  DFFX1 \mat_r_reg[0][3][2]  ( .D(n157), .CLK(clk), .Q(\mat_r[0][3][2] ) );
  DFFX1 \mat_r_reg[0][3][1]  ( .D(n156), .CLK(clk), .Q(\mat_r[0][3][1] ) );
  DFFX1 \mat_r_reg[0][3][0]  ( .D(n155), .CLK(clk), .Q(\mat_r[0][3][0] ) );
  DFFX1 \mat_r_reg[1][0][11]  ( .D(n154), .CLK(clk), .Q(\mat_r[1][0][11] ) );
  DFFX1 \mat_r_reg[1][0][10]  ( .D(n153), .CLK(clk), .Q(\mat_r[1][0][10] ) );
  DFFX1 \mat_r_reg[1][0][9]  ( .D(n152), .CLK(clk), .Q(\mat_r[1][0][9] ) );
  DFFX1 \mat_r_reg[1][0][8]  ( .D(n151), .CLK(clk), .Q(\mat_r[1][0][8] ) );
  DFFX1 \mat_r_reg[1][0][7]  ( .D(n150), .CLK(clk), .Q(\mat_r[1][0][7] ) );
  DFFX1 \mat_r_reg[1][0][6]  ( .D(n149), .CLK(clk), .Q(\mat_r[1][0][6] ) );
  DFFX1 \mat_r_reg[1][0][5]  ( .D(n148), .CLK(clk), .Q(\mat_r[1][0][5] ) );
  DFFX1 \mat_r_reg[1][0][4]  ( .D(n147), .CLK(clk), .Q(\mat_r[1][0][4] ) );
  DFFX1 \mat_r_reg[1][0][3]  ( .D(n146), .CLK(clk), .Q(\mat_r[1][0][3] ) );
  DFFX1 \mat_r_reg[1][0][2]  ( .D(n145), .CLK(clk), .Q(\mat_r[1][0][2] ) );
  DFFX1 \mat_r_reg[1][0][1]  ( .D(n144), .CLK(clk), .Q(\mat_r[1][0][1] ) );
  DFFX1 \mat_r_reg[1][0][0]  ( .D(n143), .CLK(clk), .Q(\mat_r[1][0][0] ) );
  DFFX1 \mat_r_reg[1][1][11]  ( .D(n142), .CLK(clk), .Q(\mat_r[1][1][11] ) );
  DFFX1 \mat_r_reg[1][1][10]  ( .D(n141), .CLK(clk), .Q(\mat_r[1][1][10] ) );
  DFFX1 \mat_r_reg[1][1][9]  ( .D(n140), .CLK(clk), .Q(\mat_r[1][1][9] ) );
  DFFX1 \mat_r_reg[1][1][8]  ( .D(n139), .CLK(clk), .Q(\mat_r[1][1][8] ) );
  DFFX1 \mat_r_reg[1][1][7]  ( .D(n138), .CLK(clk), .Q(\mat_r[1][1][7] ) );
  DFFX1 \mat_r_reg[1][1][6]  ( .D(n137), .CLK(clk), .Q(\mat_r[1][1][6] ) );
  DFFX1 \mat_r_reg[1][1][5]  ( .D(n136), .CLK(clk), .Q(\mat_r[1][1][5] ) );
  DFFX1 \mat_r_reg[1][1][4]  ( .D(n135), .CLK(clk), .Q(\mat_r[1][1][4] ) );
  DFFX1 \mat_r_reg[1][1][3]  ( .D(n134), .CLK(clk), .Q(\mat_r[1][1][3] ) );
  DFFX1 \mat_r_reg[1][1][2]  ( .D(n133), .CLK(clk), .Q(\mat_r[1][1][2] ) );
  DFFX1 \mat_r_reg[1][1][1]  ( .D(n132), .CLK(clk), .Q(\mat_r[1][1][1] ) );
  DFFX1 \mat_r_reg[1][1][0]  ( .D(n131), .CLK(clk), .Q(\mat_r[1][1][0] ) );
  DFFX1 \mat_r_reg[1][2][11]  ( .D(n130), .CLK(clk), .Q(\mat_r[1][2][11] ) );
  DFFX1 \mat_r_reg[1][2][10]  ( .D(n129), .CLK(clk), .Q(\mat_r[1][2][10] ) );
  DFFX1 \mat_r_reg[1][2][9]  ( .D(n128), .CLK(clk), .Q(\mat_r[1][2][9] ) );
  DFFX1 \mat_r_reg[1][2][8]  ( .D(n127), .CLK(clk), .Q(\mat_r[1][2][8] ) );
  DFFX1 \mat_r_reg[1][2][7]  ( .D(n126), .CLK(clk), .Q(\mat_r[1][2][7] ) );
  DFFX1 \mat_r_reg[1][2][6]  ( .D(n125), .CLK(clk), .Q(\mat_r[1][2][6] ) );
  DFFX1 \mat_r_reg[1][2][5]  ( .D(n124), .CLK(clk), .Q(\mat_r[1][2][5] ) );
  DFFX1 \mat_r_reg[1][2][4]  ( .D(n123), .CLK(clk), .Q(\mat_r[1][2][4] ) );
  DFFX1 \mat_r_reg[1][2][3]  ( .D(n122), .CLK(clk), .Q(\mat_r[1][2][3] ) );
  DFFX1 \mat_r_reg[1][2][2]  ( .D(n121), .CLK(clk), .Q(\mat_r[1][2][2] ) );
  DFFX1 \mat_r_reg[1][2][1]  ( .D(n120), .CLK(clk), .Q(\mat_r[1][2][1] ) );
  DFFX1 \mat_r_reg[1][2][0]  ( .D(n119), .CLK(clk), .Q(\mat_r[1][2][0] ) );
  DFFX1 \mat_r_reg[1][3][11]  ( .D(n118), .CLK(clk), .Q(\mat_r[1][3][11] ) );
  DFFX1 \mat_r_reg[1][3][10]  ( .D(n117), .CLK(clk), .Q(\mat_r[1][3][10] ) );
  DFFX1 \mat_r_reg[1][3][9]  ( .D(n116), .CLK(clk), .Q(\mat_r[1][3][9] ) );
  DFFX1 \mat_r_reg[1][3][8]  ( .D(n115), .CLK(clk), .Q(\mat_r[1][3][8] ) );
  DFFX1 \mat_r_reg[1][3][7]  ( .D(n114), .CLK(clk), .Q(\mat_r[1][3][7] ) );
  DFFX1 \mat_r_reg[1][3][6]  ( .D(n113), .CLK(clk), .Q(\mat_r[1][3][6] ) );
  DFFX1 \mat_r_reg[1][3][5]  ( .D(n112), .CLK(clk), .Q(\mat_r[1][3][5] ) );
  DFFX1 \mat_r_reg[1][3][4]  ( .D(n111), .CLK(clk), .Q(\mat_r[1][3][4] ) );
  DFFX1 \mat_r_reg[1][3][3]  ( .D(n110), .CLK(clk), .Q(\mat_r[1][3][3] ) );
  DFFX1 \mat_r_reg[1][3][2]  ( .D(n109), .CLK(clk), .Q(\mat_r[1][3][2] ) );
  DFFX1 \mat_r_reg[1][3][1]  ( .D(n108), .CLK(clk), .Q(\mat_r[1][3][1] ) );
  DFFX1 \mat_r_reg[1][3][0]  ( .D(n107), .CLK(clk), .Q(\mat_r[1][3][0] ) );
  DFFX1 \mat_r_reg[2][0][11]  ( .D(n106), .CLK(clk), .Q(\mat_r[2][0][11] ) );
  DFFX1 \mat_r_reg[2][0][10]  ( .D(n105), .CLK(clk), .Q(\mat_r[2][0][10] ) );
  DFFX1 \mat_r_reg[2][0][9]  ( .D(n104), .CLK(clk), .Q(\mat_r[2][0][9] ) );
  DFFX1 \mat_r_reg[2][0][8]  ( .D(n103), .CLK(clk), .Q(\mat_r[2][0][8] ) );
  DFFX1 \mat_r_reg[2][0][7]  ( .D(n102), .CLK(clk), .Q(\mat_r[2][0][7] ) );
  DFFX1 \mat_r_reg[2][0][6]  ( .D(n101), .CLK(clk), .Q(\mat_r[2][0][6] ) );
  DFFX1 \mat_r_reg[2][0][5]  ( .D(n100), .CLK(clk), .Q(\mat_r[2][0][5] ) );
  DFFX1 \mat_r_reg[2][0][4]  ( .D(n99), .CLK(clk), .Q(\mat_r[2][0][4] ) );
  DFFX1 \mat_r_reg[2][0][3]  ( .D(n98), .CLK(clk), .Q(\mat_r[2][0][3] ) );
  DFFX1 \mat_r_reg[2][0][2]  ( .D(n97), .CLK(clk), .Q(\mat_r[2][0][2] ) );
  DFFX1 \mat_r_reg[2][0][1]  ( .D(n96), .CLK(clk), .Q(\mat_r[2][0][1] ) );
  DFFX1 \mat_r_reg[2][0][0]  ( .D(n95), .CLK(clk), .Q(\mat_r[2][0][0] ) );
  DFFX1 \mat_r_reg[2][1][11]  ( .D(n94), .CLK(clk), .Q(\mat_r[2][1][11] ) );
  DFFX1 \mat_r_reg[2][1][10]  ( .D(n93), .CLK(clk), .Q(\mat_r[2][1][10] ) );
  DFFX1 \mat_r_reg[2][1][9]  ( .D(n92), .CLK(clk), .Q(\mat_r[2][1][9] ) );
  DFFX1 \mat_r_reg[2][1][8]  ( .D(n91), .CLK(clk), .Q(\mat_r[2][1][8] ) );
  DFFX1 \mat_r_reg[2][1][7]  ( .D(n90), .CLK(clk), .Q(\mat_r[2][1][7] ) );
  DFFX1 \mat_r_reg[2][1][6]  ( .D(n89), .CLK(clk), .Q(\mat_r[2][1][6] ) );
  DFFX1 \mat_r_reg[2][1][5]  ( .D(n88), .CLK(clk), .Q(\mat_r[2][1][5] ) );
  DFFX1 \mat_r_reg[2][1][4]  ( .D(n87), .CLK(clk), .Q(\mat_r[2][1][4] ) );
  DFFX1 \mat_r_reg[2][1][3]  ( .D(n86), .CLK(clk), .Q(\mat_r[2][1][3] ) );
  DFFX1 \mat_r_reg[2][1][2]  ( .D(n85), .CLK(clk), .Q(\mat_r[2][1][2] ) );
  DFFX1 \mat_r_reg[2][1][1]  ( .D(n84), .CLK(clk), .Q(\mat_r[2][1][1] ) );
  DFFX1 \mat_r_reg[2][1][0]  ( .D(n83), .CLK(clk), .Q(\mat_r[2][1][0] ) );
  DFFX1 \mat_r_reg[2][2][11]  ( .D(n82), .CLK(clk), .Q(\mat_r[2][2][11] ) );
  DFFX1 \mat_r_reg[2][2][10]  ( .D(n81), .CLK(clk), .Q(\mat_r[2][2][10] ) );
  DFFX1 \mat_r_reg[2][2][9]  ( .D(n80), .CLK(clk), .Q(\mat_r[2][2][9] ) );
  DFFX1 \mat_r_reg[2][2][8]  ( .D(n79), .CLK(clk), .Q(\mat_r[2][2][8] ) );
  DFFX1 \mat_r_reg[2][2][7]  ( .D(n78), .CLK(clk), .Q(\mat_r[2][2][7] ) );
  DFFX1 \mat_r_reg[2][2][6]  ( .D(n77), .CLK(clk), .Q(\mat_r[2][2][6] ) );
  DFFX1 \mat_r_reg[2][2][5]  ( .D(n76), .CLK(clk), .Q(\mat_r[2][2][5] ) );
  DFFX1 \mat_r_reg[2][2][4]  ( .D(n75), .CLK(clk), .Q(\mat_r[2][2][4] ) );
  DFFX1 \mat_r_reg[2][2][3]  ( .D(n74), .CLK(clk), .Q(\mat_r[2][2][3] ) );
  DFFX1 \mat_r_reg[2][2][2]  ( .D(n73), .CLK(clk), .Q(\mat_r[2][2][2] ) );
  DFFX1 \mat_r_reg[2][2][1]  ( .D(n72), .CLK(clk), .Q(\mat_r[2][2][1] ) );
  DFFX1 \mat_r_reg[2][2][0]  ( .D(n71), .CLK(clk), .Q(\mat_r[2][2][0] ) );
  DFFX1 \mat_r_reg[2][3][11]  ( .D(n70), .CLK(clk), .Q(\mat_r[2][3][11] ) );
  DFFX1 \mat_r_reg[2][3][10]  ( .D(n69), .CLK(clk), .Q(\mat_r[2][3][10] ) );
  DFFX1 \mat_r_reg[2][3][9]  ( .D(n68), .CLK(clk), .Q(\mat_r[2][3][9] ) );
  DFFX1 \mat_r_reg[2][3][8]  ( .D(n67), .CLK(clk), .Q(\mat_r[2][3][8] ) );
  DFFX1 \mat_r_reg[2][3][7]  ( .D(n66), .CLK(clk), .Q(\mat_r[2][3][7] ) );
  DFFX1 \mat_r_reg[2][3][6]  ( .D(n65), .CLK(clk), .Q(\mat_r[2][3][6] ) );
  DFFX1 \mat_r_reg[2][3][5]  ( .D(n64), .CLK(clk), .Q(\mat_r[2][3][5] ) );
  DFFX1 \mat_r_reg[2][3][4]  ( .D(n63), .CLK(clk), .Q(\mat_r[2][3][4] ) );
  DFFX1 \mat_r_reg[2][3][3]  ( .D(n62), .CLK(clk), .Q(\mat_r[2][3][3] ) );
  DFFX1 \mat_r_reg[2][3][2]  ( .D(n61), .CLK(clk), .Q(\mat_r[2][3][2] ) );
  DFFX1 \mat_r_reg[2][3][1]  ( .D(n60), .CLK(clk), .Q(\mat_r[2][3][1] ) );
  DFFX1 \mat_r_reg[2][3][0]  ( .D(n59), .CLK(clk), .Q(\mat_r[2][3][0] ) );
  DFFX1 \mat_r_reg[3][0][11]  ( .D(n58), .CLK(clk), .Q(\mat_r[3][0][11] ) );
  DFFX1 \mat_r_reg[3][0][10]  ( .D(n57), .CLK(clk), .Q(\mat_r[3][0][10] ) );
  DFFX1 \mat_r_reg[3][0][9]  ( .D(n56), .CLK(clk), .Q(\mat_r[3][0][9] ) );
  DFFX1 \mat_r_reg[3][0][8]  ( .D(n55), .CLK(clk), .Q(\mat_r[3][0][8] ) );
  DFFX1 \mat_r_reg[3][0][7]  ( .D(n54), .CLK(clk), .Q(\mat_r[3][0][7] ) );
  DFFX1 \mat_r_reg[3][0][6]  ( .D(n53), .CLK(clk), .Q(\mat_r[3][0][6] ) );
  DFFX1 \mat_r_reg[3][0][5]  ( .D(n52), .CLK(clk), .Q(\mat_r[3][0][5] ) );
  DFFX1 \mat_r_reg[3][0][4]  ( .D(n51), .CLK(clk), .Q(\mat_r[3][0][4] ) );
  DFFX1 \mat_r_reg[3][0][3]  ( .D(n50), .CLK(clk), .Q(\mat_r[3][0][3] ) );
  DFFX1 \mat_r_reg[3][0][2]  ( .D(n49), .CLK(clk), .Q(\mat_r[3][0][2] ) );
  DFFX1 \mat_r_reg[3][0][1]  ( .D(n48), .CLK(clk), .Q(\mat_r[3][0][1] ) );
  DFFX1 \mat_r_reg[3][0][0]  ( .D(n47), .CLK(clk), .Q(\mat_r[3][0][0] ) );
  DFFX1 \mat_r_reg[3][1][11]  ( .D(n46), .CLK(clk), .Q(\mat_r[3][1][11] ) );
  DFFX1 \mat_r_reg[3][1][10]  ( .D(n45), .CLK(clk), .Q(\mat_r[3][1][10] ) );
  DFFX1 \mat_r_reg[3][1][9]  ( .D(n44), .CLK(clk), .Q(\mat_r[3][1][9] ) );
  DFFX1 \mat_r_reg[3][1][8]  ( .D(n43), .CLK(clk), .Q(\mat_r[3][1][8] ) );
  DFFX1 \mat_r_reg[3][1][7]  ( .D(n42), .CLK(clk), .Q(\mat_r[3][1][7] ) );
  DFFX1 \mat_r_reg[3][1][6]  ( .D(n41), .CLK(clk), .Q(\mat_r[3][1][6] ) );
  DFFX1 \mat_r_reg[3][1][5]  ( .D(n40), .CLK(clk), .Q(\mat_r[3][1][5] ) );
  DFFX1 \mat_r_reg[3][1][4]  ( .D(n39), .CLK(clk), .Q(\mat_r[3][1][4] ) );
  DFFX1 \mat_r_reg[3][1][3]  ( .D(n38), .CLK(clk), .Q(\mat_r[3][1][3] ) );
  DFFX1 \mat_r_reg[3][1][2]  ( .D(n37), .CLK(clk), .Q(\mat_r[3][1][2] ) );
  DFFX1 \mat_r_reg[3][1][1]  ( .D(n36), .CLK(clk), .Q(\mat_r[3][1][1] ) );
  DFFX1 \mat_r_reg[3][1][0]  ( .D(n35), .CLK(clk), .Q(\mat_r[3][1][0] ) );
  DFFX1 \mat_r_reg[3][2][11]  ( .D(n34), .CLK(clk), .Q(\mat_r[3][2][11] ) );
  DFFX1 \mat_r_reg[3][2][10]  ( .D(n33), .CLK(clk), .Q(\mat_r[3][2][10] ) );
  DFFX1 \mat_r_reg[3][2][9]  ( .D(n32), .CLK(clk), .Q(\mat_r[3][2][9] ) );
  DFFX1 \mat_r_reg[3][2][8]  ( .D(n31), .CLK(clk), .Q(\mat_r[3][2][8] ) );
  DFFX1 \mat_r_reg[3][2][7]  ( .D(n30), .CLK(clk), .Q(\mat_r[3][2][7] ) );
  DFFX1 \mat_r_reg[3][2][6]  ( .D(n29), .CLK(clk), .Q(\mat_r[3][2][6] ) );
  DFFX1 \mat_r_reg[3][2][5]  ( .D(n28), .CLK(clk), .Q(\mat_r[3][2][5] ) );
  DFFX1 \mat_r_reg[3][2][4]  ( .D(n27), .CLK(clk), .Q(\mat_r[3][2][4] ) );
  DFFX1 \mat_r_reg[3][2][3]  ( .D(n26), .CLK(clk), .Q(\mat_r[3][2][3] ) );
  DFFX1 \mat_r_reg[3][2][2]  ( .D(n25), .CLK(clk), .Q(\mat_r[3][2][2] ) );
  DFFX1 \mat_r_reg[3][2][1]  ( .D(n24), .CLK(clk), .Q(\mat_r[3][2][1] ) );
  DFFX1 \mat_r_reg[3][2][0]  ( .D(n23), .CLK(clk), .Q(\mat_r[3][2][0] ) );
  DFFX1 \mat_r_reg[3][3][11]  ( .D(n22), .CLK(clk), .Q(\mat_r[3][3][11] ) );
  DFFX1 \mat_r_reg[3][3][10]  ( .D(n21), .CLK(clk), .Q(\mat_r[3][3][10] ) );
  DFFX1 \mat_r_reg[3][3][9]  ( .D(n20), .CLK(clk), .Q(\mat_r[3][3][9] ) );
  DFFX1 \mat_r_reg[3][3][8]  ( .D(n19), .CLK(clk), .Q(\mat_r[3][3][8] ) );
  DFFX1 \mat_r_reg[3][3][7]  ( .D(n18), .CLK(clk), .Q(\mat_r[3][3][7] ) );
  DFFX1 \mat_r_reg[3][3][6]  ( .D(n17), .CLK(clk), .Q(\mat_r[3][3][6] ) );
  DFFX1 \mat_r_reg[3][3][5]  ( .D(n16), .CLK(clk), .Q(\mat_r[3][3][5] ) );
  DFFX1 \mat_r_reg[3][3][4]  ( .D(n15), .CLK(clk), .Q(\mat_r[3][3][4] ) );
  DFFX1 \mat_r_reg[3][3][3]  ( .D(n14), .CLK(clk), .Q(\mat_r[3][3][3] ) );
  DFFX1 \mat_r_reg[3][3][2]  ( .D(n13), .CLK(clk), .Q(\mat_r[3][3][2] ) );
  DFFX1 \mat_r_reg[3][3][1]  ( .D(n12), .CLK(clk), .Q(\mat_r[3][3][1] ) );
  DFFX1 \mat_r_reg[3][3][0]  ( .D(n11), .CLK(clk), .Q(\mat_r[3][3][0] ) );
  NBUFFX2 U2 ( .INP(n1), .Z(n449) );
  NBUFFX2 U3 ( .INP(n1), .Z(n450) );
  NBUFFX2 U4 ( .INP(n1), .Z(n451) );
  NBUFFX2 U5 ( .INP(n1), .Z(n452) );
  NBUFFX2 U6 ( .INP(n1), .Z(n445) );
  NBUFFX2 U7 ( .INP(n1), .Z(n446) );
  NBUFFX2 U8 ( .INP(n1), .Z(n447) );
  NBUFFX2 U9 ( .INP(n1), .Z(n448) );
  NBUFFX2 U10 ( .INP(n2), .Z(n441) );
  NBUFFX2 U11 ( .INP(n2), .Z(n442) );
  NBUFFX2 U12 ( .INP(n2), .Z(n443) );
  NBUFFX2 U13 ( .INP(n2), .Z(n444) );
  NBUFFX2 U14 ( .INP(n3), .Z(n433) );
  NBUFFX2 U15 ( .INP(n3), .Z(n434) );
  NBUFFX2 U16 ( .INP(n3), .Z(n435) );
  NBUFFX2 U17 ( .INP(n3), .Z(n436) );
  NBUFFX2 U18 ( .INP(n2), .Z(n437) );
  NBUFFX2 U19 ( .INP(n2), .Z(n438) );
  NBUFFX2 U20 ( .INP(n2), .Z(n439) );
  NBUFFX2 U21 ( .INP(n2), .Z(n440) );
  NBUFFX2 U22 ( .INP(n3), .Z(n429) );
  NBUFFX2 U23 ( .INP(n3), .Z(n430) );
  NBUFFX2 U24 ( .INP(n3), .Z(n431) );
  NBUFFX2 U25 ( .INP(n3), .Z(n432) );
  NBUFFX2 U26 ( .INP(n4), .Z(n457) );
  NBUFFX2 U27 ( .INP(n4), .Z(n458) );
  NBUFFX2 U28 ( .INP(n4), .Z(n459) );
  NBUFFX2 U29 ( .INP(n4), .Z(n460) );
  NBUFFX2 U30 ( .INP(n4), .Z(n453) );
  NBUFFX2 U31 ( .INP(n4), .Z(n454) );
  NBUFFX2 U32 ( .INP(n4), .Z(n455) );
  NBUFFX2 U33 ( .INP(n4), .Z(n456) );
  AND3X1 U34 ( .IN1(wr_enable), .IN2(w_col_sel[1]), .IN3(n462), .Q(n1) );
  AND3X1 U35 ( .IN1(wr_enable), .IN2(w_col_sel[0]), .IN3(n461), .Q(n2) );
  AND3X1 U36 ( .IN1(wr_enable), .IN2(n462), .IN3(n461), .Q(n3) );
  AND3X1 U37 ( .IN1(w_col_sel[1]), .IN2(w_col_sel[0]), .IN3(wr_enable), .Q(n4)
         );
  INVX0 U38 ( .INP(w_col_sel[1]), .ZN(n461) );
  INVX0 U39 ( .INP(w_col_sel[0]), .ZN(n462) );
  NBUFFX4 U40 ( .INP(N6), .Z(n398) );
  NBUFFX4 U41 ( .INP(N6), .Z(n402) );
  NBUFFX4 U42 ( .INP(N6), .Z(n397) );
  NBUFFX4 U43 ( .INP(N6), .Z(n401) );
  NBUFFX4 U44 ( .INP(N6), .Z(n400) );
  NBUFFX4 U45 ( .INP(N6), .Z(n404) );
  NBUFFX4 U46 ( .INP(N6), .Z(n399) );
  NBUFFX4 U47 ( .INP(N6), .Z(n403) );
  NBUFFX4 U48 ( .INP(N10), .Z(n423) );
  NBUFFX4 U49 ( .INP(N10), .Z(n424) );
  NBUFFX4 U50 ( .INP(N12), .Z(n428) );
  NBUFFX4 U51 ( .INP(N12), .Z(n427) );
  NBUFFX2 U52 ( .INP(N11), .Z(n421) );
  NBUFFX2 U53 ( .INP(N11), .Z(n422) );
  NBUFFX2 U54 ( .INP(N13), .Z(n426) );
  NBUFFX2 U55 ( .INP(N13), .Z(n425) );
  MUX41X1 U56 ( .IN1(\mat_i[0][3][0] ), .IN3(\mat_i[2][3][0] ), .IN2(
        \mat_i[1][3][0] ), .IN4(\mat_i[3][3][0] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][0] ) );
  MUX41X1 U57 ( .IN1(\mat_i[0][3][1] ), .IN3(\mat_i[2][3][1] ), .IN2(
        \mat_i[1][3][1] ), .IN4(\mat_i[3][3][1] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][1] ) );
  MUX41X1 U58 ( .IN1(\mat_i[0][3][2] ), .IN3(\mat_i[2][3][2] ), .IN2(
        \mat_i[1][3][2] ), .IN4(\mat_i[3][3][2] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][2] ) );
  MUX41X1 U59 ( .IN1(\mat_i[0][3][3] ), .IN3(\mat_i[2][3][3] ), .IN2(
        \mat_i[1][3][3] ), .IN4(\mat_i[3][3][3] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][3] ) );
  MUX41X1 U60 ( .IN1(\mat_i[0][3][4] ), .IN3(\mat_i[2][3][4] ), .IN2(
        \mat_i[1][3][4] ), .IN4(\mat_i[3][3][4] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][4] ) );
  MUX41X1 U61 ( .IN1(\mat_i[0][3][5] ), .IN3(\mat_i[2][3][5] ), .IN2(
        \mat_i[1][3][5] ), .IN4(\mat_i[3][3][5] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][5] ) );
  MUX41X1 U62 ( .IN1(\mat_i[0][3][6] ), .IN3(\mat_i[2][3][6] ), .IN2(
        \mat_i[1][3][6] ), .IN4(\mat_i[3][3][6] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][6] ) );
  MUX41X1 U63 ( .IN1(\mat_i[0][3][7] ), .IN3(\mat_i[2][3][7] ), .IN2(
        \mat_i[1][3][7] ), .IN4(\mat_i[3][3][7] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][7] ) );
  MUX41X1 U64 ( .IN1(\mat_i[0][3][8] ), .IN3(\mat_i[2][3][8] ), .IN2(
        \mat_i[1][3][8] ), .IN4(\mat_i[3][3][8] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][8] ) );
  MUX41X1 U65 ( .IN1(\mat_i[0][3][9] ), .IN3(\mat_i[2][3][9] ), .IN2(
        \mat_i[1][3][9] ), .IN4(\mat_i[3][3][9] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][9] ) );
  MUX41X1 U66 ( .IN1(\mat_i[0][3][10] ), .IN3(\mat_i[2][3][10] ), .IN2(
        \mat_i[1][3][10] ), .IN4(\mat_i[3][3][10] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][10] ) );
  MUX41X1 U67 ( .IN1(\mat_i[0][3][11] ), .IN3(\mat_i[2][3][11] ), .IN2(
        \mat_i[1][3][11] ), .IN4(\mat_i[3][3][11] ), .S0(n5), .S1(n397), .Q(
        \vector_out_i[3][11] ) );
  MUX41X1 U68 ( .IN1(\mat_i[0][2][0] ), .IN3(\mat_i[2][2][0] ), .IN2(
        \mat_i[1][2][0] ), .IN4(\mat_i[3][2][0] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][0] ) );
  MUX41X1 U69 ( .IN1(\mat_i[0][2][1] ), .IN3(\mat_i[2][2][1] ), .IN2(
        \mat_i[1][2][1] ), .IN4(\mat_i[3][2][1] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][1] ) );
  MUX41X1 U70 ( .IN1(\mat_i[0][2][2] ), .IN3(\mat_i[2][2][2] ), .IN2(
        \mat_i[1][2][2] ), .IN4(\mat_i[3][2][2] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][2] ) );
  MUX41X1 U71 ( .IN1(\mat_i[0][2][3] ), .IN3(\mat_i[2][2][3] ), .IN2(
        \mat_i[1][2][3] ), .IN4(\mat_i[3][2][3] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][3] ) );
  MUX41X1 U72 ( .IN1(\mat_i[0][2][4] ), .IN3(\mat_i[2][2][4] ), .IN2(
        \mat_i[1][2][4] ), .IN4(\mat_i[3][2][4] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][4] ) );
  MUX41X1 U73 ( .IN1(\mat_i[0][2][5] ), .IN3(\mat_i[2][2][5] ), .IN2(
        \mat_i[1][2][5] ), .IN4(\mat_i[3][2][5] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][5] ) );
  MUX41X1 U74 ( .IN1(\mat_i[0][2][6] ), .IN3(\mat_i[2][2][6] ), .IN2(
        \mat_i[1][2][6] ), .IN4(\mat_i[3][2][6] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][6] ) );
  MUX41X1 U75 ( .IN1(\mat_i[0][2][7] ), .IN3(\mat_i[2][2][7] ), .IN2(
        \mat_i[1][2][7] ), .IN4(\mat_i[3][2][7] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][7] ) );
  MUX41X1 U76 ( .IN1(\mat_i[0][2][8] ), .IN3(\mat_i[2][2][8] ), .IN2(
        \mat_i[1][2][8] ), .IN4(\mat_i[3][2][8] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][8] ) );
  MUX41X1 U77 ( .IN1(\mat_i[0][2][9] ), .IN3(\mat_i[2][2][9] ), .IN2(
        \mat_i[1][2][9] ), .IN4(\mat_i[3][2][9] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][9] ) );
  MUX41X1 U78 ( .IN1(\mat_i[0][2][10] ), .IN3(\mat_i[2][2][10] ), .IN2(
        \mat_i[1][2][10] ), .IN4(\mat_i[3][2][10] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][10] ) );
  MUX41X1 U79 ( .IN1(\mat_i[0][2][11] ), .IN3(\mat_i[2][2][11] ), .IN2(
        \mat_i[1][2][11] ), .IN4(\mat_i[3][2][11] ), .S0(n6), .S1(n398), .Q(
        \vector_out_i[2][11] ) );
  MUX41X1 U80 ( .IN1(\mat_i[0][1][0] ), .IN3(\mat_i[2][1][0] ), .IN2(
        \mat_i[1][1][0] ), .IN4(\mat_i[3][1][0] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][0] ) );
  MUX41X1 U81 ( .IN1(\mat_i[0][1][1] ), .IN3(\mat_i[2][1][1] ), .IN2(
        \mat_i[1][1][1] ), .IN4(\mat_i[3][1][1] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][1] ) );
  MUX41X1 U82 ( .IN1(\mat_i[0][1][2] ), .IN3(\mat_i[2][1][2] ), .IN2(
        \mat_i[1][1][2] ), .IN4(\mat_i[3][1][2] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][2] ) );
  MUX41X1 U83 ( .IN1(\mat_i[0][1][3] ), .IN3(\mat_i[2][1][3] ), .IN2(
        \mat_i[1][1][3] ), .IN4(\mat_i[3][1][3] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][3] ) );
  MUX41X1 U84 ( .IN1(\mat_i[0][1][4] ), .IN3(\mat_i[2][1][4] ), .IN2(
        \mat_i[1][1][4] ), .IN4(\mat_i[3][1][4] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][4] ) );
  MUX41X1 U85 ( .IN1(\mat_i[0][1][5] ), .IN3(\mat_i[2][1][5] ), .IN2(
        \mat_i[1][1][5] ), .IN4(\mat_i[3][1][5] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][5] ) );
  MUX41X1 U86 ( .IN1(\mat_i[0][1][6] ), .IN3(\mat_i[2][1][6] ), .IN2(
        \mat_i[1][1][6] ), .IN4(\mat_i[3][1][6] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][6] ) );
  MUX41X1 U87 ( .IN1(\mat_i[0][1][7] ), .IN3(\mat_i[2][1][7] ), .IN2(
        \mat_i[1][1][7] ), .IN4(\mat_i[3][1][7] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][7] ) );
  MUX41X1 U88 ( .IN1(\mat_i[0][1][8] ), .IN3(\mat_i[2][1][8] ), .IN2(
        \mat_i[1][1][8] ), .IN4(\mat_i[3][1][8] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][8] ) );
  MUX41X1 U89 ( .IN1(\mat_i[0][1][9] ), .IN3(\mat_i[2][1][9] ), .IN2(
        \mat_i[1][1][9] ), .IN4(\mat_i[3][1][9] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][9] ) );
  MUX41X1 U90 ( .IN1(\mat_i[0][1][10] ), .IN3(\mat_i[2][1][10] ), .IN2(
        \mat_i[1][1][10] ), .IN4(\mat_i[3][1][10] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][10] ) );
  MUX41X1 U91 ( .IN1(\mat_i[0][1][11] ), .IN3(\mat_i[2][1][11] ), .IN2(
        \mat_i[1][1][11] ), .IN4(\mat_i[3][1][11] ), .S0(n7), .S1(n399), .Q(
        \vector_out_i[1][11] ) );
  MUX41X1 U92 ( .IN1(\mat_i[0][0][0] ), .IN3(\mat_i[2][0][0] ), .IN2(
        \mat_i[1][0][0] ), .IN4(\mat_i[3][0][0] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][0] ) );
  MUX41X1 U93 ( .IN1(\mat_i[0][0][1] ), .IN3(\mat_i[2][0][1] ), .IN2(
        \mat_i[1][0][1] ), .IN4(\mat_i[3][0][1] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][1] ) );
  MUX41X1 U94 ( .IN1(\mat_i[0][0][2] ), .IN3(\mat_i[2][0][2] ), .IN2(
        \mat_i[1][0][2] ), .IN4(\mat_i[3][0][2] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][2] ) );
  MUX41X1 U95 ( .IN1(\mat_i[0][0][3] ), .IN3(\mat_i[2][0][3] ), .IN2(
        \mat_i[1][0][3] ), .IN4(\mat_i[3][0][3] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][3] ) );
  MUX41X1 U96 ( .IN1(\mat_i[0][0][4] ), .IN3(\mat_i[2][0][4] ), .IN2(
        \mat_i[1][0][4] ), .IN4(\mat_i[3][0][4] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][4] ) );
  MUX41X1 U97 ( .IN1(\mat_i[0][0][5] ), .IN3(\mat_i[2][0][5] ), .IN2(
        \mat_i[1][0][5] ), .IN4(\mat_i[3][0][5] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][5] ) );
  MUX41X1 U98 ( .IN1(\mat_i[0][0][6] ), .IN3(\mat_i[2][0][6] ), .IN2(
        \mat_i[1][0][6] ), .IN4(\mat_i[3][0][6] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][6] ) );
  MUX41X1 U99 ( .IN1(\mat_i[0][0][7] ), .IN3(\mat_i[2][0][7] ), .IN2(
        \mat_i[1][0][7] ), .IN4(\mat_i[3][0][7] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][7] ) );
  MUX41X1 U100 ( .IN1(\mat_i[0][0][8] ), .IN3(\mat_i[2][0][8] ), .IN2(
        \mat_i[1][0][8] ), .IN4(\mat_i[3][0][8] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][8] ) );
  MUX41X1 U101 ( .IN1(\mat_i[0][0][9] ), .IN3(\mat_i[2][0][9] ), .IN2(
        \mat_i[1][0][9] ), .IN4(\mat_i[3][0][9] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][9] ) );
  MUX41X1 U102 ( .IN1(\mat_i[0][0][10] ), .IN3(\mat_i[2][0][10] ), .IN2(
        \mat_i[1][0][10] ), .IN4(\mat_i[3][0][10] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][10] ) );
  MUX41X1 U103 ( .IN1(\mat_i[0][0][11] ), .IN3(\mat_i[2][0][11] ), .IN2(
        \mat_i[1][0][11] ), .IN4(\mat_i[3][0][11] ), .S0(n8), .S1(n400), .Q(
        \vector_out_i[0][11] ) );
  MUX41X1 U104 ( .IN1(\mat_r[0][3][0] ), .IN3(\mat_r[2][3][0] ), .IN2(
        \mat_r[1][3][0] ), .IN4(\mat_r[3][3][0] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][0] ) );
  MUX41X1 U105 ( .IN1(\mat_r[0][3][1] ), .IN3(\mat_r[2][3][1] ), .IN2(
        \mat_r[1][3][1] ), .IN4(\mat_r[3][3][1] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][1] ) );
  MUX41X1 U106 ( .IN1(\mat_r[0][3][2] ), .IN3(\mat_r[2][3][2] ), .IN2(
        \mat_r[1][3][2] ), .IN4(\mat_r[3][3][2] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][2] ) );
  MUX41X1 U107 ( .IN1(\mat_r[0][3][3] ), .IN3(\mat_r[2][3][3] ), .IN2(
        \mat_r[1][3][3] ), .IN4(\mat_r[3][3][3] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][3] ) );
  MUX41X1 U108 ( .IN1(\mat_r[0][3][4] ), .IN3(\mat_r[2][3][4] ), .IN2(
        \mat_r[1][3][4] ), .IN4(\mat_r[3][3][4] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][4] ) );
  MUX41X1 U109 ( .IN1(\mat_r[0][3][5] ), .IN3(\mat_r[2][3][5] ), .IN2(
        \mat_r[1][3][5] ), .IN4(\mat_r[3][3][5] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][5] ) );
  MUX41X1 U110 ( .IN1(\mat_r[0][3][6] ), .IN3(\mat_r[2][3][6] ), .IN2(
        \mat_r[1][3][6] ), .IN4(\mat_r[3][3][6] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][6] ) );
  MUX41X1 U111 ( .IN1(\mat_r[0][3][7] ), .IN3(\mat_r[2][3][7] ), .IN2(
        \mat_r[1][3][7] ), .IN4(\mat_r[3][3][7] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][7] ) );
  MUX41X1 U112 ( .IN1(\mat_r[0][3][8] ), .IN3(\mat_r[2][3][8] ), .IN2(
        \mat_r[1][3][8] ), .IN4(\mat_r[3][3][8] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][8] ) );
  MUX41X1 U113 ( .IN1(\mat_r[0][3][9] ), .IN3(\mat_r[2][3][9] ), .IN2(
        \mat_r[1][3][9] ), .IN4(\mat_r[3][3][9] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][9] ) );
  MUX41X1 U114 ( .IN1(\mat_r[0][3][10] ), .IN3(\mat_r[2][3][10] ), .IN2(
        \mat_r[1][3][10] ), .IN4(\mat_r[3][3][10] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][10] ) );
  MUX41X1 U115 ( .IN1(\mat_r[0][3][11] ), .IN3(\mat_r[2][3][11] ), .IN2(
        \mat_r[1][3][11] ), .IN4(\mat_r[3][3][11] ), .S0(n9), .S1(n401), .Q(
        \vector_out_r[3][11] ) );
  MUX41X1 U116 ( .IN1(\mat_r[0][2][0] ), .IN3(\mat_r[2][2][0] ), .IN2(
        \mat_r[1][2][0] ), .IN4(\mat_r[3][2][0] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][0] ) );
  MUX41X1 U117 ( .IN1(\mat_r[0][2][1] ), .IN3(\mat_r[2][2][1] ), .IN2(
        \mat_r[1][2][1] ), .IN4(\mat_r[3][2][1] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][1] ) );
  MUX41X1 U118 ( .IN1(\mat_r[0][2][2] ), .IN3(\mat_r[2][2][2] ), .IN2(
        \mat_r[1][2][2] ), .IN4(\mat_r[3][2][2] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][2] ) );
  MUX41X1 U119 ( .IN1(\mat_r[0][2][3] ), .IN3(\mat_r[2][2][3] ), .IN2(
        \mat_r[1][2][3] ), .IN4(\mat_r[3][2][3] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][3] ) );
  MUX41X1 U120 ( .IN1(\mat_r[0][2][4] ), .IN3(\mat_r[2][2][4] ), .IN2(
        \mat_r[1][2][4] ), .IN4(\mat_r[3][2][4] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][4] ) );
  MUX41X1 U121 ( .IN1(\mat_r[0][2][5] ), .IN3(\mat_r[2][2][5] ), .IN2(
        \mat_r[1][2][5] ), .IN4(\mat_r[3][2][5] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][5] ) );
  MUX41X1 U122 ( .IN1(\mat_r[0][2][6] ), .IN3(\mat_r[2][2][6] ), .IN2(
        \mat_r[1][2][6] ), .IN4(\mat_r[3][2][6] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][6] ) );
  MUX41X1 U123 ( .IN1(\mat_r[0][2][7] ), .IN3(\mat_r[2][2][7] ), .IN2(
        \mat_r[1][2][7] ), .IN4(\mat_r[3][2][7] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][7] ) );
  MUX41X1 U124 ( .IN1(\mat_r[0][2][8] ), .IN3(\mat_r[2][2][8] ), .IN2(
        \mat_r[1][2][8] ), .IN4(\mat_r[3][2][8] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][8] ) );
  MUX41X1 U125 ( .IN1(\mat_r[0][2][9] ), .IN3(\mat_r[2][2][9] ), .IN2(
        \mat_r[1][2][9] ), .IN4(\mat_r[3][2][9] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][9] ) );
  MUX41X1 U126 ( .IN1(\mat_r[0][2][10] ), .IN3(\mat_r[2][2][10] ), .IN2(
        \mat_r[1][2][10] ), .IN4(\mat_r[3][2][10] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][10] ) );
  MUX41X1 U127 ( .IN1(\mat_r[0][2][11] ), .IN3(\mat_r[2][2][11] ), .IN2(
        \mat_r[1][2][11] ), .IN4(\mat_r[3][2][11] ), .S0(n10), .S1(n402), .Q(
        \vector_out_r[2][11] ) );
  MUX41X1 U128 ( .IN1(\mat_r[0][1][0] ), .IN3(\mat_r[2][1][0] ), .IN2(
        \mat_r[1][1][0] ), .IN4(\mat_r[3][1][0] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][0] ) );
  MUX41X1 U129 ( .IN1(\mat_r[0][1][1] ), .IN3(\mat_r[2][1][1] ), .IN2(
        \mat_r[1][1][1] ), .IN4(\mat_r[3][1][1] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][1] ) );
  MUX41X1 U130 ( .IN1(\mat_r[0][1][2] ), .IN3(\mat_r[2][1][2] ), .IN2(
        \mat_r[1][1][2] ), .IN4(\mat_r[3][1][2] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][2] ) );
  MUX41X1 U131 ( .IN1(\mat_r[0][1][3] ), .IN3(\mat_r[2][1][3] ), .IN2(
        \mat_r[1][1][3] ), .IN4(\mat_r[3][1][3] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][3] ) );
  MUX41X1 U132 ( .IN1(\mat_r[0][1][4] ), .IN3(\mat_r[2][1][4] ), .IN2(
        \mat_r[1][1][4] ), .IN4(\mat_r[3][1][4] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][4] ) );
  MUX41X1 U133 ( .IN1(\mat_r[0][1][5] ), .IN3(\mat_r[2][1][5] ), .IN2(
        \mat_r[1][1][5] ), .IN4(\mat_r[3][1][5] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][5] ) );
  MUX41X1 U134 ( .IN1(\mat_r[0][1][6] ), .IN3(\mat_r[2][1][6] ), .IN2(
        \mat_r[1][1][6] ), .IN4(\mat_r[3][1][6] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][6] ) );
  MUX41X1 U135 ( .IN1(\mat_r[0][1][7] ), .IN3(\mat_r[2][1][7] ), .IN2(
        \mat_r[1][1][7] ), .IN4(\mat_r[3][1][7] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][7] ) );
  MUX41X1 U136 ( .IN1(\mat_r[0][1][8] ), .IN3(\mat_r[2][1][8] ), .IN2(
        \mat_r[1][1][8] ), .IN4(\mat_r[3][1][8] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][8] ) );
  MUX41X1 U137 ( .IN1(\mat_r[0][1][9] ), .IN3(\mat_r[2][1][9] ), .IN2(
        \mat_r[1][1][9] ), .IN4(\mat_r[3][1][9] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][9] ) );
  MUX41X1 U138 ( .IN1(\mat_r[0][1][10] ), .IN3(\mat_r[2][1][10] ), .IN2(
        \mat_r[1][1][10] ), .IN4(\mat_r[3][1][10] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][10] ) );
  MUX41X1 U139 ( .IN1(\mat_r[0][1][11] ), .IN3(\mat_r[2][1][11] ), .IN2(
        \mat_r[1][1][11] ), .IN4(\mat_r[3][1][11] ), .S0(n395), .S1(n403), .Q(
        \vector_out_r[1][11] ) );
  MUX41X1 U140 ( .IN1(\mat_r[0][0][0] ), .IN3(\mat_r[2][0][0] ), .IN2(
        \mat_r[1][0][0] ), .IN4(\mat_r[3][0][0] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][0] ) );
  MUX41X1 U141 ( .IN1(\mat_r[0][0][1] ), .IN3(\mat_r[2][0][1] ), .IN2(
        \mat_r[1][0][1] ), .IN4(\mat_r[3][0][1] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][1] ) );
  MUX41X1 U142 ( .IN1(\mat_r[0][0][2] ), .IN3(\mat_r[2][0][2] ), .IN2(
        \mat_r[1][0][2] ), .IN4(\mat_r[3][0][2] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][2] ) );
  MUX41X1 U143 ( .IN1(\mat_r[0][0][3] ), .IN3(\mat_r[2][0][3] ), .IN2(
        \mat_r[1][0][3] ), .IN4(\mat_r[3][0][3] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][3] ) );
  MUX41X1 U144 ( .IN1(\mat_r[0][0][4] ), .IN3(\mat_r[2][0][4] ), .IN2(
        \mat_r[1][0][4] ), .IN4(\mat_r[3][0][4] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][4] ) );
  MUX41X1 U145 ( .IN1(\mat_r[0][0][5] ), .IN3(\mat_r[2][0][5] ), .IN2(
        \mat_r[1][0][5] ), .IN4(\mat_r[3][0][5] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][5] ) );
  MUX41X1 U146 ( .IN1(\mat_r[0][0][6] ), .IN3(\mat_r[2][0][6] ), .IN2(
        \mat_r[1][0][6] ), .IN4(\mat_r[3][0][6] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][6] ) );
  MUX41X1 U147 ( .IN1(\mat_r[0][0][7] ), .IN3(\mat_r[2][0][7] ), .IN2(
        \mat_r[1][0][7] ), .IN4(\mat_r[3][0][7] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][7] ) );
  MUX41X1 U148 ( .IN1(\mat_r[0][0][8] ), .IN3(\mat_r[2][0][8] ), .IN2(
        \mat_r[1][0][8] ), .IN4(\mat_r[3][0][8] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][8] ) );
  MUX41X1 U149 ( .IN1(\mat_r[0][0][9] ), .IN3(\mat_r[2][0][9] ), .IN2(
        \mat_r[1][0][9] ), .IN4(\mat_r[3][0][9] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][9] ) );
  MUX41X1 U150 ( .IN1(\mat_r[0][0][10] ), .IN3(\mat_r[2][0][10] ), .IN2(
        \mat_r[1][0][10] ), .IN4(\mat_r[3][0][10] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][10] ) );
  MUX41X1 U151 ( .IN1(\mat_r[0][0][11] ), .IN3(\mat_r[2][0][11] ), .IN2(
        \mat_r[1][0][11] ), .IN4(\mat_r[3][0][11] ), .S0(n396), .S1(n404), .Q(
        \vector_out_r[0][11] ) );
  DELLN2X2 U152 ( .INP(N7), .Z(n5) );
  DELLN2X2 U153 ( .INP(N7), .Z(n6) );
  DELLN2X2 U154 ( .INP(N7), .Z(n7) );
  DELLN2X2 U155 ( .INP(N7), .Z(n8) );
  DELLN2X2 U156 ( .INP(N7), .Z(n9) );
  DELLN2X2 U157 ( .INP(N7), .Z(n10) );
  DELLN2X2 U158 ( .INP(N7), .Z(n395) );
  DELLN2X2 U159 ( .INP(N7), .Z(n396) );
  MUX41X1 U160 ( .IN1(\mat_i[0][3][0] ), .IN3(\mat_i[2][3][0] ), .IN2(
        \mat_i[1][3][0] ), .IN4(\mat_i[3][3][0] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][0] ) );
  MUX41X1 U161 ( .IN1(\mat_i[0][3][1] ), .IN3(\mat_i[2][3][1] ), .IN2(
        \mat_i[1][3][1] ), .IN4(\mat_i[3][3][1] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][1] ) );
  MUX41X1 U162 ( .IN1(\mat_i[0][3][2] ), .IN3(\mat_i[2][3][2] ), .IN2(
        \mat_i[1][3][2] ), .IN4(\mat_i[3][3][2] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][2] ) );
  MUX41X1 U163 ( .IN1(\mat_i[0][3][3] ), .IN3(\mat_i[2][3][3] ), .IN2(
        \mat_i[1][3][3] ), .IN4(\mat_i[3][3][3] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][3] ) );
  MUX41X1 U164 ( .IN1(\mat_i[0][3][4] ), .IN3(\mat_i[2][3][4] ), .IN2(
        \mat_i[1][3][4] ), .IN4(\mat_i[3][3][4] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][4] ) );
  MUX41X1 U165 ( .IN1(\mat_i[0][3][5] ), .IN3(\mat_i[2][3][5] ), .IN2(
        \mat_i[1][3][5] ), .IN4(\mat_i[3][3][5] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][5] ) );
  MUX41X1 U166 ( .IN1(\mat_i[0][3][6] ), .IN3(\mat_i[2][3][6] ), .IN2(
        \mat_i[1][3][6] ), .IN4(\mat_i[3][3][6] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][6] ) );
  MUX41X1 U167 ( .IN1(\mat_i[0][3][7] ), .IN3(\mat_i[2][3][7] ), .IN2(
        \mat_i[1][3][7] ), .IN4(\mat_i[3][3][7] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][7] ) );
  MUX41X1 U168 ( .IN1(\mat_i[0][3][8] ), .IN3(\mat_i[2][3][8] ), .IN2(
        \mat_i[1][3][8] ), .IN4(\mat_i[3][3][8] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][8] ) );
  MUX41X1 U169 ( .IN1(\mat_i[0][3][9] ), .IN3(\mat_i[2][3][9] ), .IN2(
        \mat_i[1][3][9] ), .IN4(\mat_i[3][3][9] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][9] ) );
  MUX41X1 U170 ( .IN1(\mat_i[0][3][10] ), .IN3(\mat_i[2][3][10] ), .IN2(
        \mat_i[1][3][10] ), .IN4(\mat_i[3][3][10] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][10] ) );
  MUX41X1 U171 ( .IN1(\mat_i[0][3][11] ), .IN3(\mat_i[2][3][11] ), .IN2(
        \mat_i[1][3][11] ), .IN4(\mat_i[3][3][11] ), .S0(n405), .S1(n413), .Q(
        \vector_out_i2[3][11] ) );
  MUX41X1 U172 ( .IN1(\mat_i[0][2][0] ), .IN3(\mat_i[2][2][0] ), .IN2(
        \mat_i[1][2][0] ), .IN4(\mat_i[3][2][0] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][0] ) );
  MUX41X1 U173 ( .IN1(\mat_i[0][2][1] ), .IN3(\mat_i[2][2][1] ), .IN2(
        \mat_i[1][2][1] ), .IN4(\mat_i[3][2][1] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][1] ) );
  MUX41X1 U174 ( .IN1(\mat_i[0][2][2] ), .IN3(\mat_i[2][2][2] ), .IN2(
        \mat_i[1][2][2] ), .IN4(\mat_i[3][2][2] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][2] ) );
  MUX41X1 U175 ( .IN1(\mat_i[0][2][3] ), .IN3(\mat_i[2][2][3] ), .IN2(
        \mat_i[1][2][3] ), .IN4(\mat_i[3][2][3] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][3] ) );
  MUX41X1 U176 ( .IN1(\mat_i[0][2][4] ), .IN3(\mat_i[2][2][4] ), .IN2(
        \mat_i[1][2][4] ), .IN4(\mat_i[3][2][4] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][4] ) );
  MUX41X1 U177 ( .IN1(\mat_i[0][2][5] ), .IN3(\mat_i[2][2][5] ), .IN2(
        \mat_i[1][2][5] ), .IN4(\mat_i[3][2][5] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][5] ) );
  MUX41X1 U178 ( .IN1(\mat_i[0][2][6] ), .IN3(\mat_i[2][2][6] ), .IN2(
        \mat_i[1][2][6] ), .IN4(\mat_i[3][2][6] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][6] ) );
  MUX41X1 U179 ( .IN1(\mat_i[0][2][7] ), .IN3(\mat_i[2][2][7] ), .IN2(
        \mat_i[1][2][7] ), .IN4(\mat_i[3][2][7] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][7] ) );
  MUX41X1 U180 ( .IN1(\mat_i[0][2][8] ), .IN3(\mat_i[2][2][8] ), .IN2(
        \mat_i[1][2][8] ), .IN4(\mat_i[3][2][8] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][8] ) );
  MUX41X1 U181 ( .IN1(\mat_i[0][2][9] ), .IN3(\mat_i[2][2][9] ), .IN2(
        \mat_i[1][2][9] ), .IN4(\mat_i[3][2][9] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][9] ) );
  MUX41X1 U182 ( .IN1(\mat_i[0][2][10] ), .IN3(\mat_i[2][2][10] ), .IN2(
        \mat_i[1][2][10] ), .IN4(\mat_i[3][2][10] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][10] ) );
  MUX41X1 U183 ( .IN1(\mat_i[0][2][11] ), .IN3(\mat_i[2][2][11] ), .IN2(
        \mat_i[1][2][11] ), .IN4(\mat_i[3][2][11] ), .S0(n406), .S1(n414), .Q(
        \vector_out_i2[2][11] ) );
  MUX41X1 U184 ( .IN1(\mat_i[0][1][0] ), .IN3(\mat_i[2][1][0] ), .IN2(
        \mat_i[1][1][0] ), .IN4(\mat_i[3][1][0] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][0] ) );
  MUX41X1 U185 ( .IN1(\mat_i[0][1][1] ), .IN3(\mat_i[2][1][1] ), .IN2(
        \mat_i[1][1][1] ), .IN4(\mat_i[3][1][1] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][1] ) );
  MUX41X1 U186 ( .IN1(\mat_i[0][1][2] ), .IN3(\mat_i[2][1][2] ), .IN2(
        \mat_i[1][1][2] ), .IN4(\mat_i[3][1][2] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][2] ) );
  MUX41X1 U187 ( .IN1(\mat_i[0][1][3] ), .IN3(\mat_i[2][1][3] ), .IN2(
        \mat_i[1][1][3] ), .IN4(\mat_i[3][1][3] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][3] ) );
  MUX41X1 U188 ( .IN1(\mat_i[0][1][4] ), .IN3(\mat_i[2][1][4] ), .IN2(
        \mat_i[1][1][4] ), .IN4(\mat_i[3][1][4] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][4] ) );
  MUX41X1 U189 ( .IN1(\mat_i[0][1][5] ), .IN3(\mat_i[2][1][5] ), .IN2(
        \mat_i[1][1][5] ), .IN4(\mat_i[3][1][5] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][5] ) );
  MUX41X1 U190 ( .IN1(\mat_i[0][1][6] ), .IN3(\mat_i[2][1][6] ), .IN2(
        \mat_i[1][1][6] ), .IN4(\mat_i[3][1][6] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][6] ) );
  MUX41X1 U191 ( .IN1(\mat_i[0][1][7] ), .IN3(\mat_i[2][1][7] ), .IN2(
        \mat_i[1][1][7] ), .IN4(\mat_i[3][1][7] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][7] ) );
  MUX41X1 U192 ( .IN1(\mat_i[0][1][8] ), .IN3(\mat_i[2][1][8] ), .IN2(
        \mat_i[1][1][8] ), .IN4(\mat_i[3][1][8] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][8] ) );
  MUX41X1 U193 ( .IN1(\mat_i[0][1][9] ), .IN3(\mat_i[2][1][9] ), .IN2(
        \mat_i[1][1][9] ), .IN4(\mat_i[3][1][9] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][9] ) );
  MUX41X1 U194 ( .IN1(\mat_i[0][1][10] ), .IN3(\mat_i[2][1][10] ), .IN2(
        \mat_i[1][1][10] ), .IN4(\mat_i[3][1][10] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][10] ) );
  MUX41X1 U195 ( .IN1(\mat_i[0][1][11] ), .IN3(\mat_i[2][1][11] ), .IN2(
        \mat_i[1][1][11] ), .IN4(\mat_i[3][1][11] ), .S0(n407), .S1(n415), .Q(
        \vector_out_i2[1][11] ) );
  MUX41X1 U196 ( .IN1(\mat_i[0][0][0] ), .IN3(\mat_i[2][0][0] ), .IN2(
        \mat_i[1][0][0] ), .IN4(\mat_i[3][0][0] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][0] ) );
  MUX41X1 U197 ( .IN1(\mat_i[0][0][1] ), .IN3(\mat_i[2][0][1] ), .IN2(
        \mat_i[1][0][1] ), .IN4(\mat_i[3][0][1] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][1] ) );
  MUX41X1 U198 ( .IN1(\mat_i[0][0][2] ), .IN3(\mat_i[2][0][2] ), .IN2(
        \mat_i[1][0][2] ), .IN4(\mat_i[3][0][2] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][2] ) );
  MUX41X1 U199 ( .IN1(\mat_i[0][0][3] ), .IN3(\mat_i[2][0][3] ), .IN2(
        \mat_i[1][0][3] ), .IN4(\mat_i[3][0][3] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][3] ) );
  MUX41X1 U200 ( .IN1(\mat_i[0][0][4] ), .IN3(\mat_i[2][0][4] ), .IN2(
        \mat_i[1][0][4] ), .IN4(\mat_i[3][0][4] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][4] ) );
  MUX41X1 U201 ( .IN1(\mat_i[0][0][5] ), .IN3(\mat_i[2][0][5] ), .IN2(
        \mat_i[1][0][5] ), .IN4(\mat_i[3][0][5] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][5] ) );
  MUX41X1 U202 ( .IN1(\mat_i[0][0][6] ), .IN3(\mat_i[2][0][6] ), .IN2(
        \mat_i[1][0][6] ), .IN4(\mat_i[3][0][6] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][6] ) );
  MUX41X1 U203 ( .IN1(\mat_i[0][0][7] ), .IN3(\mat_i[2][0][7] ), .IN2(
        \mat_i[1][0][7] ), .IN4(\mat_i[3][0][7] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][7] ) );
  MUX41X1 U204 ( .IN1(\mat_i[0][0][8] ), .IN3(\mat_i[2][0][8] ), .IN2(
        \mat_i[1][0][8] ), .IN4(\mat_i[3][0][8] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][8] ) );
  MUX41X1 U205 ( .IN1(\mat_i[0][0][9] ), .IN3(\mat_i[2][0][9] ), .IN2(
        \mat_i[1][0][9] ), .IN4(\mat_i[3][0][9] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][9] ) );
  MUX41X1 U206 ( .IN1(\mat_i[0][0][10] ), .IN3(\mat_i[2][0][10] ), .IN2(
        \mat_i[1][0][10] ), .IN4(\mat_i[3][0][10] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][10] ) );
  MUX41X1 U207 ( .IN1(\mat_i[0][0][11] ), .IN3(\mat_i[2][0][11] ), .IN2(
        \mat_i[1][0][11] ), .IN4(\mat_i[3][0][11] ), .S0(n408), .S1(n416), .Q(
        \vector_out_i2[0][11] ) );
  MUX41X1 U208 ( .IN1(\mat_r[0][3][0] ), .IN3(\mat_r[2][3][0] ), .IN2(
        \mat_r[1][3][0] ), .IN4(\mat_r[3][3][0] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][0] ) );
  MUX41X1 U209 ( .IN1(\mat_r[0][3][1] ), .IN3(\mat_r[2][3][1] ), .IN2(
        \mat_r[1][3][1] ), .IN4(\mat_r[3][3][1] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][1] ) );
  MUX41X1 U210 ( .IN1(\mat_r[0][3][2] ), .IN3(\mat_r[2][3][2] ), .IN2(
        \mat_r[1][3][2] ), .IN4(\mat_r[3][3][2] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][2] ) );
  MUX41X1 U211 ( .IN1(\mat_r[0][3][3] ), .IN3(\mat_r[2][3][3] ), .IN2(
        \mat_r[1][3][3] ), .IN4(\mat_r[3][3][3] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][3] ) );
  MUX41X1 U212 ( .IN1(\mat_r[0][3][4] ), .IN3(\mat_r[2][3][4] ), .IN2(
        \mat_r[1][3][4] ), .IN4(\mat_r[3][3][4] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][4] ) );
  MUX41X1 U213 ( .IN1(\mat_r[0][3][5] ), .IN3(\mat_r[2][3][5] ), .IN2(
        \mat_r[1][3][5] ), .IN4(\mat_r[3][3][5] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][5] ) );
  MUX41X1 U214 ( .IN1(\mat_r[0][3][6] ), .IN3(\mat_r[2][3][6] ), .IN2(
        \mat_r[1][3][6] ), .IN4(\mat_r[3][3][6] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][6] ) );
  MUX41X1 U215 ( .IN1(\mat_r[0][3][7] ), .IN3(\mat_r[2][3][7] ), .IN2(
        \mat_r[1][3][7] ), .IN4(\mat_r[3][3][7] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][7] ) );
  MUX41X1 U216 ( .IN1(\mat_r[0][3][8] ), .IN3(\mat_r[2][3][8] ), .IN2(
        \mat_r[1][3][8] ), .IN4(\mat_r[3][3][8] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][8] ) );
  MUX41X1 U217 ( .IN1(\mat_r[0][3][9] ), .IN3(\mat_r[2][3][9] ), .IN2(
        \mat_r[1][3][9] ), .IN4(\mat_r[3][3][9] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][9] ) );
  MUX41X1 U218 ( .IN1(\mat_r[0][3][10] ), .IN3(\mat_r[2][3][10] ), .IN2(
        \mat_r[1][3][10] ), .IN4(\mat_r[3][3][10] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][10] ) );
  MUX41X1 U219 ( .IN1(\mat_r[0][3][11] ), .IN3(\mat_r[2][3][11] ), .IN2(
        \mat_r[1][3][11] ), .IN4(\mat_r[3][3][11] ), .S0(n409), .S1(n417), .Q(
        \vector_out_r2[3][11] ) );
  MUX41X1 U220 ( .IN1(\mat_r[0][2][0] ), .IN3(\mat_r[2][2][0] ), .IN2(
        \mat_r[1][2][0] ), .IN4(\mat_r[3][2][0] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][0] ) );
  MUX41X1 U221 ( .IN1(\mat_r[0][2][1] ), .IN3(\mat_r[2][2][1] ), .IN2(
        \mat_r[1][2][1] ), .IN4(\mat_r[3][2][1] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][1] ) );
  MUX41X1 U222 ( .IN1(\mat_r[0][2][2] ), .IN3(\mat_r[2][2][2] ), .IN2(
        \mat_r[1][2][2] ), .IN4(\mat_r[3][2][2] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][2] ) );
  MUX41X1 U223 ( .IN1(\mat_r[0][2][3] ), .IN3(\mat_r[2][2][3] ), .IN2(
        \mat_r[1][2][3] ), .IN4(\mat_r[3][2][3] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][3] ) );
  MUX41X1 U224 ( .IN1(\mat_r[0][2][4] ), .IN3(\mat_r[2][2][4] ), .IN2(
        \mat_r[1][2][4] ), .IN4(\mat_r[3][2][4] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][4] ) );
  MUX41X1 U225 ( .IN1(\mat_r[0][2][5] ), .IN3(\mat_r[2][2][5] ), .IN2(
        \mat_r[1][2][5] ), .IN4(\mat_r[3][2][5] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][5] ) );
  MUX41X1 U226 ( .IN1(\mat_r[0][2][6] ), .IN3(\mat_r[2][2][6] ), .IN2(
        \mat_r[1][2][6] ), .IN4(\mat_r[3][2][6] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][6] ) );
  MUX41X1 U227 ( .IN1(\mat_r[0][2][7] ), .IN3(\mat_r[2][2][7] ), .IN2(
        \mat_r[1][2][7] ), .IN4(\mat_r[3][2][7] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][7] ) );
  MUX41X1 U228 ( .IN1(\mat_r[0][2][8] ), .IN3(\mat_r[2][2][8] ), .IN2(
        \mat_r[1][2][8] ), .IN4(\mat_r[3][2][8] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][8] ) );
  MUX41X1 U229 ( .IN1(\mat_r[0][2][9] ), .IN3(\mat_r[2][2][9] ), .IN2(
        \mat_r[1][2][9] ), .IN4(\mat_r[3][2][9] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][9] ) );
  MUX41X1 U230 ( .IN1(\mat_r[0][2][10] ), .IN3(\mat_r[2][2][10] ), .IN2(
        \mat_r[1][2][10] ), .IN4(\mat_r[3][2][10] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][10] ) );
  MUX41X1 U231 ( .IN1(\mat_r[0][2][11] ), .IN3(\mat_r[2][2][11] ), .IN2(
        \mat_r[1][2][11] ), .IN4(\mat_r[3][2][11] ), .S0(n410), .S1(n418), .Q(
        \vector_out_r2[2][11] ) );
  MUX41X1 U232 ( .IN1(\mat_r[0][1][0] ), .IN3(\mat_r[2][1][0] ), .IN2(
        \mat_r[1][1][0] ), .IN4(\mat_r[3][1][0] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][0] ) );
  MUX41X1 U233 ( .IN1(\mat_r[0][1][1] ), .IN3(\mat_r[2][1][1] ), .IN2(
        \mat_r[1][1][1] ), .IN4(\mat_r[3][1][1] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][1] ) );
  MUX41X1 U234 ( .IN1(\mat_r[0][1][2] ), .IN3(\mat_r[2][1][2] ), .IN2(
        \mat_r[1][1][2] ), .IN4(\mat_r[3][1][2] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][2] ) );
  MUX41X1 U235 ( .IN1(\mat_r[0][1][3] ), .IN3(\mat_r[2][1][3] ), .IN2(
        \mat_r[1][1][3] ), .IN4(\mat_r[3][1][3] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][3] ) );
  MUX41X1 U236 ( .IN1(\mat_r[0][1][4] ), .IN3(\mat_r[2][1][4] ), .IN2(
        \mat_r[1][1][4] ), .IN4(\mat_r[3][1][4] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][4] ) );
  MUX41X1 U237 ( .IN1(\mat_r[0][1][5] ), .IN3(\mat_r[2][1][5] ), .IN2(
        \mat_r[1][1][5] ), .IN4(\mat_r[3][1][5] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][5] ) );
  MUX41X1 U238 ( .IN1(\mat_r[0][1][6] ), .IN3(\mat_r[2][1][6] ), .IN2(
        \mat_r[1][1][6] ), .IN4(\mat_r[3][1][6] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][6] ) );
  MUX41X1 U239 ( .IN1(\mat_r[0][1][7] ), .IN3(\mat_r[2][1][7] ), .IN2(
        \mat_r[1][1][7] ), .IN4(\mat_r[3][1][7] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][7] ) );
  MUX41X1 U240 ( .IN1(\mat_r[0][1][8] ), .IN3(\mat_r[2][1][8] ), .IN2(
        \mat_r[1][1][8] ), .IN4(\mat_r[3][1][8] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][8] ) );
  MUX41X1 U241 ( .IN1(\mat_r[0][1][9] ), .IN3(\mat_r[2][1][9] ), .IN2(
        \mat_r[1][1][9] ), .IN4(\mat_r[3][1][9] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][9] ) );
  MUX41X1 U242 ( .IN1(\mat_r[0][1][10] ), .IN3(\mat_r[2][1][10] ), .IN2(
        \mat_r[1][1][10] ), .IN4(\mat_r[3][1][10] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][10] ) );
  MUX41X1 U243 ( .IN1(\mat_r[0][1][11] ), .IN3(\mat_r[2][1][11] ), .IN2(
        \mat_r[1][1][11] ), .IN4(\mat_r[3][1][11] ), .S0(n411), .S1(n419), .Q(
        \vector_out_r2[1][11] ) );
  MUX41X1 U244 ( .IN1(\mat_r[0][0][0] ), .IN3(\mat_r[2][0][0] ), .IN2(
        \mat_r[1][0][0] ), .IN4(\mat_r[3][0][0] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][0] ) );
  MUX41X1 U245 ( .IN1(\mat_r[0][0][1] ), .IN3(\mat_r[2][0][1] ), .IN2(
        \mat_r[1][0][1] ), .IN4(\mat_r[3][0][1] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][1] ) );
  MUX41X1 U246 ( .IN1(\mat_r[0][0][2] ), .IN3(\mat_r[2][0][2] ), .IN2(
        \mat_r[1][0][2] ), .IN4(\mat_r[3][0][2] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][2] ) );
  MUX41X1 U247 ( .IN1(\mat_r[0][0][3] ), .IN3(\mat_r[2][0][3] ), .IN2(
        \mat_r[1][0][3] ), .IN4(\mat_r[3][0][3] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][3] ) );
  MUX41X1 U248 ( .IN1(\mat_r[0][0][4] ), .IN3(\mat_r[2][0][4] ), .IN2(
        \mat_r[1][0][4] ), .IN4(\mat_r[3][0][4] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][4] ) );
  MUX41X1 U249 ( .IN1(\mat_r[0][0][5] ), .IN3(\mat_r[2][0][5] ), .IN2(
        \mat_r[1][0][5] ), .IN4(\mat_r[3][0][5] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][5] ) );
  MUX41X1 U250 ( .IN1(\mat_r[0][0][6] ), .IN3(\mat_r[2][0][6] ), .IN2(
        \mat_r[1][0][6] ), .IN4(\mat_r[3][0][6] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][6] ) );
  MUX41X1 U251 ( .IN1(\mat_r[0][0][7] ), .IN3(\mat_r[2][0][7] ), .IN2(
        \mat_r[1][0][7] ), .IN4(\mat_r[3][0][7] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][7] ) );
  MUX41X1 U252 ( .IN1(\mat_r[0][0][8] ), .IN3(\mat_r[2][0][8] ), .IN2(
        \mat_r[1][0][8] ), .IN4(\mat_r[3][0][8] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][8] ) );
  MUX41X1 U253 ( .IN1(\mat_r[0][0][9] ), .IN3(\mat_r[2][0][9] ), .IN2(
        \mat_r[1][0][9] ), .IN4(\mat_r[3][0][9] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][9] ) );
  MUX41X1 U254 ( .IN1(\mat_r[0][0][10] ), .IN3(\mat_r[2][0][10] ), .IN2(
        \mat_r[1][0][10] ), .IN4(\mat_r[3][0][10] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][10] ) );
  MUX41X1 U255 ( .IN1(\mat_r[0][0][11] ), .IN3(\mat_r[2][0][11] ), .IN2(
        \mat_r[1][0][11] ), .IN4(\mat_r[3][0][11] ), .S0(n412), .S1(n420), .Q(
        \vector_out_r2[0][11] ) );
  DELLN2X2 U256 ( .INP(N9), .Z(n405) );
  DELLN2X2 U257 ( .INP(N9), .Z(n406) );
  DELLN2X2 U258 ( .INP(N9), .Z(n407) );
  DELLN2X2 U259 ( .INP(N9), .Z(n408) );
  DELLN2X2 U260 ( .INP(N9), .Z(n409) );
  DELLN2X2 U261 ( .INP(N9), .Z(n410) );
  DELLN2X2 U262 ( .INP(N9), .Z(n411) );
  DELLN2X2 U263 ( .INP(N9), .Z(n412) );
  DELLN1X2 U264 ( .INP(N8), .Z(n413) );
  DELLN1X2 U265 ( .INP(N8), .Z(n414) );
  DELLN1X2 U266 ( .INP(N8), .Z(n415) );
  DELLN1X2 U267 ( .INP(N8), .Z(n416) );
  DELLN1X2 U268 ( .INP(N8), .Z(n417) );
  DELLN1X2 U269 ( .INP(N8), .Z(n418) );
  DELLN1X2 U270 ( .INP(N8), .Z(n419) );
  DELLN1X2 U271 ( .INP(N8), .Z(n420) );
  MUX41X1 U272 ( .IN1(\vector_out_i[0][0] ), .IN3(\vector_out_i[2][0] ), .IN2(
        \vector_out_i[1][0] ), .IN4(\vector_out_i[3][0] ), .S0(n421), .S1(n423), .Q(single_out_i[0]) );
  MUX41X1 U273 ( .IN1(\vector_out_i[0][1] ), .IN3(\vector_out_i[2][1] ), .IN2(
        \vector_out_i[1][1] ), .IN4(\vector_out_i[3][1] ), .S0(n421), .S1(n423), .Q(single_out_i[1]) );
  MUX41X1 U274 ( .IN1(\vector_out_i[0][2] ), .IN3(\vector_out_i[2][2] ), .IN2(
        \vector_out_i[1][2] ), .IN4(\vector_out_i[3][2] ), .S0(n421), .S1(n423), .Q(single_out_i[2]) );
  MUX41X1 U275 ( .IN1(\vector_out_i[0][3] ), .IN3(\vector_out_i[2][3] ), .IN2(
        \vector_out_i[1][3] ), .IN4(\vector_out_i[3][3] ), .S0(n421), .S1(n423), .Q(single_out_i[3]) );
  MUX41X1 U276 ( .IN1(\vector_out_i[0][4] ), .IN3(\vector_out_i[2][4] ), .IN2(
        \vector_out_i[1][4] ), .IN4(\vector_out_i[3][4] ), .S0(n421), .S1(n423), .Q(single_out_i[4]) );
  MUX41X1 U277 ( .IN1(\vector_out_i[0][5] ), .IN3(\vector_out_i[2][5] ), .IN2(
        \vector_out_i[1][5] ), .IN4(\vector_out_i[3][5] ), .S0(n421), .S1(n423), .Q(single_out_i[5]) );
  MUX41X1 U278 ( .IN1(\vector_out_i[0][6] ), .IN3(\vector_out_i[2][6] ), .IN2(
        \vector_out_i[1][6] ), .IN4(\vector_out_i[3][6] ), .S0(n421), .S1(n423), .Q(single_out_i[6]) );
  MUX41X1 U279 ( .IN1(\vector_out_i[0][7] ), .IN3(\vector_out_i[2][7] ), .IN2(
        \vector_out_i[1][7] ), .IN4(\vector_out_i[3][7] ), .S0(n421), .S1(n423), .Q(single_out_i[7]) );
  MUX41X1 U280 ( .IN1(\vector_out_i[0][8] ), .IN3(\vector_out_i[2][8] ), .IN2(
        \vector_out_i[1][8] ), .IN4(\vector_out_i[3][8] ), .S0(n421), .S1(n423), .Q(single_out_i[8]) );
  MUX41X1 U281 ( .IN1(\vector_out_i[0][9] ), .IN3(\vector_out_i[2][9] ), .IN2(
        \vector_out_i[1][9] ), .IN4(\vector_out_i[3][9] ), .S0(n421), .S1(n423), .Q(single_out_i[9]) );
  MUX41X1 U282 ( .IN1(\vector_out_i[0][10] ), .IN3(\vector_out_i[2][10] ), 
        .IN2(\vector_out_i[1][10] ), .IN4(\vector_out_i[3][10] ), .S0(n421), 
        .S1(n423), .Q(single_out_i[10]) );
  MUX41X1 U283 ( .IN1(\vector_out_i[0][11] ), .IN3(\vector_out_i[2][11] ), 
        .IN2(\vector_out_i[1][11] ), .IN4(\vector_out_i[3][11] ), .S0(n421), 
        .S1(n423), .Q(single_out_i[11]) );
  MUX41X1 U284 ( .IN1(\vector_out_r[0][0] ), .IN3(\vector_out_r[2][0] ), .IN2(
        \vector_out_r[1][0] ), .IN4(\vector_out_r[3][0] ), .S0(n422), .S1(n424), .Q(single_out_r[0]) );
  MUX41X1 U285 ( .IN1(\vector_out_r[0][1] ), .IN3(\vector_out_r[2][1] ), .IN2(
        \vector_out_r[1][1] ), .IN4(\vector_out_r[3][1] ), .S0(n422), .S1(n424), .Q(single_out_r[1]) );
  MUX41X1 U286 ( .IN1(\vector_out_r[0][2] ), .IN3(\vector_out_r[2][2] ), .IN2(
        \vector_out_r[1][2] ), .IN4(\vector_out_r[3][2] ), .S0(n422), .S1(n424), .Q(single_out_r[2]) );
  MUX41X1 U287 ( .IN1(\vector_out_r[0][3] ), .IN3(\vector_out_r[2][3] ), .IN2(
        \vector_out_r[1][3] ), .IN4(\vector_out_r[3][3] ), .S0(n422), .S1(n424), .Q(single_out_r[3]) );
  MUX41X1 U288 ( .IN1(\vector_out_r[0][4] ), .IN3(\vector_out_r[2][4] ), .IN2(
        \vector_out_r[1][4] ), .IN4(\vector_out_r[3][4] ), .S0(n422), .S1(n424), .Q(single_out_r[4]) );
  MUX41X1 U289 ( .IN1(\vector_out_r[0][5] ), .IN3(\vector_out_r[2][5] ), .IN2(
        \vector_out_r[1][5] ), .IN4(\vector_out_r[3][5] ), .S0(n422), .S1(n424), .Q(single_out_r[5]) );
  MUX41X1 U290 ( .IN1(\vector_out_r[0][6] ), .IN3(\vector_out_r[2][6] ), .IN2(
        \vector_out_r[1][6] ), .IN4(\vector_out_r[3][6] ), .S0(n422), .S1(n424), .Q(single_out_r[6]) );
  MUX41X1 U291 ( .IN1(\vector_out_r[0][7] ), .IN3(\vector_out_r[2][7] ), .IN2(
        \vector_out_r[1][7] ), .IN4(\vector_out_r[3][7] ), .S0(n422), .S1(n424), .Q(single_out_r[7]) );
  MUX41X1 U292 ( .IN1(\vector_out_r[0][8] ), .IN3(\vector_out_r[2][8] ), .IN2(
        \vector_out_r[1][8] ), .IN4(\vector_out_r[3][8] ), .S0(n422), .S1(n424), .Q(single_out_r[8]) );
  MUX41X1 U293 ( .IN1(\vector_out_r[0][9] ), .IN3(\vector_out_r[2][9] ), .IN2(
        \vector_out_r[1][9] ), .IN4(\vector_out_r[3][9] ), .S0(n422), .S1(n424), .Q(single_out_r[9]) );
  MUX41X1 U294 ( .IN1(\vector_out_r[0][10] ), .IN3(\vector_out_r[2][10] ), 
        .IN2(\vector_out_r[1][10] ), .IN4(\vector_out_r[3][10] ), .S0(n422), 
        .S1(n424), .Q(single_out_r[10]) );
  MUX41X1 U295 ( .IN1(\vector_out_r[0][11] ), .IN3(\vector_out_r[2][11] ), 
        .IN2(\vector_out_r[1][11] ), .IN4(\vector_out_r[3][11] ), .S0(n422), 
        .S1(n424), .Q(single_out_r[11]) );
  MUX41X1 U296 ( .IN1(\vector_out_i2[0][0] ), .IN3(\vector_out_i2[2][0] ), 
        .IN2(\vector_out_i2[1][0] ), .IN4(\vector_out_i2[3][0] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[0]) );
  MUX41X1 U297 ( .IN1(\vector_out_i2[0][1] ), .IN3(\vector_out_i2[2][1] ), 
        .IN2(\vector_out_i2[1][1] ), .IN4(\vector_out_i2[3][1] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[1]) );
  MUX41X1 U298 ( .IN1(\vector_out_i2[0][2] ), .IN3(\vector_out_i2[2][2] ), 
        .IN2(\vector_out_i2[1][2] ), .IN4(\vector_out_i2[3][2] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[2]) );
  MUX41X1 U299 ( .IN1(\vector_out_i2[0][3] ), .IN3(\vector_out_i2[2][3] ), 
        .IN2(\vector_out_i2[1][3] ), .IN4(\vector_out_i2[3][3] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[3]) );
  MUX41X1 U300 ( .IN1(\vector_out_i2[0][4] ), .IN3(\vector_out_i2[2][4] ), 
        .IN2(\vector_out_i2[1][4] ), .IN4(\vector_out_i2[3][4] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[4]) );
  MUX41X1 U301 ( .IN1(\vector_out_i2[0][5] ), .IN3(\vector_out_i2[2][5] ), 
        .IN2(\vector_out_i2[1][5] ), .IN4(\vector_out_i2[3][5] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[5]) );
  MUX41X1 U302 ( .IN1(\vector_out_i2[0][6] ), .IN3(\vector_out_i2[2][6] ), 
        .IN2(\vector_out_i2[1][6] ), .IN4(\vector_out_i2[3][6] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[6]) );
  MUX41X1 U303 ( .IN1(\vector_out_i2[0][7] ), .IN3(\vector_out_i2[2][7] ), 
        .IN2(\vector_out_i2[1][7] ), .IN4(\vector_out_i2[3][7] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[7]) );
  MUX41X1 U304 ( .IN1(\vector_out_i2[0][8] ), .IN3(\vector_out_i2[2][8] ), 
        .IN2(\vector_out_i2[1][8] ), .IN4(\vector_out_i2[3][8] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[8]) );
  MUX41X1 U305 ( .IN1(\vector_out_i2[0][9] ), .IN3(\vector_out_i2[2][9] ), 
        .IN2(\vector_out_i2[1][9] ), .IN4(\vector_out_i2[3][9] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[9]) );
  MUX41X1 U306 ( .IN1(\vector_out_i2[0][10] ), .IN3(\vector_out_i2[2][10] ), 
        .IN2(\vector_out_i2[1][10] ), .IN4(\vector_out_i2[3][10] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[10]) );
  MUX41X1 U307 ( .IN1(\vector_out_i2[0][11] ), .IN3(\vector_out_i2[2][11] ), 
        .IN2(\vector_out_i2[1][11] ), .IN4(\vector_out_i2[3][11] ), .S0(n425), 
        .S1(n427), .Q(single_out_i2[11]) );
  MUX41X1 U308 ( .IN1(\vector_out_r2[0][0] ), .IN3(\vector_out_r2[2][0] ), 
        .IN2(\vector_out_r2[1][0] ), .IN4(\vector_out_r2[3][0] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[0]) );
  MUX41X1 U309 ( .IN1(\vector_out_r2[0][1] ), .IN3(\vector_out_r2[2][1] ), 
        .IN2(\vector_out_r2[1][1] ), .IN4(\vector_out_r2[3][1] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[1]) );
  MUX41X1 U310 ( .IN1(\vector_out_r2[0][2] ), .IN3(\vector_out_r2[2][2] ), 
        .IN2(\vector_out_r2[1][2] ), .IN4(\vector_out_r2[3][2] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[2]) );
  MUX41X1 U311 ( .IN1(\vector_out_r2[0][3] ), .IN3(\vector_out_r2[2][3] ), 
        .IN2(\vector_out_r2[1][3] ), .IN4(\vector_out_r2[3][3] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[3]) );
  MUX41X1 U312 ( .IN1(\vector_out_r2[0][4] ), .IN3(\vector_out_r2[2][4] ), 
        .IN2(\vector_out_r2[1][4] ), .IN4(\vector_out_r2[3][4] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[4]) );
  MUX41X1 U313 ( .IN1(\vector_out_r2[0][5] ), .IN3(\vector_out_r2[2][5] ), 
        .IN2(\vector_out_r2[1][5] ), .IN4(\vector_out_r2[3][5] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[5]) );
  MUX41X1 U314 ( .IN1(\vector_out_r2[0][6] ), .IN3(\vector_out_r2[2][6] ), 
        .IN2(\vector_out_r2[1][6] ), .IN4(\vector_out_r2[3][6] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[6]) );
  MUX41X1 U315 ( .IN1(\vector_out_r2[0][7] ), .IN3(\vector_out_r2[2][7] ), 
        .IN2(\vector_out_r2[1][7] ), .IN4(\vector_out_r2[3][7] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[7]) );
  MUX41X1 U316 ( .IN1(\vector_out_r2[0][8] ), .IN3(\vector_out_r2[2][8] ), 
        .IN2(\vector_out_r2[1][8] ), .IN4(\vector_out_r2[3][8] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[8]) );
  MUX41X1 U317 ( .IN1(\vector_out_r2[0][9] ), .IN3(\vector_out_r2[2][9] ), 
        .IN2(\vector_out_r2[1][9] ), .IN4(\vector_out_r2[3][9] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[9]) );
  MUX41X1 U318 ( .IN1(\vector_out_r2[0][10] ), .IN3(\vector_out_r2[2][10] ), 
        .IN2(\vector_out_r2[1][10] ), .IN4(\vector_out_r2[3][10] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[10]) );
  MUX41X1 U319 ( .IN1(\vector_out_r2[0][11] ), .IN3(\vector_out_r2[2][11] ), 
        .IN2(\vector_out_r2[1][11] ), .IN4(\vector_out_r2[3][11] ), .S0(n426), 
        .S1(n428), .Q(single_out_r2[11]) );
  MUX21X1 U320 ( .IN1(\mat_i[0][3][0] ), .IN2(\vector_in_i[3][0] ), .S(n429), 
        .Q(n347) );
  MUX21X1 U321 ( .IN1(\mat_i[0][3][1] ), .IN2(\vector_in_i[3][1] ), .S(n429), 
        .Q(n348) );
  MUX21X1 U322 ( .IN1(\mat_i[0][3][2] ), .IN2(\vector_in_i[3][2] ), .S(n429), 
        .Q(n349) );
  MUX21X1 U323 ( .IN1(\mat_i[0][3][3] ), .IN2(\vector_in_i[3][3] ), .S(n429), 
        .Q(n350) );
  MUX21X1 U324 ( .IN1(\mat_i[0][3][4] ), .IN2(\vector_in_i[3][4] ), .S(n429), 
        .Q(n351) );
  MUX21X1 U325 ( .IN1(\mat_i[0][3][5] ), .IN2(\vector_in_i[3][5] ), .S(n429), 
        .Q(n352) );
  MUX21X1 U326 ( .IN1(\mat_i[0][3][6] ), .IN2(\vector_in_i[3][6] ), .S(n429), 
        .Q(n353) );
  MUX21X1 U327 ( .IN1(\mat_i[0][3][7] ), .IN2(\vector_in_i[3][7] ), .S(n429), 
        .Q(n354) );
  MUX21X1 U328 ( .IN1(\mat_i[0][3][8] ), .IN2(\vector_in_i[3][8] ), .S(n429), 
        .Q(n355) );
  MUX21X1 U329 ( .IN1(\mat_i[0][3][9] ), .IN2(\vector_in_i[3][9] ), .S(n429), 
        .Q(n356) );
  MUX21X1 U330 ( .IN1(\mat_i[0][3][10] ), .IN2(\vector_in_i[3][10] ), .S(n429), 
        .Q(n357) );
  MUX21X1 U331 ( .IN1(\mat_i[0][3][11] ), .IN2(\vector_in_i[3][11] ), .S(n429), 
        .Q(n358) );
  MUX21X1 U332 ( .IN1(\mat_i[0][2][0] ), .IN2(\vector_in_i[2][0] ), .S(n430), 
        .Q(n359) );
  MUX21X1 U333 ( .IN1(\mat_i[0][2][1] ), .IN2(\vector_in_i[2][1] ), .S(n430), 
        .Q(n360) );
  MUX21X1 U334 ( .IN1(\mat_i[0][2][2] ), .IN2(\vector_in_i[2][2] ), .S(n430), 
        .Q(n361) );
  MUX21X1 U335 ( .IN1(\mat_i[0][2][3] ), .IN2(\vector_in_i[2][3] ), .S(n430), 
        .Q(n362) );
  MUX21X1 U336 ( .IN1(\mat_i[0][2][4] ), .IN2(\vector_in_i[2][4] ), .S(n430), 
        .Q(n363) );
  MUX21X1 U337 ( .IN1(\mat_i[0][2][5] ), .IN2(\vector_in_i[2][5] ), .S(n430), 
        .Q(n364) );
  MUX21X1 U338 ( .IN1(\mat_i[0][2][6] ), .IN2(\vector_in_i[2][6] ), .S(n430), 
        .Q(n365) );
  MUX21X1 U339 ( .IN1(\mat_i[0][2][7] ), .IN2(\vector_in_i[2][7] ), .S(n430), 
        .Q(n366) );
  MUX21X1 U340 ( .IN1(\mat_i[0][2][8] ), .IN2(\vector_in_i[2][8] ), .S(n430), 
        .Q(n367) );
  MUX21X1 U341 ( .IN1(\mat_i[0][2][9] ), .IN2(\vector_in_i[2][9] ), .S(n430), 
        .Q(n368) );
  MUX21X1 U342 ( .IN1(\mat_i[0][2][10] ), .IN2(\vector_in_i[2][10] ), .S(n430), 
        .Q(n369) );
  MUX21X1 U343 ( .IN1(\mat_i[0][2][11] ), .IN2(\vector_in_i[2][11] ), .S(n430), 
        .Q(n370) );
  MUX21X1 U344 ( .IN1(\mat_i[0][1][0] ), .IN2(\vector_in_i[1][0] ), .S(n431), 
        .Q(n371) );
  MUX21X1 U345 ( .IN1(\mat_i[0][1][1] ), .IN2(\vector_in_i[1][1] ), .S(n431), 
        .Q(n372) );
  MUX21X1 U346 ( .IN1(\mat_i[0][1][2] ), .IN2(\vector_in_i[1][2] ), .S(n431), 
        .Q(n373) );
  MUX21X1 U347 ( .IN1(\mat_i[0][1][3] ), .IN2(\vector_in_i[1][3] ), .S(n431), 
        .Q(n374) );
  MUX21X1 U348 ( .IN1(\mat_i[0][1][4] ), .IN2(\vector_in_i[1][4] ), .S(n431), 
        .Q(n375) );
  MUX21X1 U349 ( .IN1(\mat_i[0][1][5] ), .IN2(\vector_in_i[1][5] ), .S(n431), 
        .Q(n376) );
  MUX21X1 U350 ( .IN1(\mat_i[0][1][6] ), .IN2(\vector_in_i[1][6] ), .S(n431), 
        .Q(n377) );
  MUX21X1 U351 ( .IN1(\mat_i[0][1][7] ), .IN2(\vector_in_i[1][7] ), .S(n431), 
        .Q(n378) );
  MUX21X1 U352 ( .IN1(\mat_i[0][1][8] ), .IN2(\vector_in_i[1][8] ), .S(n431), 
        .Q(n379) );
  MUX21X1 U353 ( .IN1(\mat_i[0][1][9] ), .IN2(\vector_in_i[1][9] ), .S(n431), 
        .Q(n380) );
  MUX21X1 U354 ( .IN1(\mat_i[0][1][10] ), .IN2(\vector_in_i[1][10] ), .S(n431), 
        .Q(n381) );
  MUX21X1 U355 ( .IN1(\mat_i[0][1][11] ), .IN2(\vector_in_i[1][11] ), .S(n431), 
        .Q(n382) );
  MUX21X1 U356 ( .IN1(\mat_i[0][0][0] ), .IN2(\vector_in_i[0][0] ), .S(n432), 
        .Q(n383) );
  MUX21X1 U357 ( .IN1(\mat_i[0][0][1] ), .IN2(\vector_in_i[0][1] ), .S(n432), 
        .Q(n384) );
  MUX21X1 U358 ( .IN1(\mat_i[0][0][2] ), .IN2(\vector_in_i[0][2] ), .S(n432), 
        .Q(n385) );
  MUX21X1 U359 ( .IN1(\mat_i[0][0][3] ), .IN2(\vector_in_i[0][3] ), .S(n432), 
        .Q(n386) );
  MUX21X1 U360 ( .IN1(\mat_i[0][0][4] ), .IN2(\vector_in_i[0][4] ), .S(n432), 
        .Q(n387) );
  MUX21X1 U361 ( .IN1(\mat_i[0][0][5] ), .IN2(\vector_in_i[0][5] ), .S(n432), 
        .Q(n388) );
  MUX21X1 U362 ( .IN1(\mat_i[0][0][6] ), .IN2(\vector_in_i[0][6] ), .S(n432), 
        .Q(n389) );
  MUX21X1 U363 ( .IN1(\mat_i[0][0][7] ), .IN2(\vector_in_i[0][7] ), .S(n432), 
        .Q(n390) );
  MUX21X1 U364 ( .IN1(\mat_i[0][0][8] ), .IN2(\vector_in_i[0][8] ), .S(n432), 
        .Q(n391) );
  MUX21X1 U365 ( .IN1(\mat_i[0][0][9] ), .IN2(\vector_in_i[0][9] ), .S(n432), 
        .Q(n392) );
  MUX21X1 U366 ( .IN1(\mat_i[0][0][10] ), .IN2(\vector_in_i[0][10] ), .S(n432), 
        .Q(n393) );
  MUX21X1 U367 ( .IN1(\mat_i[0][0][11] ), .IN2(\vector_in_i[0][11] ), .S(n432), 
        .Q(n394) );
  MUX21X1 U368 ( .IN1(\mat_r[0][3][0] ), .IN2(\vector_in_r[3][0] ), .S(n433), 
        .Q(n155) );
  MUX21X1 U369 ( .IN1(\mat_r[0][3][1] ), .IN2(\vector_in_r[3][1] ), .S(n433), 
        .Q(n156) );
  MUX21X1 U370 ( .IN1(\mat_r[0][3][2] ), .IN2(\vector_in_r[3][2] ), .S(n433), 
        .Q(n157) );
  MUX21X1 U371 ( .IN1(\mat_r[0][3][3] ), .IN2(\vector_in_r[3][3] ), .S(n433), 
        .Q(n158) );
  MUX21X1 U372 ( .IN1(\mat_r[0][3][4] ), .IN2(\vector_in_r[3][4] ), .S(n433), 
        .Q(n159) );
  MUX21X1 U373 ( .IN1(\mat_r[0][3][5] ), .IN2(\vector_in_r[3][5] ), .S(n433), 
        .Q(n160) );
  MUX21X1 U374 ( .IN1(\mat_r[0][3][6] ), .IN2(\vector_in_r[3][6] ), .S(n433), 
        .Q(n161) );
  MUX21X1 U375 ( .IN1(\mat_r[0][3][7] ), .IN2(\vector_in_r[3][7] ), .S(n433), 
        .Q(n162) );
  MUX21X1 U376 ( .IN1(\mat_r[0][3][8] ), .IN2(\vector_in_r[3][8] ), .S(n433), 
        .Q(n163) );
  MUX21X1 U377 ( .IN1(\mat_r[0][3][9] ), .IN2(\vector_in_r[3][9] ), .S(n433), 
        .Q(n164) );
  MUX21X1 U378 ( .IN1(\mat_r[0][3][10] ), .IN2(\vector_in_r[3][10] ), .S(n433), 
        .Q(n165) );
  MUX21X1 U379 ( .IN1(\mat_r[0][3][11] ), .IN2(\vector_in_r[3][11] ), .S(n433), 
        .Q(n166) );
  MUX21X1 U380 ( .IN1(\mat_r[0][2][0] ), .IN2(\vector_in_r[2][0] ), .S(n434), 
        .Q(n167) );
  MUX21X1 U381 ( .IN1(\mat_r[0][2][1] ), .IN2(\vector_in_r[2][1] ), .S(n434), 
        .Q(n168) );
  MUX21X1 U382 ( .IN1(\mat_r[0][2][2] ), .IN2(\vector_in_r[2][2] ), .S(n434), 
        .Q(n169) );
  MUX21X1 U383 ( .IN1(\mat_r[0][2][3] ), .IN2(\vector_in_r[2][3] ), .S(n434), 
        .Q(n170) );
  MUX21X1 U384 ( .IN1(\mat_r[0][2][4] ), .IN2(\vector_in_r[2][4] ), .S(n434), 
        .Q(n171) );
  MUX21X1 U385 ( .IN1(\mat_r[0][2][5] ), .IN2(\vector_in_r[2][5] ), .S(n434), 
        .Q(n172) );
  MUX21X1 U386 ( .IN1(\mat_r[0][2][6] ), .IN2(\vector_in_r[2][6] ), .S(n434), 
        .Q(n173) );
  MUX21X1 U387 ( .IN1(\mat_r[0][2][7] ), .IN2(\vector_in_r[2][7] ), .S(n434), 
        .Q(n174) );
  MUX21X1 U388 ( .IN1(\mat_r[0][2][8] ), .IN2(\vector_in_r[2][8] ), .S(n434), 
        .Q(n175) );
  MUX21X1 U389 ( .IN1(\mat_r[0][2][9] ), .IN2(\vector_in_r[2][9] ), .S(n434), 
        .Q(n176) );
  MUX21X1 U390 ( .IN1(\mat_r[0][2][10] ), .IN2(\vector_in_r[2][10] ), .S(n434), 
        .Q(n177) );
  MUX21X1 U391 ( .IN1(\mat_r[0][2][11] ), .IN2(\vector_in_r[2][11] ), .S(n434), 
        .Q(n178) );
  MUX21X1 U392 ( .IN1(\mat_r[0][1][0] ), .IN2(\vector_in_r[1][0] ), .S(n435), 
        .Q(n179) );
  MUX21X1 U393 ( .IN1(\mat_r[0][1][1] ), .IN2(\vector_in_r[1][1] ), .S(n435), 
        .Q(n180) );
  MUX21X1 U394 ( .IN1(\mat_r[0][1][2] ), .IN2(\vector_in_r[1][2] ), .S(n435), 
        .Q(n181) );
  MUX21X1 U395 ( .IN1(\mat_r[0][1][3] ), .IN2(\vector_in_r[1][3] ), .S(n435), 
        .Q(n182) );
  MUX21X1 U396 ( .IN1(\mat_r[0][1][4] ), .IN2(\vector_in_r[1][4] ), .S(n435), 
        .Q(n183) );
  MUX21X1 U397 ( .IN1(\mat_r[0][1][5] ), .IN2(\vector_in_r[1][5] ), .S(n435), 
        .Q(n184) );
  MUX21X1 U398 ( .IN1(\mat_r[0][1][6] ), .IN2(\vector_in_r[1][6] ), .S(n435), 
        .Q(n185) );
  MUX21X1 U399 ( .IN1(\mat_r[0][1][7] ), .IN2(\vector_in_r[1][7] ), .S(n435), 
        .Q(n186) );
  MUX21X1 U400 ( .IN1(\mat_r[0][1][8] ), .IN2(\vector_in_r[1][8] ), .S(n435), 
        .Q(n187) );
  MUX21X1 U401 ( .IN1(\mat_r[0][1][9] ), .IN2(\vector_in_r[1][9] ), .S(n435), 
        .Q(n188) );
  MUX21X1 U402 ( .IN1(\mat_r[0][1][10] ), .IN2(\vector_in_r[1][10] ), .S(n435), 
        .Q(n189) );
  MUX21X1 U403 ( .IN1(\mat_r[0][1][11] ), .IN2(\vector_in_r[1][11] ), .S(n435), 
        .Q(n190) );
  MUX21X1 U404 ( .IN1(\mat_r[0][0][0] ), .IN2(\vector_in_r[0][0] ), .S(n436), 
        .Q(n191) );
  MUX21X1 U405 ( .IN1(\mat_r[0][0][1] ), .IN2(\vector_in_r[0][1] ), .S(n436), 
        .Q(n192) );
  MUX21X1 U406 ( .IN1(\mat_r[0][0][2] ), .IN2(\vector_in_r[0][2] ), .S(n436), 
        .Q(n193) );
  MUX21X1 U407 ( .IN1(\mat_r[0][0][3] ), .IN2(\vector_in_r[0][3] ), .S(n436), 
        .Q(n194) );
  MUX21X1 U408 ( .IN1(\mat_r[0][0][4] ), .IN2(\vector_in_r[0][4] ), .S(n436), 
        .Q(n195) );
  MUX21X1 U409 ( .IN1(\mat_r[0][0][5] ), .IN2(\vector_in_r[0][5] ), .S(n436), 
        .Q(n196) );
  MUX21X1 U410 ( .IN1(\mat_r[0][0][6] ), .IN2(\vector_in_r[0][6] ), .S(n436), 
        .Q(n197) );
  MUX21X1 U411 ( .IN1(\mat_r[0][0][7] ), .IN2(\vector_in_r[0][7] ), .S(n436), 
        .Q(n198) );
  MUX21X1 U412 ( .IN1(\mat_r[0][0][8] ), .IN2(\vector_in_r[0][8] ), .S(n436), 
        .Q(n199) );
  MUX21X1 U413 ( .IN1(\mat_r[0][0][9] ), .IN2(\vector_in_r[0][9] ), .S(n436), 
        .Q(n200) );
  MUX21X1 U414 ( .IN1(\mat_r[0][0][10] ), .IN2(\vector_in_r[0][10] ), .S(n436), 
        .Q(n201) );
  MUX21X1 U415 ( .IN1(\mat_r[0][0][11] ), .IN2(\vector_in_r[0][11] ), .S(n436), 
        .Q(n202) );
  MUX21X1 U416 ( .IN1(\mat_i[1][3][0] ), .IN2(\vector_in_i[3][0] ), .S(n437), 
        .Q(n299) );
  MUX21X1 U417 ( .IN1(\mat_i[1][3][1] ), .IN2(\vector_in_i[3][1] ), .S(n437), 
        .Q(n300) );
  MUX21X1 U418 ( .IN1(\mat_i[1][3][2] ), .IN2(\vector_in_i[3][2] ), .S(n437), 
        .Q(n301) );
  MUX21X1 U419 ( .IN1(\mat_i[1][3][3] ), .IN2(\vector_in_i[3][3] ), .S(n437), 
        .Q(n302) );
  MUX21X1 U420 ( .IN1(\mat_i[1][3][4] ), .IN2(\vector_in_i[3][4] ), .S(n437), 
        .Q(n303) );
  MUX21X1 U421 ( .IN1(\mat_i[1][3][5] ), .IN2(\vector_in_i[3][5] ), .S(n437), 
        .Q(n304) );
  MUX21X1 U422 ( .IN1(\mat_i[1][3][6] ), .IN2(\vector_in_i[3][6] ), .S(n437), 
        .Q(n305) );
  MUX21X1 U423 ( .IN1(\mat_i[1][3][7] ), .IN2(\vector_in_i[3][7] ), .S(n437), 
        .Q(n306) );
  MUX21X1 U424 ( .IN1(\mat_i[1][3][8] ), .IN2(\vector_in_i[3][8] ), .S(n437), 
        .Q(n307) );
  MUX21X1 U425 ( .IN1(\mat_i[1][3][9] ), .IN2(\vector_in_i[3][9] ), .S(n437), 
        .Q(n308) );
  MUX21X1 U426 ( .IN1(\mat_i[1][3][10] ), .IN2(\vector_in_i[3][10] ), .S(n437), 
        .Q(n309) );
  MUX21X1 U427 ( .IN1(\mat_i[1][3][11] ), .IN2(\vector_in_i[3][11] ), .S(n437), 
        .Q(n310) );
  MUX21X1 U428 ( .IN1(\mat_i[1][2][0] ), .IN2(\vector_in_i[2][0] ), .S(n438), 
        .Q(n311) );
  MUX21X1 U429 ( .IN1(\mat_i[1][2][1] ), .IN2(\vector_in_i[2][1] ), .S(n438), 
        .Q(n312) );
  MUX21X1 U430 ( .IN1(\mat_i[1][2][2] ), .IN2(\vector_in_i[2][2] ), .S(n438), 
        .Q(n313) );
  MUX21X1 U431 ( .IN1(\mat_i[1][2][3] ), .IN2(\vector_in_i[2][3] ), .S(n438), 
        .Q(n314) );
  MUX21X1 U432 ( .IN1(\mat_i[1][2][4] ), .IN2(\vector_in_i[2][4] ), .S(n438), 
        .Q(n315) );
  MUX21X1 U433 ( .IN1(\mat_i[1][2][5] ), .IN2(\vector_in_i[2][5] ), .S(n438), 
        .Q(n316) );
  MUX21X1 U434 ( .IN1(\mat_i[1][2][6] ), .IN2(\vector_in_i[2][6] ), .S(n438), 
        .Q(n317) );
  MUX21X1 U435 ( .IN1(\mat_i[1][2][7] ), .IN2(\vector_in_i[2][7] ), .S(n438), 
        .Q(n318) );
  MUX21X1 U436 ( .IN1(\mat_i[1][2][8] ), .IN2(\vector_in_i[2][8] ), .S(n438), 
        .Q(n319) );
  MUX21X1 U437 ( .IN1(\mat_i[1][2][9] ), .IN2(\vector_in_i[2][9] ), .S(n438), 
        .Q(n320) );
  MUX21X1 U438 ( .IN1(\mat_i[1][2][10] ), .IN2(\vector_in_i[2][10] ), .S(n438), 
        .Q(n321) );
  MUX21X1 U439 ( .IN1(\mat_i[1][2][11] ), .IN2(\vector_in_i[2][11] ), .S(n438), 
        .Q(n322) );
  MUX21X1 U440 ( .IN1(\mat_i[1][1][0] ), .IN2(\vector_in_i[1][0] ), .S(n439), 
        .Q(n323) );
  MUX21X1 U441 ( .IN1(\mat_i[1][1][1] ), .IN2(\vector_in_i[1][1] ), .S(n439), 
        .Q(n324) );
  MUX21X1 U442 ( .IN1(\mat_i[1][1][2] ), .IN2(\vector_in_i[1][2] ), .S(n439), 
        .Q(n325) );
  MUX21X1 U443 ( .IN1(\mat_i[1][1][3] ), .IN2(\vector_in_i[1][3] ), .S(n439), 
        .Q(n326) );
  MUX21X1 U444 ( .IN1(\mat_i[1][1][4] ), .IN2(\vector_in_i[1][4] ), .S(n439), 
        .Q(n327) );
  MUX21X1 U445 ( .IN1(\mat_i[1][1][5] ), .IN2(\vector_in_i[1][5] ), .S(n439), 
        .Q(n328) );
  MUX21X1 U446 ( .IN1(\mat_i[1][1][6] ), .IN2(\vector_in_i[1][6] ), .S(n439), 
        .Q(n329) );
  MUX21X1 U447 ( .IN1(\mat_i[1][1][7] ), .IN2(\vector_in_i[1][7] ), .S(n439), 
        .Q(n330) );
  MUX21X1 U448 ( .IN1(\mat_i[1][1][8] ), .IN2(\vector_in_i[1][8] ), .S(n439), 
        .Q(n331) );
  MUX21X1 U449 ( .IN1(\mat_i[1][1][9] ), .IN2(\vector_in_i[1][9] ), .S(n439), 
        .Q(n332) );
  MUX21X1 U450 ( .IN1(\mat_i[1][1][10] ), .IN2(\vector_in_i[1][10] ), .S(n439), 
        .Q(n333) );
  MUX21X1 U451 ( .IN1(\mat_i[1][1][11] ), .IN2(\vector_in_i[1][11] ), .S(n439), 
        .Q(n334) );
  MUX21X1 U452 ( .IN1(\mat_i[1][0][0] ), .IN2(\vector_in_i[0][0] ), .S(n440), 
        .Q(n335) );
  MUX21X1 U453 ( .IN1(\mat_i[1][0][1] ), .IN2(\vector_in_i[0][1] ), .S(n440), 
        .Q(n336) );
  MUX21X1 U454 ( .IN1(\mat_i[1][0][2] ), .IN2(\vector_in_i[0][2] ), .S(n440), 
        .Q(n337) );
  MUX21X1 U455 ( .IN1(\mat_i[1][0][3] ), .IN2(\vector_in_i[0][3] ), .S(n440), 
        .Q(n338) );
  MUX21X1 U456 ( .IN1(\mat_i[1][0][4] ), .IN2(\vector_in_i[0][4] ), .S(n440), 
        .Q(n339) );
  MUX21X1 U457 ( .IN1(\mat_i[1][0][5] ), .IN2(\vector_in_i[0][5] ), .S(n440), 
        .Q(n340) );
  MUX21X1 U458 ( .IN1(\mat_i[1][0][6] ), .IN2(\vector_in_i[0][6] ), .S(n440), 
        .Q(n341) );
  MUX21X1 U459 ( .IN1(\mat_i[1][0][7] ), .IN2(\vector_in_i[0][7] ), .S(n440), 
        .Q(n342) );
  MUX21X1 U460 ( .IN1(\mat_i[1][0][8] ), .IN2(\vector_in_i[0][8] ), .S(n440), 
        .Q(n343) );
  MUX21X1 U461 ( .IN1(\mat_i[1][0][9] ), .IN2(\vector_in_i[0][9] ), .S(n440), 
        .Q(n344) );
  MUX21X1 U462 ( .IN1(\mat_i[1][0][10] ), .IN2(\vector_in_i[0][10] ), .S(n440), 
        .Q(n345) );
  MUX21X1 U463 ( .IN1(\mat_i[1][0][11] ), .IN2(\vector_in_i[0][11] ), .S(n440), 
        .Q(n346) );
  MUX21X1 U464 ( .IN1(\mat_r[1][3][0] ), .IN2(\vector_in_r[3][0] ), .S(n441), 
        .Q(n107) );
  MUX21X1 U465 ( .IN1(\mat_r[1][3][1] ), .IN2(\vector_in_r[3][1] ), .S(n441), 
        .Q(n108) );
  MUX21X1 U466 ( .IN1(\mat_r[1][3][2] ), .IN2(\vector_in_r[3][2] ), .S(n441), 
        .Q(n109) );
  MUX21X1 U467 ( .IN1(\mat_r[1][3][3] ), .IN2(\vector_in_r[3][3] ), .S(n441), 
        .Q(n110) );
  MUX21X1 U468 ( .IN1(\mat_r[1][3][4] ), .IN2(\vector_in_r[3][4] ), .S(n441), 
        .Q(n111) );
  MUX21X1 U469 ( .IN1(\mat_r[1][3][5] ), .IN2(\vector_in_r[3][5] ), .S(n441), 
        .Q(n112) );
  MUX21X1 U470 ( .IN1(\mat_r[1][3][6] ), .IN2(\vector_in_r[3][6] ), .S(n441), 
        .Q(n113) );
  MUX21X1 U471 ( .IN1(\mat_r[1][3][7] ), .IN2(\vector_in_r[3][7] ), .S(n441), 
        .Q(n114) );
  MUX21X1 U472 ( .IN1(\mat_r[1][3][8] ), .IN2(\vector_in_r[3][8] ), .S(n441), 
        .Q(n115) );
  MUX21X1 U473 ( .IN1(\mat_r[1][3][9] ), .IN2(\vector_in_r[3][9] ), .S(n441), 
        .Q(n116) );
  MUX21X1 U474 ( .IN1(\mat_r[1][3][10] ), .IN2(\vector_in_r[3][10] ), .S(n441), 
        .Q(n117) );
  MUX21X1 U475 ( .IN1(\mat_r[1][3][11] ), .IN2(\vector_in_r[3][11] ), .S(n441), 
        .Q(n118) );
  MUX21X1 U476 ( .IN1(\mat_r[1][2][0] ), .IN2(\vector_in_r[2][0] ), .S(n442), 
        .Q(n119) );
  MUX21X1 U477 ( .IN1(\mat_r[1][2][1] ), .IN2(\vector_in_r[2][1] ), .S(n442), 
        .Q(n120) );
  MUX21X1 U478 ( .IN1(\mat_r[1][2][2] ), .IN2(\vector_in_r[2][2] ), .S(n442), 
        .Q(n121) );
  MUX21X1 U479 ( .IN1(\mat_r[1][2][3] ), .IN2(\vector_in_r[2][3] ), .S(n442), 
        .Q(n122) );
  MUX21X1 U480 ( .IN1(\mat_r[1][2][4] ), .IN2(\vector_in_r[2][4] ), .S(n442), 
        .Q(n123) );
  MUX21X1 U481 ( .IN1(\mat_r[1][2][5] ), .IN2(\vector_in_r[2][5] ), .S(n442), 
        .Q(n124) );
  MUX21X1 U482 ( .IN1(\mat_r[1][2][6] ), .IN2(\vector_in_r[2][6] ), .S(n442), 
        .Q(n125) );
  MUX21X1 U483 ( .IN1(\mat_r[1][2][7] ), .IN2(\vector_in_r[2][7] ), .S(n442), 
        .Q(n126) );
  MUX21X1 U484 ( .IN1(\mat_r[1][2][8] ), .IN2(\vector_in_r[2][8] ), .S(n442), 
        .Q(n127) );
  MUX21X1 U485 ( .IN1(\mat_r[1][2][9] ), .IN2(\vector_in_r[2][9] ), .S(n442), 
        .Q(n128) );
  MUX21X1 U486 ( .IN1(\mat_r[1][2][10] ), .IN2(\vector_in_r[2][10] ), .S(n442), 
        .Q(n129) );
  MUX21X1 U487 ( .IN1(\mat_r[1][2][11] ), .IN2(\vector_in_r[2][11] ), .S(n442), 
        .Q(n130) );
  MUX21X1 U488 ( .IN1(\mat_r[1][1][0] ), .IN2(\vector_in_r[1][0] ), .S(n443), 
        .Q(n131) );
  MUX21X1 U489 ( .IN1(\mat_r[1][1][1] ), .IN2(\vector_in_r[1][1] ), .S(n443), 
        .Q(n132) );
  MUX21X1 U490 ( .IN1(\mat_r[1][1][2] ), .IN2(\vector_in_r[1][2] ), .S(n443), 
        .Q(n133) );
  MUX21X1 U491 ( .IN1(\mat_r[1][1][3] ), .IN2(\vector_in_r[1][3] ), .S(n443), 
        .Q(n134) );
  MUX21X1 U492 ( .IN1(\mat_r[1][1][4] ), .IN2(\vector_in_r[1][4] ), .S(n443), 
        .Q(n135) );
  MUX21X1 U493 ( .IN1(\mat_r[1][1][5] ), .IN2(\vector_in_r[1][5] ), .S(n443), 
        .Q(n136) );
  MUX21X1 U494 ( .IN1(\mat_r[1][1][6] ), .IN2(\vector_in_r[1][6] ), .S(n443), 
        .Q(n137) );
  MUX21X1 U495 ( .IN1(\mat_r[1][1][7] ), .IN2(\vector_in_r[1][7] ), .S(n443), 
        .Q(n138) );
  MUX21X1 U496 ( .IN1(\mat_r[1][1][8] ), .IN2(\vector_in_r[1][8] ), .S(n443), 
        .Q(n139) );
  MUX21X1 U497 ( .IN1(\mat_r[1][1][9] ), .IN2(\vector_in_r[1][9] ), .S(n443), 
        .Q(n140) );
  MUX21X1 U498 ( .IN1(\mat_r[1][1][10] ), .IN2(\vector_in_r[1][10] ), .S(n443), 
        .Q(n141) );
  MUX21X1 U499 ( .IN1(\mat_r[1][1][11] ), .IN2(\vector_in_r[1][11] ), .S(n443), 
        .Q(n142) );
  MUX21X1 U500 ( .IN1(\mat_r[1][0][0] ), .IN2(\vector_in_r[0][0] ), .S(n444), 
        .Q(n143) );
  MUX21X1 U501 ( .IN1(\mat_r[1][0][1] ), .IN2(\vector_in_r[0][1] ), .S(n444), 
        .Q(n144) );
  MUX21X1 U502 ( .IN1(\mat_r[1][0][2] ), .IN2(\vector_in_r[0][2] ), .S(n444), 
        .Q(n145) );
  MUX21X1 U503 ( .IN1(\mat_r[1][0][3] ), .IN2(\vector_in_r[0][3] ), .S(n444), 
        .Q(n146) );
  MUX21X1 U504 ( .IN1(\mat_r[1][0][4] ), .IN2(\vector_in_r[0][4] ), .S(n444), 
        .Q(n147) );
  MUX21X1 U505 ( .IN1(\mat_r[1][0][5] ), .IN2(\vector_in_r[0][5] ), .S(n444), 
        .Q(n148) );
  MUX21X1 U506 ( .IN1(\mat_r[1][0][6] ), .IN2(\vector_in_r[0][6] ), .S(n444), 
        .Q(n149) );
  MUX21X1 U507 ( .IN1(\mat_r[1][0][7] ), .IN2(\vector_in_r[0][7] ), .S(n444), 
        .Q(n150) );
  MUX21X1 U508 ( .IN1(\mat_r[1][0][8] ), .IN2(\vector_in_r[0][8] ), .S(n444), 
        .Q(n151) );
  MUX21X1 U509 ( .IN1(\mat_r[1][0][9] ), .IN2(\vector_in_r[0][9] ), .S(n444), 
        .Q(n152) );
  MUX21X1 U510 ( .IN1(\mat_r[1][0][10] ), .IN2(\vector_in_r[0][10] ), .S(n444), 
        .Q(n153) );
  MUX21X1 U511 ( .IN1(\mat_r[1][0][11] ), .IN2(\vector_in_r[0][11] ), .S(n444), 
        .Q(n154) );
  MUX21X1 U512 ( .IN1(\mat_i[2][3][0] ), .IN2(\vector_in_i[3][0] ), .S(n445), 
        .Q(n251) );
  MUX21X1 U513 ( .IN1(\mat_i[2][3][1] ), .IN2(\vector_in_i[3][1] ), .S(n445), 
        .Q(n252) );
  MUX21X1 U514 ( .IN1(\mat_i[2][3][2] ), .IN2(\vector_in_i[3][2] ), .S(n445), 
        .Q(n253) );
  MUX21X1 U515 ( .IN1(\mat_i[2][3][3] ), .IN2(\vector_in_i[3][3] ), .S(n445), 
        .Q(n254) );
  MUX21X1 U516 ( .IN1(\mat_i[2][3][4] ), .IN2(\vector_in_i[3][4] ), .S(n445), 
        .Q(n255) );
  MUX21X1 U517 ( .IN1(\mat_i[2][3][5] ), .IN2(\vector_in_i[3][5] ), .S(n445), 
        .Q(n256) );
  MUX21X1 U518 ( .IN1(\mat_i[2][3][6] ), .IN2(\vector_in_i[3][6] ), .S(n445), 
        .Q(n257) );
  MUX21X1 U519 ( .IN1(\mat_i[2][3][7] ), .IN2(\vector_in_i[3][7] ), .S(n445), 
        .Q(n258) );
  MUX21X1 U520 ( .IN1(\mat_i[2][3][8] ), .IN2(\vector_in_i[3][8] ), .S(n445), 
        .Q(n259) );
  MUX21X1 U521 ( .IN1(\mat_i[2][3][9] ), .IN2(\vector_in_i[3][9] ), .S(n445), 
        .Q(n260) );
  MUX21X1 U522 ( .IN1(\mat_i[2][3][10] ), .IN2(\vector_in_i[3][10] ), .S(n445), 
        .Q(n261) );
  MUX21X1 U523 ( .IN1(\mat_i[2][3][11] ), .IN2(\vector_in_i[3][11] ), .S(n445), 
        .Q(n262) );
  MUX21X1 U524 ( .IN1(\mat_i[2][2][0] ), .IN2(\vector_in_i[2][0] ), .S(n446), 
        .Q(n263) );
  MUX21X1 U525 ( .IN1(\mat_i[2][2][1] ), .IN2(\vector_in_i[2][1] ), .S(n446), 
        .Q(n264) );
  MUX21X1 U526 ( .IN1(\mat_i[2][2][2] ), .IN2(\vector_in_i[2][2] ), .S(n446), 
        .Q(n265) );
  MUX21X1 U527 ( .IN1(\mat_i[2][2][3] ), .IN2(\vector_in_i[2][3] ), .S(n446), 
        .Q(n266) );
  MUX21X1 U528 ( .IN1(\mat_i[2][2][4] ), .IN2(\vector_in_i[2][4] ), .S(n446), 
        .Q(n267) );
  MUX21X1 U529 ( .IN1(\mat_i[2][2][5] ), .IN2(\vector_in_i[2][5] ), .S(n446), 
        .Q(n268) );
  MUX21X1 U530 ( .IN1(\mat_i[2][2][6] ), .IN2(\vector_in_i[2][6] ), .S(n446), 
        .Q(n269) );
  MUX21X1 U531 ( .IN1(\mat_i[2][2][7] ), .IN2(\vector_in_i[2][7] ), .S(n446), 
        .Q(n270) );
  MUX21X1 U532 ( .IN1(\mat_i[2][2][8] ), .IN2(\vector_in_i[2][8] ), .S(n446), 
        .Q(n271) );
  MUX21X1 U533 ( .IN1(\mat_i[2][2][9] ), .IN2(\vector_in_i[2][9] ), .S(n446), 
        .Q(n272) );
  MUX21X1 U534 ( .IN1(\mat_i[2][2][10] ), .IN2(\vector_in_i[2][10] ), .S(n446), 
        .Q(n273) );
  MUX21X1 U535 ( .IN1(\mat_i[2][2][11] ), .IN2(\vector_in_i[2][11] ), .S(n446), 
        .Q(n274) );
  MUX21X1 U536 ( .IN1(\mat_i[2][1][0] ), .IN2(\vector_in_i[1][0] ), .S(n447), 
        .Q(n275) );
  MUX21X1 U537 ( .IN1(\mat_i[2][1][1] ), .IN2(\vector_in_i[1][1] ), .S(n447), 
        .Q(n276) );
  MUX21X1 U538 ( .IN1(\mat_i[2][1][2] ), .IN2(\vector_in_i[1][2] ), .S(n447), 
        .Q(n277) );
  MUX21X1 U539 ( .IN1(\mat_i[2][1][3] ), .IN2(\vector_in_i[1][3] ), .S(n447), 
        .Q(n278) );
  MUX21X1 U540 ( .IN1(\mat_i[2][1][4] ), .IN2(\vector_in_i[1][4] ), .S(n447), 
        .Q(n279) );
  MUX21X1 U541 ( .IN1(\mat_i[2][1][5] ), .IN2(\vector_in_i[1][5] ), .S(n447), 
        .Q(n280) );
  MUX21X1 U542 ( .IN1(\mat_i[2][1][6] ), .IN2(\vector_in_i[1][6] ), .S(n447), 
        .Q(n281) );
  MUX21X1 U543 ( .IN1(\mat_i[2][1][7] ), .IN2(\vector_in_i[1][7] ), .S(n447), 
        .Q(n282) );
  MUX21X1 U544 ( .IN1(\mat_i[2][1][8] ), .IN2(\vector_in_i[1][8] ), .S(n447), 
        .Q(n283) );
  MUX21X1 U545 ( .IN1(\mat_i[2][1][9] ), .IN2(\vector_in_i[1][9] ), .S(n447), 
        .Q(n284) );
  MUX21X1 U546 ( .IN1(\mat_i[2][1][10] ), .IN2(\vector_in_i[1][10] ), .S(n447), 
        .Q(n285) );
  MUX21X1 U547 ( .IN1(\mat_i[2][1][11] ), .IN2(\vector_in_i[1][11] ), .S(n447), 
        .Q(n286) );
  MUX21X1 U548 ( .IN1(\mat_i[2][0][0] ), .IN2(\vector_in_i[0][0] ), .S(n448), 
        .Q(n287) );
  MUX21X1 U549 ( .IN1(\mat_i[2][0][1] ), .IN2(\vector_in_i[0][1] ), .S(n448), 
        .Q(n288) );
  MUX21X1 U550 ( .IN1(\mat_i[2][0][2] ), .IN2(\vector_in_i[0][2] ), .S(n448), 
        .Q(n289) );
  MUX21X1 U551 ( .IN1(\mat_i[2][0][3] ), .IN2(\vector_in_i[0][3] ), .S(n448), 
        .Q(n290) );
  MUX21X1 U552 ( .IN1(\mat_i[2][0][4] ), .IN2(\vector_in_i[0][4] ), .S(n448), 
        .Q(n291) );
  MUX21X1 U553 ( .IN1(\mat_i[2][0][5] ), .IN2(\vector_in_i[0][5] ), .S(n448), 
        .Q(n292) );
  MUX21X1 U554 ( .IN1(\mat_i[2][0][6] ), .IN2(\vector_in_i[0][6] ), .S(n448), 
        .Q(n293) );
  MUX21X1 U555 ( .IN1(\mat_i[2][0][7] ), .IN2(\vector_in_i[0][7] ), .S(n448), 
        .Q(n294) );
  MUX21X1 U556 ( .IN1(\mat_i[2][0][8] ), .IN2(\vector_in_i[0][8] ), .S(n448), 
        .Q(n295) );
  MUX21X1 U557 ( .IN1(\mat_i[2][0][9] ), .IN2(\vector_in_i[0][9] ), .S(n448), 
        .Q(n296) );
  MUX21X1 U558 ( .IN1(\mat_i[2][0][10] ), .IN2(\vector_in_i[0][10] ), .S(n448), 
        .Q(n297) );
  MUX21X1 U559 ( .IN1(\mat_i[2][0][11] ), .IN2(\vector_in_i[0][11] ), .S(n448), 
        .Q(n298) );
  MUX21X1 U560 ( .IN1(\mat_r[2][3][0] ), .IN2(\vector_in_r[3][0] ), .S(n449), 
        .Q(n59) );
  MUX21X1 U561 ( .IN1(\mat_r[2][3][1] ), .IN2(\vector_in_r[3][1] ), .S(n449), 
        .Q(n60) );
  MUX21X1 U562 ( .IN1(\mat_r[2][3][2] ), .IN2(\vector_in_r[3][2] ), .S(n449), 
        .Q(n61) );
  MUX21X1 U563 ( .IN1(\mat_r[2][3][3] ), .IN2(\vector_in_r[3][3] ), .S(n449), 
        .Q(n62) );
  MUX21X1 U564 ( .IN1(\mat_r[2][3][4] ), .IN2(\vector_in_r[3][4] ), .S(n449), 
        .Q(n63) );
  MUX21X1 U565 ( .IN1(\mat_r[2][3][5] ), .IN2(\vector_in_r[3][5] ), .S(n449), 
        .Q(n64) );
  MUX21X1 U566 ( .IN1(\mat_r[2][3][6] ), .IN2(\vector_in_r[3][6] ), .S(n449), 
        .Q(n65) );
  MUX21X1 U567 ( .IN1(\mat_r[2][3][7] ), .IN2(\vector_in_r[3][7] ), .S(n449), 
        .Q(n66) );
  MUX21X1 U568 ( .IN1(\mat_r[2][3][8] ), .IN2(\vector_in_r[3][8] ), .S(n449), 
        .Q(n67) );
  MUX21X1 U569 ( .IN1(\mat_r[2][3][9] ), .IN2(\vector_in_r[3][9] ), .S(n449), 
        .Q(n68) );
  MUX21X1 U570 ( .IN1(\mat_r[2][3][10] ), .IN2(\vector_in_r[3][10] ), .S(n449), 
        .Q(n69) );
  MUX21X1 U571 ( .IN1(\mat_r[2][3][11] ), .IN2(\vector_in_r[3][11] ), .S(n449), 
        .Q(n70) );
  MUX21X1 U572 ( .IN1(\mat_r[2][2][0] ), .IN2(\vector_in_r[2][0] ), .S(n450), 
        .Q(n71) );
  MUX21X1 U573 ( .IN1(\mat_r[2][2][1] ), .IN2(\vector_in_r[2][1] ), .S(n450), 
        .Q(n72) );
  MUX21X1 U574 ( .IN1(\mat_r[2][2][2] ), .IN2(\vector_in_r[2][2] ), .S(n450), 
        .Q(n73) );
  MUX21X1 U575 ( .IN1(\mat_r[2][2][3] ), .IN2(\vector_in_r[2][3] ), .S(n450), 
        .Q(n74) );
  MUX21X1 U576 ( .IN1(\mat_r[2][2][4] ), .IN2(\vector_in_r[2][4] ), .S(n450), 
        .Q(n75) );
  MUX21X1 U577 ( .IN1(\mat_r[2][2][5] ), .IN2(\vector_in_r[2][5] ), .S(n450), 
        .Q(n76) );
  MUX21X1 U578 ( .IN1(\mat_r[2][2][6] ), .IN2(\vector_in_r[2][6] ), .S(n450), 
        .Q(n77) );
  MUX21X1 U579 ( .IN1(\mat_r[2][2][7] ), .IN2(\vector_in_r[2][7] ), .S(n450), 
        .Q(n78) );
  MUX21X1 U580 ( .IN1(\mat_r[2][2][8] ), .IN2(\vector_in_r[2][8] ), .S(n450), 
        .Q(n79) );
  MUX21X1 U581 ( .IN1(\mat_r[2][2][9] ), .IN2(\vector_in_r[2][9] ), .S(n450), 
        .Q(n80) );
  MUX21X1 U582 ( .IN1(\mat_r[2][2][10] ), .IN2(\vector_in_r[2][10] ), .S(n450), 
        .Q(n81) );
  MUX21X1 U583 ( .IN1(\mat_r[2][2][11] ), .IN2(\vector_in_r[2][11] ), .S(n450), 
        .Q(n82) );
  MUX21X1 U584 ( .IN1(\mat_r[2][1][0] ), .IN2(\vector_in_r[1][0] ), .S(n451), 
        .Q(n83) );
  MUX21X1 U585 ( .IN1(\mat_r[2][1][1] ), .IN2(\vector_in_r[1][1] ), .S(n451), 
        .Q(n84) );
  MUX21X1 U586 ( .IN1(\mat_r[2][1][2] ), .IN2(\vector_in_r[1][2] ), .S(n451), 
        .Q(n85) );
  MUX21X1 U587 ( .IN1(\mat_r[2][1][3] ), .IN2(\vector_in_r[1][3] ), .S(n451), 
        .Q(n86) );
  MUX21X1 U588 ( .IN1(\mat_r[2][1][4] ), .IN2(\vector_in_r[1][4] ), .S(n451), 
        .Q(n87) );
  MUX21X1 U589 ( .IN1(\mat_r[2][1][5] ), .IN2(\vector_in_r[1][5] ), .S(n451), 
        .Q(n88) );
  MUX21X1 U590 ( .IN1(\mat_r[2][1][6] ), .IN2(\vector_in_r[1][6] ), .S(n451), 
        .Q(n89) );
  MUX21X1 U591 ( .IN1(\mat_r[2][1][7] ), .IN2(\vector_in_r[1][7] ), .S(n451), 
        .Q(n90) );
  MUX21X1 U592 ( .IN1(\mat_r[2][1][8] ), .IN2(\vector_in_r[1][8] ), .S(n451), 
        .Q(n91) );
  MUX21X1 U593 ( .IN1(\mat_r[2][1][9] ), .IN2(\vector_in_r[1][9] ), .S(n451), 
        .Q(n92) );
  MUX21X1 U594 ( .IN1(\mat_r[2][1][10] ), .IN2(\vector_in_r[1][10] ), .S(n451), 
        .Q(n93) );
  MUX21X1 U595 ( .IN1(\mat_r[2][1][11] ), .IN2(\vector_in_r[1][11] ), .S(n451), 
        .Q(n94) );
  MUX21X1 U596 ( .IN1(\mat_r[2][0][0] ), .IN2(\vector_in_r[0][0] ), .S(n452), 
        .Q(n95) );
  MUX21X1 U597 ( .IN1(\mat_r[2][0][1] ), .IN2(\vector_in_r[0][1] ), .S(n452), 
        .Q(n96) );
  MUX21X1 U598 ( .IN1(\mat_r[2][0][2] ), .IN2(\vector_in_r[0][2] ), .S(n452), 
        .Q(n97) );
  MUX21X1 U599 ( .IN1(\mat_r[2][0][3] ), .IN2(\vector_in_r[0][3] ), .S(n452), 
        .Q(n98) );
  MUX21X1 U600 ( .IN1(\mat_r[2][0][4] ), .IN2(\vector_in_r[0][4] ), .S(n452), 
        .Q(n99) );
  MUX21X1 U601 ( .IN1(\mat_r[2][0][5] ), .IN2(\vector_in_r[0][5] ), .S(n452), 
        .Q(n100) );
  MUX21X1 U602 ( .IN1(\mat_r[2][0][6] ), .IN2(\vector_in_r[0][6] ), .S(n452), 
        .Q(n101) );
  MUX21X1 U603 ( .IN1(\mat_r[2][0][7] ), .IN2(\vector_in_r[0][7] ), .S(n452), 
        .Q(n102) );
  MUX21X1 U604 ( .IN1(\mat_r[2][0][8] ), .IN2(\vector_in_r[0][8] ), .S(n452), 
        .Q(n103) );
  MUX21X1 U605 ( .IN1(\mat_r[2][0][9] ), .IN2(\vector_in_r[0][9] ), .S(n452), 
        .Q(n104) );
  MUX21X1 U606 ( .IN1(\mat_r[2][0][10] ), .IN2(\vector_in_r[0][10] ), .S(n452), 
        .Q(n105) );
  MUX21X1 U607 ( .IN1(\mat_r[2][0][11] ), .IN2(\vector_in_r[0][11] ), .S(n452), 
        .Q(n106) );
  MUX21X1 U608 ( .IN1(\mat_i[3][3][0] ), .IN2(\vector_in_i[3][0] ), .S(n453), 
        .Q(n203) );
  MUX21X1 U609 ( .IN1(\mat_i[3][3][1] ), .IN2(\vector_in_i[3][1] ), .S(n453), 
        .Q(n204) );
  MUX21X1 U610 ( .IN1(\mat_i[3][3][2] ), .IN2(\vector_in_i[3][2] ), .S(n453), 
        .Q(n205) );
  MUX21X1 U611 ( .IN1(\mat_i[3][3][3] ), .IN2(\vector_in_i[3][3] ), .S(n453), 
        .Q(n206) );
  MUX21X1 U612 ( .IN1(\mat_i[3][3][4] ), .IN2(\vector_in_i[3][4] ), .S(n453), 
        .Q(n207) );
  MUX21X1 U613 ( .IN1(\mat_i[3][3][5] ), .IN2(\vector_in_i[3][5] ), .S(n453), 
        .Q(n208) );
  MUX21X1 U614 ( .IN1(\mat_i[3][3][6] ), .IN2(\vector_in_i[3][6] ), .S(n453), 
        .Q(n209) );
  MUX21X1 U615 ( .IN1(\mat_i[3][3][7] ), .IN2(\vector_in_i[3][7] ), .S(n453), 
        .Q(n210) );
  MUX21X1 U616 ( .IN1(\mat_i[3][3][8] ), .IN2(\vector_in_i[3][8] ), .S(n453), 
        .Q(n211) );
  MUX21X1 U617 ( .IN1(\mat_i[3][3][9] ), .IN2(\vector_in_i[3][9] ), .S(n453), 
        .Q(n212) );
  MUX21X1 U618 ( .IN1(\mat_i[3][3][10] ), .IN2(\vector_in_i[3][10] ), .S(n453), 
        .Q(n213) );
  MUX21X1 U619 ( .IN1(\mat_i[3][3][11] ), .IN2(\vector_in_i[3][11] ), .S(n453), 
        .Q(n214) );
  MUX21X1 U620 ( .IN1(\mat_i[3][2][0] ), .IN2(\vector_in_i[2][0] ), .S(n454), 
        .Q(n215) );
  MUX21X1 U621 ( .IN1(\mat_i[3][2][1] ), .IN2(\vector_in_i[2][1] ), .S(n454), 
        .Q(n216) );
  MUX21X1 U622 ( .IN1(\mat_i[3][2][2] ), .IN2(\vector_in_i[2][2] ), .S(n454), 
        .Q(n217) );
  MUX21X1 U623 ( .IN1(\mat_i[3][2][3] ), .IN2(\vector_in_i[2][3] ), .S(n454), 
        .Q(n218) );
  MUX21X1 U624 ( .IN1(\mat_i[3][2][4] ), .IN2(\vector_in_i[2][4] ), .S(n454), 
        .Q(n219) );
  MUX21X1 U625 ( .IN1(\mat_i[3][2][5] ), .IN2(\vector_in_i[2][5] ), .S(n454), 
        .Q(n220) );
  MUX21X1 U626 ( .IN1(\mat_i[3][2][6] ), .IN2(\vector_in_i[2][6] ), .S(n454), 
        .Q(n221) );
  MUX21X1 U627 ( .IN1(\mat_i[3][2][7] ), .IN2(\vector_in_i[2][7] ), .S(n454), 
        .Q(n222) );
  MUX21X1 U628 ( .IN1(\mat_i[3][2][8] ), .IN2(\vector_in_i[2][8] ), .S(n454), 
        .Q(n223) );
  MUX21X1 U629 ( .IN1(\mat_i[3][2][9] ), .IN2(\vector_in_i[2][9] ), .S(n454), 
        .Q(n224) );
  MUX21X1 U630 ( .IN1(\mat_i[3][2][10] ), .IN2(\vector_in_i[2][10] ), .S(n454), 
        .Q(n225) );
  MUX21X1 U631 ( .IN1(\mat_i[3][2][11] ), .IN2(\vector_in_i[2][11] ), .S(n454), 
        .Q(n226) );
  MUX21X1 U632 ( .IN1(\mat_i[3][1][0] ), .IN2(\vector_in_i[1][0] ), .S(n455), 
        .Q(n227) );
  MUX21X1 U633 ( .IN1(\mat_i[3][1][1] ), .IN2(\vector_in_i[1][1] ), .S(n455), 
        .Q(n228) );
  MUX21X1 U634 ( .IN1(\mat_i[3][1][2] ), .IN2(\vector_in_i[1][2] ), .S(n455), 
        .Q(n229) );
  MUX21X1 U635 ( .IN1(\mat_i[3][1][3] ), .IN2(\vector_in_i[1][3] ), .S(n455), 
        .Q(n230) );
  MUX21X1 U636 ( .IN1(\mat_i[3][1][4] ), .IN2(\vector_in_i[1][4] ), .S(n455), 
        .Q(n231) );
  MUX21X1 U637 ( .IN1(\mat_i[3][1][5] ), .IN2(\vector_in_i[1][5] ), .S(n455), 
        .Q(n232) );
  MUX21X1 U638 ( .IN1(\mat_i[3][1][6] ), .IN2(\vector_in_i[1][6] ), .S(n455), 
        .Q(n233) );
  MUX21X1 U639 ( .IN1(\mat_i[3][1][7] ), .IN2(\vector_in_i[1][7] ), .S(n455), 
        .Q(n234) );
  MUX21X1 U640 ( .IN1(\mat_i[3][1][8] ), .IN2(\vector_in_i[1][8] ), .S(n455), 
        .Q(n235) );
  MUX21X1 U641 ( .IN1(\mat_i[3][1][9] ), .IN2(\vector_in_i[1][9] ), .S(n455), 
        .Q(n236) );
  MUX21X1 U642 ( .IN1(\mat_i[3][1][10] ), .IN2(\vector_in_i[1][10] ), .S(n455), 
        .Q(n237) );
  MUX21X1 U643 ( .IN1(\mat_i[3][1][11] ), .IN2(\vector_in_i[1][11] ), .S(n455), 
        .Q(n238) );
  MUX21X1 U644 ( .IN1(\mat_i[3][0][0] ), .IN2(\vector_in_i[0][0] ), .S(n456), 
        .Q(n239) );
  MUX21X1 U645 ( .IN1(\mat_i[3][0][1] ), .IN2(\vector_in_i[0][1] ), .S(n456), 
        .Q(n240) );
  MUX21X1 U646 ( .IN1(\mat_i[3][0][2] ), .IN2(\vector_in_i[0][2] ), .S(n456), 
        .Q(n241) );
  MUX21X1 U647 ( .IN1(\mat_i[3][0][3] ), .IN2(\vector_in_i[0][3] ), .S(n456), 
        .Q(n242) );
  MUX21X1 U648 ( .IN1(\mat_i[3][0][4] ), .IN2(\vector_in_i[0][4] ), .S(n456), 
        .Q(n243) );
  MUX21X1 U649 ( .IN1(\mat_i[3][0][5] ), .IN2(\vector_in_i[0][5] ), .S(n456), 
        .Q(n244) );
  MUX21X1 U650 ( .IN1(\mat_i[3][0][6] ), .IN2(\vector_in_i[0][6] ), .S(n456), 
        .Q(n245) );
  MUX21X1 U651 ( .IN1(\mat_i[3][0][7] ), .IN2(\vector_in_i[0][7] ), .S(n456), 
        .Q(n246) );
  MUX21X1 U652 ( .IN1(\mat_i[3][0][8] ), .IN2(\vector_in_i[0][8] ), .S(n456), 
        .Q(n247) );
  MUX21X1 U653 ( .IN1(\mat_i[3][0][9] ), .IN2(\vector_in_i[0][9] ), .S(n456), 
        .Q(n248) );
  MUX21X1 U654 ( .IN1(\mat_i[3][0][10] ), .IN2(\vector_in_i[0][10] ), .S(n456), 
        .Q(n249) );
  MUX21X1 U655 ( .IN1(\mat_i[3][0][11] ), .IN2(\vector_in_i[0][11] ), .S(n456), 
        .Q(n250) );
  MUX21X1 U656 ( .IN1(\mat_r[3][3][0] ), .IN2(\vector_in_r[3][0] ), .S(n457), 
        .Q(n11) );
  MUX21X1 U657 ( .IN1(\mat_r[3][3][1] ), .IN2(\vector_in_r[3][1] ), .S(n457), 
        .Q(n12) );
  MUX21X1 U658 ( .IN1(\mat_r[3][3][2] ), .IN2(\vector_in_r[3][2] ), .S(n457), 
        .Q(n13) );
  MUX21X1 U659 ( .IN1(\mat_r[3][3][3] ), .IN2(\vector_in_r[3][3] ), .S(n457), 
        .Q(n14) );
  MUX21X1 U660 ( .IN1(\mat_r[3][3][4] ), .IN2(\vector_in_r[3][4] ), .S(n457), 
        .Q(n15) );
  MUX21X1 U661 ( .IN1(\mat_r[3][3][5] ), .IN2(\vector_in_r[3][5] ), .S(n457), 
        .Q(n16) );
  MUX21X1 U662 ( .IN1(\mat_r[3][3][6] ), .IN2(\vector_in_r[3][6] ), .S(n457), 
        .Q(n17) );
  MUX21X1 U663 ( .IN1(\mat_r[3][3][7] ), .IN2(\vector_in_r[3][7] ), .S(n457), 
        .Q(n18) );
  MUX21X1 U664 ( .IN1(\mat_r[3][3][8] ), .IN2(\vector_in_r[3][8] ), .S(n457), 
        .Q(n19) );
  MUX21X1 U665 ( .IN1(\mat_r[3][3][9] ), .IN2(\vector_in_r[3][9] ), .S(n457), 
        .Q(n20) );
  MUX21X1 U666 ( .IN1(\mat_r[3][3][10] ), .IN2(\vector_in_r[3][10] ), .S(n457), 
        .Q(n21) );
  MUX21X1 U667 ( .IN1(\mat_r[3][3][11] ), .IN2(\vector_in_r[3][11] ), .S(n457), 
        .Q(n22) );
  MUX21X1 U668 ( .IN1(\mat_r[3][2][0] ), .IN2(\vector_in_r[2][0] ), .S(n458), 
        .Q(n23) );
  MUX21X1 U669 ( .IN1(\mat_r[3][2][1] ), .IN2(\vector_in_r[2][1] ), .S(n458), 
        .Q(n24) );
  MUX21X1 U670 ( .IN1(\mat_r[3][2][2] ), .IN2(\vector_in_r[2][2] ), .S(n458), 
        .Q(n25) );
  MUX21X1 U671 ( .IN1(\mat_r[3][2][3] ), .IN2(\vector_in_r[2][3] ), .S(n458), 
        .Q(n26) );
  MUX21X1 U672 ( .IN1(\mat_r[3][2][4] ), .IN2(\vector_in_r[2][4] ), .S(n458), 
        .Q(n27) );
  MUX21X1 U673 ( .IN1(\mat_r[3][2][5] ), .IN2(\vector_in_r[2][5] ), .S(n458), 
        .Q(n28) );
  MUX21X1 U674 ( .IN1(\mat_r[3][2][6] ), .IN2(\vector_in_r[2][6] ), .S(n458), 
        .Q(n29) );
  MUX21X1 U675 ( .IN1(\mat_r[3][2][7] ), .IN2(\vector_in_r[2][7] ), .S(n458), 
        .Q(n30) );
  MUX21X1 U676 ( .IN1(\mat_r[3][2][8] ), .IN2(\vector_in_r[2][8] ), .S(n458), 
        .Q(n31) );
  MUX21X1 U677 ( .IN1(\mat_r[3][2][9] ), .IN2(\vector_in_r[2][9] ), .S(n458), 
        .Q(n32) );
  MUX21X1 U678 ( .IN1(\mat_r[3][2][10] ), .IN2(\vector_in_r[2][10] ), .S(n458), 
        .Q(n33) );
  MUX21X1 U679 ( .IN1(\mat_r[3][2][11] ), .IN2(\vector_in_r[2][11] ), .S(n458), 
        .Q(n34) );
  MUX21X1 U680 ( .IN1(\mat_r[3][1][0] ), .IN2(\vector_in_r[1][0] ), .S(n459), 
        .Q(n35) );
  MUX21X1 U681 ( .IN1(\mat_r[3][1][1] ), .IN2(\vector_in_r[1][1] ), .S(n459), 
        .Q(n36) );
  MUX21X1 U682 ( .IN1(\mat_r[3][1][2] ), .IN2(\vector_in_r[1][2] ), .S(n459), 
        .Q(n37) );
  MUX21X1 U683 ( .IN1(\mat_r[3][1][3] ), .IN2(\vector_in_r[1][3] ), .S(n459), 
        .Q(n38) );
  MUX21X1 U684 ( .IN1(\mat_r[3][1][4] ), .IN2(\vector_in_r[1][4] ), .S(n459), 
        .Q(n39) );
  MUX21X1 U685 ( .IN1(\mat_r[3][1][5] ), .IN2(\vector_in_r[1][5] ), .S(n459), 
        .Q(n40) );
  MUX21X1 U686 ( .IN1(\mat_r[3][1][6] ), .IN2(\vector_in_r[1][6] ), .S(n459), 
        .Q(n41) );
  MUX21X1 U687 ( .IN1(\mat_r[3][1][7] ), .IN2(\vector_in_r[1][7] ), .S(n459), 
        .Q(n42) );
  MUX21X1 U688 ( .IN1(\mat_r[3][1][8] ), .IN2(\vector_in_r[1][8] ), .S(n459), 
        .Q(n43) );
  MUX21X1 U689 ( .IN1(\mat_r[3][1][9] ), .IN2(\vector_in_r[1][9] ), .S(n459), 
        .Q(n44) );
  MUX21X1 U690 ( .IN1(\mat_r[3][1][10] ), .IN2(\vector_in_r[1][10] ), .S(n459), 
        .Q(n45) );
  MUX21X1 U691 ( .IN1(\mat_r[3][1][11] ), .IN2(\vector_in_r[1][11] ), .S(n459), 
        .Q(n46) );
  MUX21X1 U692 ( .IN1(\mat_r[3][0][0] ), .IN2(\vector_in_r[0][0] ), .S(n460), 
        .Q(n47) );
  MUX21X1 U693 ( .IN1(\mat_r[3][0][1] ), .IN2(\vector_in_r[0][1] ), .S(n460), 
        .Q(n48) );
  MUX21X1 U694 ( .IN1(\mat_r[3][0][2] ), .IN2(\vector_in_r[0][2] ), .S(n460), 
        .Q(n49) );
  MUX21X1 U695 ( .IN1(\mat_r[3][0][3] ), .IN2(\vector_in_r[0][3] ), .S(n460), 
        .Q(n50) );
  MUX21X1 U696 ( .IN1(\mat_r[3][0][4] ), .IN2(\vector_in_r[0][4] ), .S(n460), 
        .Q(n51) );
  MUX21X1 U697 ( .IN1(\mat_r[3][0][5] ), .IN2(\vector_in_r[0][5] ), .S(n460), 
        .Q(n52) );
  MUX21X1 U698 ( .IN1(\mat_r[3][0][6] ), .IN2(\vector_in_r[0][6] ), .S(n460), 
        .Q(n53) );
  MUX21X1 U699 ( .IN1(\mat_r[3][0][7] ), .IN2(\vector_in_r[0][7] ), .S(n460), 
        .Q(n54) );
  MUX21X1 U700 ( .IN1(\mat_r[3][0][8] ), .IN2(\vector_in_r[0][8] ), .S(n460), 
        .Q(n55) );
  MUX21X1 U701 ( .IN1(\mat_r[3][0][9] ), .IN2(\vector_in_r[0][9] ), .S(n460), 
        .Q(n56) );
  MUX21X1 U702 ( .IN1(\mat_r[3][0][10] ), .IN2(\vector_in_r[0][10] ), .S(n460), 
        .Q(n57) );
  MUX21X1 U703 ( .IN1(\mat_r[3][0][11] ), .IN2(\vector_in_r[0][11] ), .S(n460), 
        .Q(n58) );
endmodule


module r_mat_regs_WORD_WIDTH12_N4_LOG2_N2 ( single_in_r, single_in_i, 
    .vector_out_r({\vector_out_r[0][11] , \vector_out_r[0][10] , 
        \vector_out_r[0][9] , \vector_out_r[0][8] , \vector_out_r[0][7] , 
        \vector_out_r[0][6] , \vector_out_r[0][5] , \vector_out_r[0][4] , 
        \vector_out_r[0][3] , \vector_out_r[0][2] , \vector_out_r[0][1] , 
        \vector_out_r[0][0] , \vector_out_r[1][11] , \vector_out_r[1][10] , 
        \vector_out_r[1][9] , \vector_out_r[1][8] , \vector_out_r[1][7] , 
        \vector_out_r[1][6] , \vector_out_r[1][5] , \vector_out_r[1][4] , 
        \vector_out_r[1][3] , \vector_out_r[1][2] , \vector_out_r[1][1] , 
        \vector_out_r[1][0] , \vector_out_r[2][11] , \vector_out_r[2][10] , 
        \vector_out_r[2][9] , \vector_out_r[2][8] , \vector_out_r[2][7] , 
        \vector_out_r[2][6] , \vector_out_r[2][5] , \vector_out_r[2][4] , 
        \vector_out_r[2][3] , \vector_out_r[2][2] , \vector_out_r[2][1] , 
        \vector_out_r[2][0] , \vector_out_r[3][11] , \vector_out_r[3][10] , 
        \vector_out_r[3][9] , \vector_out_r[3][8] , \vector_out_r[3][7] , 
        \vector_out_r[3][6] , \vector_out_r[3][5] , \vector_out_r[3][4] , 
        \vector_out_r[3][3] , \vector_out_r[3][2] , \vector_out_r[3][1] , 
        \vector_out_r[3][0] }), .vector_out_i({\vector_out_i[0][11] , 
        \vector_out_i[0][10] , \vector_out_i[0][9] , \vector_out_i[0][8] , 
        \vector_out_i[0][7] , \vector_out_i[0][6] , \vector_out_i[0][5] , 
        \vector_out_i[0][4] , \vector_out_i[0][3] , \vector_out_i[0][2] , 
        \vector_out_i[0][1] , \vector_out_i[0][0] , \vector_out_i[1][11] , 
        \vector_out_i[1][10] , \vector_out_i[1][9] , \vector_out_i[1][8] , 
        \vector_out_i[1][7] , \vector_out_i[1][6] , \vector_out_i[1][5] , 
        \vector_out_i[1][4] , \vector_out_i[1][3] , \vector_out_i[1][2] , 
        \vector_out_i[1][1] , \vector_out_i[1][0] , \vector_out_i[2][11] , 
        \vector_out_i[2][10] , \vector_out_i[2][9] , \vector_out_i[2][8] , 
        \vector_out_i[2][7] , \vector_out_i[2][6] , \vector_out_i[2][5] , 
        \vector_out_i[2][4] , \vector_out_i[2][3] , \vector_out_i[2][2] , 
        \vector_out_i[2][1] , \vector_out_i[2][0] , \vector_out_i[3][11] , 
        \vector_out_i[3][10] , \vector_out_i[3][9] , \vector_out_i[3][8] , 
        \vector_out_i[3][7] , \vector_out_i[3][6] , \vector_out_i[3][5] , 
        \vector_out_i[3][4] , \vector_out_i[3][3] , \vector_out_i[3][2] , 
        \vector_out_i[3][1] , \vector_out_i[3][0] }), col_sel, row_sel, clk, 
        wr_enable );
  input [11:0] single_in_r;
  input [11:0] single_in_i;
  input [1:0] col_sel;
  input [1:0] row_sel;
  input clk, wr_enable;
  output \vector_out_r[0][11] , \vector_out_r[0][10] , \vector_out_r[0][9] ,
         \vector_out_r[0][8] , \vector_out_r[0][7] , \vector_out_r[0][6] ,
         \vector_out_r[0][5] , \vector_out_r[0][4] , \vector_out_r[0][3] ,
         \vector_out_r[0][2] , \vector_out_r[0][1] , \vector_out_r[0][0] ,
         \vector_out_r[1][11] , \vector_out_r[1][10] , \vector_out_r[1][9] ,
         \vector_out_r[1][8] , \vector_out_r[1][7] , \vector_out_r[1][6] ,
         \vector_out_r[1][5] , \vector_out_r[1][4] , \vector_out_r[1][3] ,
         \vector_out_r[1][2] , \vector_out_r[1][1] , \vector_out_r[1][0] ,
         \vector_out_r[2][11] , \vector_out_r[2][10] , \vector_out_r[2][9] ,
         \vector_out_r[2][8] , \vector_out_r[2][7] , \vector_out_r[2][6] ,
         \vector_out_r[2][5] , \vector_out_r[2][4] , \vector_out_r[2][3] ,
         \vector_out_r[2][2] , \vector_out_r[2][1] , \vector_out_r[2][0] ,
         \vector_out_r[3][11] , \vector_out_r[3][10] , \vector_out_r[3][9] ,
         \vector_out_r[3][8] , \vector_out_r[3][7] , \vector_out_r[3][6] ,
         \vector_out_r[3][5] , \vector_out_r[3][4] , \vector_out_r[3][3] ,
         \vector_out_r[3][2] , \vector_out_r[3][1] , \vector_out_r[3][0] ,
         \vector_out_i[0][11] , \vector_out_i[0][10] , \vector_out_i[0][9] ,
         \vector_out_i[0][8] , \vector_out_i[0][7] , \vector_out_i[0][6] ,
         \vector_out_i[0][5] , \vector_out_i[0][4] , \vector_out_i[0][3] ,
         \vector_out_i[0][2] , \vector_out_i[0][1] , \vector_out_i[0][0] ,
         \vector_out_i[1][11] , \vector_out_i[1][10] , \vector_out_i[1][9] ,
         \vector_out_i[1][8] , \vector_out_i[1][7] , \vector_out_i[1][6] ,
         \vector_out_i[1][5] , \vector_out_i[1][4] , \vector_out_i[1][3] ,
         \vector_out_i[1][2] , \vector_out_i[1][1] , \vector_out_i[1][0] ,
         \vector_out_i[2][11] , \vector_out_i[2][10] , \vector_out_i[2][9] ,
         \vector_out_i[2][8] , \vector_out_i[2][7] , \vector_out_i[2][6] ,
         \vector_out_i[2][5] , \vector_out_i[2][4] , \vector_out_i[2][3] ,
         \vector_out_i[2][2] , \vector_out_i[2][1] , \vector_out_i[2][0] ,
         \vector_out_i[3][11] , \vector_out_i[3][10] , \vector_out_i[3][9] ,
         \vector_out_i[3][8] , \vector_out_i[3][7] , \vector_out_i[3][6] ,
         \vector_out_i[3][5] , \vector_out_i[3][4] , \vector_out_i[3][3] ,
         \vector_out_i[3][2] , \vector_out_i[3][1] , \vector_out_i[3][0] ;
  wire   N11, N12, \mat_r[0][0][11] , \mat_r[0][0][10] , \mat_r[0][0][9] ,
         \mat_r[0][0][8] , \mat_r[0][0][7] , \mat_r[0][0][6] ,
         \mat_r[0][0][5] , \mat_r[0][0][4] , \mat_r[0][0][3] ,
         \mat_r[0][0][2] , \mat_r[0][0][1] , \mat_r[0][0][0] ,
         \mat_r[1][0][11] , \mat_r[1][0][10] , \mat_r[1][0][9] ,
         \mat_r[1][0][8] , \mat_r[1][0][7] , \mat_r[1][0][6] ,
         \mat_r[1][0][5] , \mat_r[1][0][4] , \mat_r[1][0][3] ,
         \mat_r[1][0][2] , \mat_r[1][0][1] , \mat_r[1][0][0] ,
         \mat_r[1][1][11] , \mat_r[1][1][10] , \mat_r[1][1][9] ,
         \mat_r[1][1][8] , \mat_r[1][1][7] , \mat_r[1][1][6] ,
         \mat_r[1][1][5] , \mat_r[1][1][4] , \mat_r[1][1][3] ,
         \mat_r[1][1][2] , \mat_r[1][1][1] , \mat_r[1][1][0] ,
         \mat_r[2][0][11] , \mat_r[2][0][10] , \mat_r[2][0][9] ,
         \mat_r[2][0][8] , \mat_r[2][0][7] , \mat_r[2][0][6] ,
         \mat_r[2][0][5] , \mat_r[2][0][4] , \mat_r[2][0][3] ,
         \mat_r[2][0][2] , \mat_r[2][0][1] , \mat_r[2][0][0] ,
         \mat_r[2][1][11] , \mat_r[2][1][10] , \mat_r[2][1][9] ,
         \mat_r[2][1][8] , \mat_r[2][1][7] , \mat_r[2][1][6] ,
         \mat_r[2][1][5] , \mat_r[2][1][4] , \mat_r[2][1][3] ,
         \mat_r[2][1][2] , \mat_r[2][1][1] , \mat_r[2][1][0] ,
         \mat_r[2][2][11] , \mat_r[2][2][10] , \mat_r[2][2][9] ,
         \mat_r[2][2][8] , \mat_r[2][2][7] , \mat_r[2][2][6] ,
         \mat_r[2][2][5] , \mat_r[2][2][4] , \mat_r[2][2][3] ,
         \mat_r[2][2][2] , \mat_r[2][2][1] , \mat_r[2][2][0] ,
         \mat_r[3][0][11] , \mat_r[3][0][10] , \mat_r[3][0][9] ,
         \mat_r[3][0][8] , \mat_r[3][0][7] , \mat_r[3][0][6] ,
         \mat_r[3][0][5] , \mat_r[3][0][4] , \mat_r[3][0][3] ,
         \mat_r[3][0][2] , \mat_r[3][0][1] , \mat_r[3][0][0] ,
         \mat_r[3][1][11] , \mat_r[3][1][10] , \mat_r[3][1][9] ,
         \mat_r[3][1][8] , \mat_r[3][1][7] , \mat_r[3][1][6] ,
         \mat_r[3][1][5] , \mat_r[3][1][4] , \mat_r[3][1][3] ,
         \mat_r[3][1][2] , \mat_r[3][1][1] , \mat_r[3][1][0] ,
         \mat_r[3][2][11] , \mat_r[3][2][10] , \mat_r[3][2][9] ,
         \mat_r[3][2][8] , \mat_r[3][2][7] , \mat_r[3][2][6] ,
         \mat_r[3][2][5] , \mat_r[3][2][4] , \mat_r[3][2][3] ,
         \mat_r[3][2][2] , \mat_r[3][2][1] , \mat_r[3][2][0] ,
         \mat_r[3][3][11] , \mat_r[3][3][10] , \mat_r[3][3][9] ,
         \mat_r[3][3][8] , \mat_r[3][3][7] , \mat_r[3][3][6] ,
         \mat_r[3][3][5] , \mat_r[3][3][4] , \mat_r[3][3][3] ,
         \mat_r[3][3][2] , \mat_r[3][3][1] , \mat_r[3][3][0] ,
         \mat_i[1][0][11] , \mat_i[1][0][10] , \mat_i[1][0][9] ,
         \mat_i[1][0][8] , \mat_i[1][0][7] , \mat_i[1][0][6] ,
         \mat_i[1][0][5] , \mat_i[1][0][4] , \mat_i[1][0][3] ,
         \mat_i[1][0][2] , \mat_i[1][0][1] , \mat_i[1][0][0] ,
         \mat_i[2][0][11] , \mat_i[2][0][10] , \mat_i[2][0][9] ,
         \mat_i[2][0][8] , \mat_i[2][0][7] , \mat_i[2][0][6] ,
         \mat_i[2][0][5] , \mat_i[2][0][4] , \mat_i[2][0][3] ,
         \mat_i[2][0][2] , \mat_i[2][0][1] , \mat_i[2][0][0] ,
         \mat_i[2][1][11] , \mat_i[2][1][10] , \mat_i[2][1][9] ,
         \mat_i[2][1][8] , \mat_i[2][1][7] , \mat_i[2][1][6] ,
         \mat_i[2][1][5] , \mat_i[2][1][4] , \mat_i[2][1][3] ,
         \mat_i[2][1][2] , \mat_i[2][1][1] , \mat_i[2][1][0] ,
         \mat_i[3][0][11] , \mat_i[3][0][10] , \mat_i[3][0][9] ,
         \mat_i[3][0][8] , \mat_i[3][0][7] , \mat_i[3][0][6] ,
         \mat_i[3][0][5] , \mat_i[3][0][4] , \mat_i[3][0][3] ,
         \mat_i[3][0][2] , \mat_i[3][0][1] , \mat_i[3][0][0] ,
         \mat_i[3][1][11] , \mat_i[3][1][10] , \mat_i[3][1][9] ,
         \mat_i[3][1][8] , \mat_i[3][1][7] , \mat_i[3][1][6] ,
         \mat_i[3][1][5] , \mat_i[3][1][4] , \mat_i[3][1][3] ,
         \mat_i[3][1][2] , \mat_i[3][1][1] , \mat_i[3][1][0] ,
         \mat_i[3][2][11] , \mat_i[3][2][10] , \mat_i[3][2][9] ,
         \mat_i[3][2][8] , \mat_i[3][2][7] , \mat_i[3][2][6] ,
         \mat_i[3][2][5] , \mat_i[3][2][4] , \mat_i[3][2][3] ,
         \mat_i[3][2][2] , \mat_i[3][2][1] , \mat_i[3][2][0] , n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330;
  assign N11 = col_sel[0];
  assign N12 = col_sel[1];
  assign \vector_out_i[3][0]  = 1'b0;
  assign \vector_out_i[3][1]  = 1'b0;
  assign \vector_out_i[3][2]  = 1'b0;
  assign \vector_out_i[3][3]  = 1'b0;
  assign \vector_out_i[3][4]  = 1'b0;
  assign \vector_out_i[3][5]  = 1'b0;
  assign \vector_out_i[3][6]  = 1'b0;
  assign \vector_out_i[3][7]  = 1'b0;
  assign \vector_out_i[3][8]  = 1'b0;
  assign \vector_out_i[3][9]  = 1'b0;
  assign \vector_out_i[3][10]  = 1'b0;
  assign \vector_out_i[3][11]  = 1'b0;

  DFFX1 \mat_i_reg_reg[1][0][11]  ( .D(n224), .CLK(clk), .Q(\mat_i[1][0][11] )
         );
  DFFX1 \mat_i_reg_reg[1][0][10]  ( .D(n223), .CLK(clk), .Q(\mat_i[1][0][10] )
         );
  DFFX1 \mat_i_reg_reg[1][0][9]  ( .D(n222), .CLK(clk), .Q(\mat_i[1][0][9] )
         );
  DFFX1 \mat_i_reg_reg[1][0][8]  ( .D(n221), .CLK(clk), .Q(\mat_i[1][0][8] )
         );
  DFFX1 \mat_i_reg_reg[1][0][7]  ( .D(n220), .CLK(clk), .Q(\mat_i[1][0][7] )
         );
  DFFX1 \mat_i_reg_reg[1][0][6]  ( .D(n219), .CLK(clk), .Q(\mat_i[1][0][6] )
         );
  DFFX1 \mat_i_reg_reg[1][0][5]  ( .D(n218), .CLK(clk), .Q(\mat_i[1][0][5] )
         );
  DFFX1 \mat_i_reg_reg[1][0][4]  ( .D(n217), .CLK(clk), .Q(\mat_i[1][0][4] )
         );
  DFFX1 \mat_i_reg_reg[1][0][3]  ( .D(n216), .CLK(clk), .Q(\mat_i[1][0][3] )
         );
  DFFX1 \mat_i_reg_reg[1][0][2]  ( .D(n215), .CLK(clk), .Q(\mat_i[1][0][2] )
         );
  DFFX1 \mat_i_reg_reg[1][0][1]  ( .D(n214), .CLK(clk), .Q(\mat_i[1][0][1] )
         );
  DFFX1 \mat_i_reg_reg[1][0][0]  ( .D(n213), .CLK(clk), .Q(\mat_i[1][0][0] )
         );
  DFFX1 \mat_i_reg_reg[2][0][11]  ( .D(n212), .CLK(clk), .Q(\mat_i[2][0][11] )
         );
  DFFX1 \mat_i_reg_reg[2][0][10]  ( .D(n211), .CLK(clk), .Q(\mat_i[2][0][10] )
         );
  DFFX1 \mat_i_reg_reg[2][0][9]  ( .D(n210), .CLK(clk), .Q(\mat_i[2][0][9] )
         );
  DFFX1 \mat_i_reg_reg[2][0][8]  ( .D(n209), .CLK(clk), .Q(\mat_i[2][0][8] )
         );
  DFFX1 \mat_i_reg_reg[2][0][7]  ( .D(n208), .CLK(clk), .Q(\mat_i[2][0][7] )
         );
  DFFX1 \mat_i_reg_reg[2][0][6]  ( .D(n207), .CLK(clk), .Q(\mat_i[2][0][6] )
         );
  DFFX1 \mat_i_reg_reg[2][0][5]  ( .D(n206), .CLK(clk), .Q(\mat_i[2][0][5] )
         );
  DFFX1 \mat_i_reg_reg[2][0][4]  ( .D(n205), .CLK(clk), .Q(\mat_i[2][0][4] )
         );
  DFFX1 \mat_i_reg_reg[2][0][3]  ( .D(n204), .CLK(clk), .Q(\mat_i[2][0][3] )
         );
  DFFX1 \mat_i_reg_reg[2][0][2]  ( .D(n203), .CLK(clk), .Q(\mat_i[2][0][2] )
         );
  DFFX1 \mat_i_reg_reg[2][0][1]  ( .D(n202), .CLK(clk), .Q(\mat_i[2][0][1] )
         );
  DFFX1 \mat_i_reg_reg[2][0][0]  ( .D(n201), .CLK(clk), .Q(\mat_i[2][0][0] )
         );
  DFFX1 \mat_i_reg_reg[2][1][11]  ( .D(n200), .CLK(clk), .Q(\mat_i[2][1][11] )
         );
  DFFX1 \mat_i_reg_reg[2][1][10]  ( .D(n199), .CLK(clk), .Q(\mat_i[2][1][10] )
         );
  DFFX1 \mat_i_reg_reg[2][1][9]  ( .D(n198), .CLK(clk), .Q(\mat_i[2][1][9] )
         );
  DFFX1 \mat_i_reg_reg[2][1][8]  ( .D(n197), .CLK(clk), .Q(\mat_i[2][1][8] )
         );
  DFFX1 \mat_i_reg_reg[2][1][7]  ( .D(n196), .CLK(clk), .Q(\mat_i[2][1][7] )
         );
  DFFX1 \mat_i_reg_reg[2][1][6]  ( .D(n195), .CLK(clk), .Q(\mat_i[2][1][6] )
         );
  DFFX1 \mat_i_reg_reg[2][1][5]  ( .D(n194), .CLK(clk), .Q(\mat_i[2][1][5] )
         );
  DFFX1 \mat_i_reg_reg[2][1][4]  ( .D(n193), .CLK(clk), .Q(\mat_i[2][1][4] )
         );
  DFFX1 \mat_i_reg_reg[2][1][3]  ( .D(n192), .CLK(clk), .Q(\mat_i[2][1][3] )
         );
  DFFX1 \mat_i_reg_reg[2][1][2]  ( .D(n191), .CLK(clk), .Q(\mat_i[2][1][2] )
         );
  DFFX1 \mat_i_reg_reg[2][1][1]  ( .D(n190), .CLK(clk), .Q(\mat_i[2][1][1] )
         );
  DFFX1 \mat_i_reg_reg[2][1][0]  ( .D(n189), .CLK(clk), .Q(\mat_i[2][1][0] )
         );
  DFFX1 \mat_i_reg_reg[3][0][11]  ( .D(n188), .CLK(clk), .Q(\mat_i[3][0][11] )
         );
  DFFX1 \mat_i_reg_reg[3][0][10]  ( .D(n187), .CLK(clk), .Q(\mat_i[3][0][10] )
         );
  DFFX1 \mat_i_reg_reg[3][0][9]  ( .D(n186), .CLK(clk), .Q(\mat_i[3][0][9] )
         );
  DFFX1 \mat_i_reg_reg[3][0][8]  ( .D(n185), .CLK(clk), .Q(\mat_i[3][0][8] )
         );
  DFFX1 \mat_i_reg_reg[3][0][7]  ( .D(n184), .CLK(clk), .Q(\mat_i[3][0][7] )
         );
  DFFX1 \mat_i_reg_reg[3][0][6]  ( .D(n183), .CLK(clk), .Q(\mat_i[3][0][6] )
         );
  DFFX1 \mat_i_reg_reg[3][0][5]  ( .D(n182), .CLK(clk), .Q(\mat_i[3][0][5] )
         );
  DFFX1 \mat_i_reg_reg[3][0][4]  ( .D(n181), .CLK(clk), .Q(\mat_i[3][0][4] )
         );
  DFFX1 \mat_i_reg_reg[3][0][3]  ( .D(n180), .CLK(clk), .Q(\mat_i[3][0][3] )
         );
  DFFX1 \mat_i_reg_reg[3][0][2]  ( .D(n179), .CLK(clk), .Q(\mat_i[3][0][2] )
         );
  DFFX1 \mat_i_reg_reg[3][0][1]  ( .D(n178), .CLK(clk), .Q(\mat_i[3][0][1] )
         );
  DFFX1 \mat_i_reg_reg[3][0][0]  ( .D(n177), .CLK(clk), .Q(\mat_i[3][0][0] )
         );
  DFFX1 \mat_i_reg_reg[3][1][11]  ( .D(n176), .CLK(clk), .Q(\mat_i[3][1][11] )
         );
  DFFX1 \mat_i_reg_reg[3][1][10]  ( .D(n175), .CLK(clk), .Q(\mat_i[3][1][10] )
         );
  DFFX1 \mat_i_reg_reg[3][1][9]  ( .D(n174), .CLK(clk), .Q(\mat_i[3][1][9] )
         );
  DFFX1 \mat_i_reg_reg[3][1][8]  ( .D(n173), .CLK(clk), .Q(\mat_i[3][1][8] )
         );
  DFFX1 \mat_i_reg_reg[3][1][7]  ( .D(n172), .CLK(clk), .Q(\mat_i[3][1][7] )
         );
  DFFX1 \mat_i_reg_reg[3][1][6]  ( .D(n171), .CLK(clk), .Q(\mat_i[3][1][6] )
         );
  DFFX1 \mat_i_reg_reg[3][1][5]  ( .D(n170), .CLK(clk), .Q(\mat_i[3][1][5] )
         );
  DFFX1 \mat_i_reg_reg[3][1][4]  ( .D(n169), .CLK(clk), .Q(\mat_i[3][1][4] )
         );
  DFFX1 \mat_i_reg_reg[3][1][3]  ( .D(n168), .CLK(clk), .Q(\mat_i[3][1][3] )
         );
  DFFX1 \mat_i_reg_reg[3][1][2]  ( .D(n167), .CLK(clk), .Q(\mat_i[3][1][2] )
         );
  DFFX1 \mat_i_reg_reg[3][1][1]  ( .D(n166), .CLK(clk), .Q(\mat_i[3][1][1] )
         );
  DFFX1 \mat_i_reg_reg[3][1][0]  ( .D(n165), .CLK(clk), .Q(\mat_i[3][1][0] )
         );
  DFFX1 \mat_i_reg_reg[3][2][11]  ( .D(n164), .CLK(clk), .Q(\mat_i[3][2][11] )
         );
  DFFX1 \mat_i_reg_reg[3][2][10]  ( .D(n163), .CLK(clk), .Q(\mat_i[3][2][10] )
         );
  DFFX1 \mat_i_reg_reg[3][2][9]  ( .D(n162), .CLK(clk), .Q(\mat_i[3][2][9] )
         );
  DFFX1 \mat_i_reg_reg[3][2][8]  ( .D(n161), .CLK(clk), .Q(\mat_i[3][2][8] )
         );
  DFFX1 \mat_i_reg_reg[3][2][7]  ( .D(n160), .CLK(clk), .Q(\mat_i[3][2][7] )
         );
  DFFX1 \mat_i_reg_reg[3][2][6]  ( .D(n159), .CLK(clk), .Q(\mat_i[3][2][6] )
         );
  DFFX1 \mat_i_reg_reg[3][2][5]  ( .D(n158), .CLK(clk), .Q(\mat_i[3][2][5] )
         );
  DFFX1 \mat_i_reg_reg[3][2][4]  ( .D(n157), .CLK(clk), .Q(\mat_i[3][2][4] )
         );
  DFFX1 \mat_i_reg_reg[3][2][3]  ( .D(n156), .CLK(clk), .Q(\mat_i[3][2][3] )
         );
  DFFX1 \mat_i_reg_reg[3][2][2]  ( .D(n155), .CLK(clk), .Q(\mat_i[3][2][2] )
         );
  DFFX1 \mat_i_reg_reg[3][2][1]  ( .D(n154), .CLK(clk), .Q(\mat_i[3][2][1] )
         );
  DFFX1 \mat_i_reg_reg[3][2][0]  ( .D(n153), .CLK(clk), .Q(\mat_i[3][2][0] )
         );
  DFFX1 \mat_r_reg_reg[0][0][11]  ( .D(n152), .CLK(clk), .Q(\mat_r[0][0][11] )
         );
  DFFX1 \mat_r_reg_reg[0][0][10]  ( .D(n151), .CLK(clk), .Q(\mat_r[0][0][10] )
         );
  DFFX1 \mat_r_reg_reg[0][0][9]  ( .D(n150), .CLK(clk), .Q(\mat_r[0][0][9] )
         );
  DFFX1 \mat_r_reg_reg[0][0][8]  ( .D(n149), .CLK(clk), .Q(\mat_r[0][0][8] )
         );
  DFFX1 \mat_r_reg_reg[0][0][7]  ( .D(n148), .CLK(clk), .Q(\mat_r[0][0][7] )
         );
  DFFX1 \mat_r_reg_reg[0][0][6]  ( .D(n147), .CLK(clk), .Q(\mat_r[0][0][6] )
         );
  DFFX1 \mat_r_reg_reg[0][0][5]  ( .D(n146), .CLK(clk), .Q(\mat_r[0][0][5] )
         );
  DFFX1 \mat_r_reg_reg[0][0][4]  ( .D(n145), .CLK(clk), .Q(\mat_r[0][0][4] )
         );
  DFFX1 \mat_r_reg_reg[0][0][3]  ( .D(n144), .CLK(clk), .Q(\mat_r[0][0][3] )
         );
  DFFX1 \mat_r_reg_reg[0][0][2]  ( .D(n143), .CLK(clk), .Q(\mat_r[0][0][2] )
         );
  DFFX1 \mat_r_reg_reg[0][0][1]  ( .D(n142), .CLK(clk), .Q(\mat_r[0][0][1] )
         );
  DFFX1 \mat_r_reg_reg[0][0][0]  ( .D(n141), .CLK(clk), .Q(\mat_r[0][0][0] )
         );
  DFFX1 \mat_r_reg_reg[1][0][11]  ( .D(n140), .CLK(clk), .Q(\mat_r[1][0][11] )
         );
  DFFX1 \mat_r_reg_reg[1][0][10]  ( .D(n139), .CLK(clk), .Q(\mat_r[1][0][10] )
         );
  DFFX1 \mat_r_reg_reg[1][0][9]  ( .D(n138), .CLK(clk), .Q(\mat_r[1][0][9] )
         );
  DFFX1 \mat_r_reg_reg[1][0][8]  ( .D(n137), .CLK(clk), .Q(\mat_r[1][0][8] )
         );
  DFFX1 \mat_r_reg_reg[1][0][7]  ( .D(n136), .CLK(clk), .Q(\mat_r[1][0][7] )
         );
  DFFX1 \mat_r_reg_reg[1][0][6]  ( .D(n135), .CLK(clk), .Q(\mat_r[1][0][6] )
         );
  DFFX1 \mat_r_reg_reg[1][0][5]  ( .D(n134), .CLK(clk), .Q(\mat_r[1][0][5] )
         );
  DFFX1 \mat_r_reg_reg[1][0][4]  ( .D(n133), .CLK(clk), .Q(\mat_r[1][0][4] )
         );
  DFFX1 \mat_r_reg_reg[1][0][3]  ( .D(n132), .CLK(clk), .Q(\mat_r[1][0][3] )
         );
  DFFX1 \mat_r_reg_reg[1][0][2]  ( .D(n131), .CLK(clk), .Q(\mat_r[1][0][2] )
         );
  DFFX1 \mat_r_reg_reg[1][0][1]  ( .D(n130), .CLK(clk), .Q(\mat_r[1][0][1] )
         );
  DFFX1 \mat_r_reg_reg[1][0][0]  ( .D(n129), .CLK(clk), .Q(\mat_r[1][0][0] )
         );
  DFFX1 \mat_r_reg_reg[1][1][11]  ( .D(n128), .CLK(clk), .Q(\mat_r[1][1][11] )
         );
  DFFX1 \mat_r_reg_reg[1][1][10]  ( .D(n127), .CLK(clk), .Q(\mat_r[1][1][10] )
         );
  DFFX1 \mat_r_reg_reg[1][1][9]  ( .D(n126), .CLK(clk), .Q(\mat_r[1][1][9] )
         );
  DFFX1 \mat_r_reg_reg[1][1][8]  ( .D(n125), .CLK(clk), .Q(\mat_r[1][1][8] )
         );
  DFFX1 \mat_r_reg_reg[1][1][7]  ( .D(n124), .CLK(clk), .Q(\mat_r[1][1][7] )
         );
  DFFX1 \mat_r_reg_reg[1][1][6]  ( .D(n123), .CLK(clk), .Q(\mat_r[1][1][6] )
         );
  DFFX1 \mat_r_reg_reg[1][1][5]  ( .D(n122), .CLK(clk), .Q(\mat_r[1][1][5] )
         );
  DFFX1 \mat_r_reg_reg[1][1][4]  ( .D(n121), .CLK(clk), .Q(\mat_r[1][1][4] )
         );
  DFFX1 \mat_r_reg_reg[1][1][3]  ( .D(n120), .CLK(clk), .Q(\mat_r[1][1][3] )
         );
  DFFX1 \mat_r_reg_reg[1][1][2]  ( .D(n119), .CLK(clk), .Q(\mat_r[1][1][2] )
         );
  DFFX1 \mat_r_reg_reg[1][1][1]  ( .D(n118), .CLK(clk), .Q(\mat_r[1][1][1] )
         );
  DFFX1 \mat_r_reg_reg[1][1][0]  ( .D(n117), .CLK(clk), .Q(\mat_r[1][1][0] )
         );
  DFFX1 \mat_r_reg_reg[2][0][11]  ( .D(n116), .CLK(clk), .Q(\mat_r[2][0][11] )
         );
  DFFX1 \mat_r_reg_reg[2][0][10]  ( .D(n115), .CLK(clk), .Q(\mat_r[2][0][10] )
         );
  DFFX1 \mat_r_reg_reg[2][0][9]  ( .D(n114), .CLK(clk), .Q(\mat_r[2][0][9] )
         );
  DFFX1 \mat_r_reg_reg[2][0][8]  ( .D(n113), .CLK(clk), .Q(\mat_r[2][0][8] )
         );
  DFFX1 \mat_r_reg_reg[2][0][7]  ( .D(n112), .CLK(clk), .Q(\mat_r[2][0][7] )
         );
  DFFX1 \mat_r_reg_reg[2][0][6]  ( .D(n111), .CLK(clk), .Q(\mat_r[2][0][6] )
         );
  DFFX1 \mat_r_reg_reg[2][0][5]  ( .D(n110), .CLK(clk), .Q(\mat_r[2][0][5] )
         );
  DFFX1 \mat_r_reg_reg[2][0][4]  ( .D(n109), .CLK(clk), .Q(\mat_r[2][0][4] )
         );
  DFFX1 \mat_r_reg_reg[2][0][3]  ( .D(n108), .CLK(clk), .Q(\mat_r[2][0][3] )
         );
  DFFX1 \mat_r_reg_reg[2][0][2]  ( .D(n107), .CLK(clk), .Q(\mat_r[2][0][2] )
         );
  DFFX1 \mat_r_reg_reg[2][0][1]  ( .D(n106), .CLK(clk), .Q(\mat_r[2][0][1] )
         );
  DFFX1 \mat_r_reg_reg[2][0][0]  ( .D(n105), .CLK(clk), .Q(\mat_r[2][0][0] )
         );
  DFFX1 \mat_r_reg_reg[2][1][11]  ( .D(n104), .CLK(clk), .Q(\mat_r[2][1][11] )
         );
  DFFX1 \mat_r_reg_reg[2][1][10]  ( .D(n103), .CLK(clk), .Q(\mat_r[2][1][10] )
         );
  DFFX1 \mat_r_reg_reg[2][1][9]  ( .D(n102), .CLK(clk), .Q(\mat_r[2][1][9] )
         );
  DFFX1 \mat_r_reg_reg[2][1][8]  ( .D(n101), .CLK(clk), .Q(\mat_r[2][1][8] )
         );
  DFFX1 \mat_r_reg_reg[2][1][7]  ( .D(n100), .CLK(clk), .Q(\mat_r[2][1][7] )
         );
  DFFX1 \mat_r_reg_reg[2][1][6]  ( .D(n99), .CLK(clk), .Q(\mat_r[2][1][6] ) );
  DFFX1 \mat_r_reg_reg[2][1][5]  ( .D(n98), .CLK(clk), .Q(\mat_r[2][1][5] ) );
  DFFX1 \mat_r_reg_reg[2][1][4]  ( .D(n97), .CLK(clk), .Q(\mat_r[2][1][4] ) );
  DFFX1 \mat_r_reg_reg[2][1][3]  ( .D(n96), .CLK(clk), .Q(\mat_r[2][1][3] ) );
  DFFX1 \mat_r_reg_reg[2][1][2]  ( .D(n95), .CLK(clk), .Q(\mat_r[2][1][2] ) );
  DFFX1 \mat_r_reg_reg[2][1][1]  ( .D(n94), .CLK(clk), .Q(\mat_r[2][1][1] ) );
  DFFX1 \mat_r_reg_reg[2][1][0]  ( .D(n93), .CLK(clk), .Q(\mat_r[2][1][0] ) );
  DFFX1 \mat_r_reg_reg[2][2][11]  ( .D(n92), .CLK(clk), .Q(\mat_r[2][2][11] )
         );
  DFFX1 \mat_r_reg_reg[2][2][10]  ( .D(n91), .CLK(clk), .Q(\mat_r[2][2][10] )
         );
  DFFX1 \mat_r_reg_reg[2][2][9]  ( .D(n90), .CLK(clk), .Q(\mat_r[2][2][9] ) );
  DFFX1 \mat_r_reg_reg[2][2][8]  ( .D(n89), .CLK(clk), .Q(\mat_r[2][2][8] ) );
  DFFX1 \mat_r_reg_reg[2][2][7]  ( .D(n88), .CLK(clk), .Q(\mat_r[2][2][7] ) );
  DFFX1 \mat_r_reg_reg[2][2][6]  ( .D(n87), .CLK(clk), .Q(\mat_r[2][2][6] ) );
  DFFX1 \mat_r_reg_reg[2][2][5]  ( .D(n86), .CLK(clk), .Q(\mat_r[2][2][5] ) );
  DFFX1 \mat_r_reg_reg[2][2][4]  ( .D(n85), .CLK(clk), .Q(\mat_r[2][2][4] ) );
  DFFX1 \mat_r_reg_reg[2][2][3]  ( .D(n84), .CLK(clk), .Q(\mat_r[2][2][3] ) );
  DFFX1 \mat_r_reg_reg[2][2][2]  ( .D(n83), .CLK(clk), .Q(\mat_r[2][2][2] ) );
  DFFX1 \mat_r_reg_reg[2][2][1]  ( .D(n82), .CLK(clk), .Q(\mat_r[2][2][1] ) );
  DFFX1 \mat_r_reg_reg[2][2][0]  ( .D(n81), .CLK(clk), .Q(\mat_r[2][2][0] ) );
  DFFX1 \mat_r_reg_reg[3][0][11]  ( .D(n80), .CLK(clk), .Q(\mat_r[3][0][11] )
         );
  DFFX1 \mat_r_reg_reg[3][0][10]  ( .D(n79), .CLK(clk), .Q(\mat_r[3][0][10] )
         );
  DFFX1 \mat_r_reg_reg[3][0][9]  ( .D(n78), .CLK(clk), .Q(\mat_r[3][0][9] ) );
  DFFX1 \mat_r_reg_reg[3][0][8]  ( .D(n77), .CLK(clk), .Q(\mat_r[3][0][8] ) );
  DFFX1 \mat_r_reg_reg[3][0][7]  ( .D(n76), .CLK(clk), .Q(\mat_r[3][0][7] ) );
  DFFX1 \mat_r_reg_reg[3][0][6]  ( .D(n75), .CLK(clk), .Q(\mat_r[3][0][6] ) );
  DFFX1 \mat_r_reg_reg[3][0][5]  ( .D(n74), .CLK(clk), .Q(\mat_r[3][0][5] ) );
  DFFX1 \mat_r_reg_reg[3][0][4]  ( .D(n73), .CLK(clk), .Q(\mat_r[3][0][4] ) );
  DFFX1 \mat_r_reg_reg[3][0][3]  ( .D(n72), .CLK(clk), .Q(\mat_r[3][0][3] ) );
  DFFX1 \mat_r_reg_reg[3][0][2]  ( .D(n71), .CLK(clk), .Q(\mat_r[3][0][2] ) );
  DFFX1 \mat_r_reg_reg[3][0][1]  ( .D(n70), .CLK(clk), .Q(\mat_r[3][0][1] ) );
  DFFX1 \mat_r_reg_reg[3][0][0]  ( .D(n69), .CLK(clk), .Q(\mat_r[3][0][0] ) );
  DFFX1 \mat_r_reg_reg[3][1][11]  ( .D(n68), .CLK(clk), .Q(\mat_r[3][1][11] )
         );
  DFFX1 \mat_r_reg_reg[3][1][10]  ( .D(n67), .CLK(clk), .Q(\mat_r[3][1][10] )
         );
  DFFX1 \mat_r_reg_reg[3][1][9]  ( .D(n66), .CLK(clk), .Q(\mat_r[3][1][9] ) );
  DFFX1 \mat_r_reg_reg[3][1][8]  ( .D(n65), .CLK(clk), .Q(\mat_r[3][1][8] ) );
  DFFX1 \mat_r_reg_reg[3][1][7]  ( .D(n64), .CLK(clk), .Q(\mat_r[3][1][7] ) );
  DFFX1 \mat_r_reg_reg[3][1][6]  ( .D(n63), .CLK(clk), .Q(\mat_r[3][1][6] ) );
  DFFX1 \mat_r_reg_reg[3][1][5]  ( .D(n62), .CLK(clk), .Q(\mat_r[3][1][5] ) );
  DFFX1 \mat_r_reg_reg[3][1][4]  ( .D(n61), .CLK(clk), .Q(\mat_r[3][1][4] ) );
  DFFX1 \mat_r_reg_reg[3][1][3]  ( .D(n60), .CLK(clk), .Q(\mat_r[3][1][3] ) );
  DFFX1 \mat_r_reg_reg[3][1][2]  ( .D(n59), .CLK(clk), .Q(\mat_r[3][1][2] ) );
  DFFX1 \mat_r_reg_reg[3][1][1]  ( .D(n58), .CLK(clk), .Q(\mat_r[3][1][1] ) );
  DFFX1 \mat_r_reg_reg[3][1][0]  ( .D(n57), .CLK(clk), .Q(\mat_r[3][1][0] ) );
  DFFX1 \mat_r_reg_reg[3][2][11]  ( .D(n56), .CLK(clk), .Q(\mat_r[3][2][11] )
         );
  DFFX1 \mat_r_reg_reg[3][2][10]  ( .D(n55), .CLK(clk), .Q(\mat_r[3][2][10] )
         );
  DFFX1 \mat_r_reg_reg[3][2][9]  ( .D(n54), .CLK(clk), .Q(\mat_r[3][2][9] ) );
  DFFX1 \mat_r_reg_reg[3][2][8]  ( .D(n53), .CLK(clk), .Q(\mat_r[3][2][8] ) );
  DFFX1 \mat_r_reg_reg[3][2][7]  ( .D(n52), .CLK(clk), .Q(\mat_r[3][2][7] ) );
  DFFX1 \mat_r_reg_reg[3][2][6]  ( .D(n51), .CLK(clk), .Q(\mat_r[3][2][6] ) );
  DFFX1 \mat_r_reg_reg[3][2][5]  ( .D(n50), .CLK(clk), .Q(\mat_r[3][2][5] ) );
  DFFX1 \mat_r_reg_reg[3][2][4]  ( .D(n49), .CLK(clk), .Q(\mat_r[3][2][4] ) );
  DFFX1 \mat_r_reg_reg[3][2][3]  ( .D(n48), .CLK(clk), .Q(\mat_r[3][2][3] ) );
  DFFX1 \mat_r_reg_reg[3][2][2]  ( .D(n47), .CLK(clk), .Q(\mat_r[3][2][2] ) );
  DFFX1 \mat_r_reg_reg[3][2][1]  ( .D(n46), .CLK(clk), .Q(\mat_r[3][2][1] ) );
  DFFX1 \mat_r_reg_reg[3][2][0]  ( .D(n45), .CLK(clk), .Q(\mat_r[3][2][0] ) );
  DFFX1 \mat_r_reg_reg[3][3][11]  ( .D(n44), .CLK(clk), .Q(\mat_r[3][3][11] )
         );
  DFFX1 \mat_r_reg_reg[3][3][10]  ( .D(n43), .CLK(clk), .Q(\mat_r[3][3][10] )
         );
  DFFX1 \mat_r_reg_reg[3][3][9]  ( .D(n42), .CLK(clk), .Q(\mat_r[3][3][9] ) );
  DFFX1 \mat_r_reg_reg[3][3][8]  ( .D(n41), .CLK(clk), .Q(\mat_r[3][3][8] ) );
  DFFX1 \mat_r_reg_reg[3][3][7]  ( .D(n40), .CLK(clk), .Q(\mat_r[3][3][7] ) );
  DFFX1 \mat_r_reg_reg[3][3][6]  ( .D(n39), .CLK(clk), .Q(\mat_r[3][3][6] ) );
  DFFX1 \mat_r_reg_reg[3][3][5]  ( .D(n38), .CLK(clk), .Q(\mat_r[3][3][5] ) );
  DFFX1 \mat_r_reg_reg[3][3][4]  ( .D(n37), .CLK(clk), .Q(\mat_r[3][3][4] ) );
  DFFX1 \mat_r_reg_reg[3][3][3]  ( .D(n36), .CLK(clk), .Q(\mat_r[3][3][3] ) );
  DFFX1 \mat_r_reg_reg[3][3][2]  ( .D(n35), .CLK(clk), .Q(\mat_r[3][3][2] ) );
  DFFX1 \mat_r_reg_reg[3][3][1]  ( .D(n34), .CLK(clk), .Q(\mat_r[3][3][1] ) );
  DFFX1 \mat_r_reg_reg[3][3][0]  ( .D(n33), .CLK(clk), .Q(\mat_r[3][3][0] ) );
  AO22X1 U21 ( .IN1(single_in_r[0]), .IN2(n328), .IN3(\mat_r[3][3][0] ), .IN4(
        n17), .Q(n33) );
  AO22X1 U22 ( .IN1(single_in_r[1]), .IN2(n328), .IN3(\mat_r[3][3][1] ), .IN4(
        n17), .Q(n34) );
  AO22X1 U23 ( .IN1(single_in_r[2]), .IN2(n328), .IN3(\mat_r[3][3][2] ), .IN4(
        n17), .Q(n35) );
  AO22X1 U24 ( .IN1(single_in_r[3]), .IN2(n328), .IN3(\mat_r[3][3][3] ), .IN4(
        n17), .Q(n36) );
  AO22X1 U25 ( .IN1(single_in_r[4]), .IN2(n328), .IN3(\mat_r[3][3][4] ), .IN4(
        n17), .Q(n37) );
  AO22X1 U26 ( .IN1(single_in_r[5]), .IN2(n328), .IN3(\mat_r[3][3][5] ), .IN4(
        n17), .Q(n38) );
  AO22X1 U27 ( .IN1(single_in_r[6]), .IN2(n328), .IN3(\mat_r[3][3][6] ), .IN4(
        n17), .Q(n39) );
  AO22X1 U28 ( .IN1(single_in_r[7]), .IN2(n328), .IN3(\mat_r[3][3][7] ), .IN4(
        n17), .Q(n40) );
  AO22X1 U29 ( .IN1(single_in_r[8]), .IN2(n328), .IN3(\mat_r[3][3][8] ), .IN4(
        n17), .Q(n41) );
  AO22X1 U30 ( .IN1(single_in_r[9]), .IN2(n328), .IN3(\mat_r[3][3][9] ), .IN4(
        n17), .Q(n42) );
  AO22X1 U31 ( .IN1(single_in_r[10]), .IN2(n328), .IN3(\mat_r[3][3][10] ), 
        .IN4(n17), .Q(n43) );
  AO22X1 U32 ( .IN1(single_in_r[11]), .IN2(n328), .IN3(\mat_r[3][3][11] ), 
        .IN4(n17), .Q(n44) );
  AO22X1 U33 ( .IN1(n320), .IN2(single_in_r[0]), .IN3(\mat_r[3][2][0] ), .IN4(
        n319), .Q(n45) );
  AO22X1 U34 ( .IN1(n320), .IN2(single_in_r[1]), .IN3(\mat_r[3][2][1] ), .IN4(
        n319), .Q(n46) );
  AO22X1 U35 ( .IN1(n320), .IN2(single_in_r[2]), .IN3(\mat_r[3][2][2] ), .IN4(
        n319), .Q(n47) );
  AO22X1 U36 ( .IN1(n320), .IN2(single_in_r[3]), .IN3(\mat_r[3][2][3] ), .IN4(
        n319), .Q(n48) );
  AO22X1 U37 ( .IN1(n320), .IN2(single_in_r[4]), .IN3(\mat_r[3][2][4] ), .IN4(
        n319), .Q(n49) );
  AO22X1 U38 ( .IN1(n321), .IN2(single_in_r[5]), .IN3(\mat_r[3][2][5] ), .IN4(
        n319), .Q(n50) );
  AO22X1 U39 ( .IN1(n321), .IN2(single_in_r[6]), .IN3(\mat_r[3][2][6] ), .IN4(
        n319), .Q(n51) );
  AO22X1 U40 ( .IN1(n321), .IN2(single_in_r[7]), .IN3(\mat_r[3][2][7] ), .IN4(
        n319), .Q(n52) );
  AO22X1 U41 ( .IN1(n321), .IN2(single_in_r[8]), .IN3(\mat_r[3][2][8] ), .IN4(
        n319), .Q(n53) );
  AO22X1 U42 ( .IN1(n321), .IN2(single_in_r[9]), .IN3(\mat_r[3][2][9] ), .IN4(
        n319), .Q(n54) );
  AO22X1 U43 ( .IN1(n321), .IN2(single_in_r[10]), .IN3(\mat_r[3][2][10] ), 
        .IN4(n319), .Q(n55) );
  AO22X1 U44 ( .IN1(n321), .IN2(single_in_r[11]), .IN3(\mat_r[3][2][11] ), 
        .IN4(n319), .Q(n56) );
  AO22X1 U45 ( .IN1(n315), .IN2(single_in_r[0]), .IN3(\mat_r[3][1][0] ), .IN4(
        n314), .Q(n57) );
  AO22X1 U46 ( .IN1(n315), .IN2(single_in_r[1]), .IN3(\mat_r[3][1][1] ), .IN4(
        n314), .Q(n58) );
  AO22X1 U47 ( .IN1(n315), .IN2(single_in_r[2]), .IN3(\mat_r[3][1][2] ), .IN4(
        n314), .Q(n59) );
  AO22X1 U48 ( .IN1(n315), .IN2(single_in_r[3]), .IN3(\mat_r[3][1][3] ), .IN4(
        n314), .Q(n60) );
  AO22X1 U49 ( .IN1(n315), .IN2(single_in_r[4]), .IN3(\mat_r[3][1][4] ), .IN4(
        n314), .Q(n61) );
  AO22X1 U50 ( .IN1(n316), .IN2(single_in_r[5]), .IN3(\mat_r[3][1][5] ), .IN4(
        n314), .Q(n62) );
  AO22X1 U51 ( .IN1(n316), .IN2(single_in_r[6]), .IN3(\mat_r[3][1][6] ), .IN4(
        n314), .Q(n63) );
  AO22X1 U52 ( .IN1(n316), .IN2(single_in_r[7]), .IN3(\mat_r[3][1][7] ), .IN4(
        n314), .Q(n64) );
  AO22X1 U53 ( .IN1(n316), .IN2(single_in_r[8]), .IN3(\mat_r[3][1][8] ), .IN4(
        n314), .Q(n65) );
  AO22X1 U54 ( .IN1(n316), .IN2(single_in_r[9]), .IN3(\mat_r[3][1][9] ), .IN4(
        n314), .Q(n66) );
  AO22X1 U55 ( .IN1(n316), .IN2(single_in_r[10]), .IN3(\mat_r[3][1][10] ), 
        .IN4(n314), .Q(n67) );
  AO22X1 U56 ( .IN1(n316), .IN2(single_in_r[11]), .IN3(\mat_r[3][1][11] ), 
        .IN4(n314), .Q(n68) );
  AO22X1 U57 ( .IN1(n310), .IN2(single_in_r[0]), .IN3(\mat_r[3][0][0] ), .IN4(
        n309), .Q(n69) );
  AO22X1 U58 ( .IN1(n310), .IN2(single_in_r[1]), .IN3(\mat_r[3][0][1] ), .IN4(
        n309), .Q(n70) );
  AO22X1 U59 ( .IN1(n310), .IN2(single_in_r[2]), .IN3(\mat_r[3][0][2] ), .IN4(
        n309), .Q(n71) );
  AO22X1 U60 ( .IN1(n310), .IN2(single_in_r[3]), .IN3(\mat_r[3][0][3] ), .IN4(
        n309), .Q(n72) );
  AO22X1 U61 ( .IN1(n310), .IN2(single_in_r[4]), .IN3(\mat_r[3][0][4] ), .IN4(
        n309), .Q(n73) );
  AO22X1 U62 ( .IN1(n311), .IN2(single_in_r[5]), .IN3(\mat_r[3][0][5] ), .IN4(
        n309), .Q(n74) );
  AO22X1 U63 ( .IN1(n311), .IN2(single_in_r[6]), .IN3(\mat_r[3][0][6] ), .IN4(
        n309), .Q(n75) );
  AO22X1 U64 ( .IN1(n311), .IN2(single_in_r[7]), .IN3(\mat_r[3][0][7] ), .IN4(
        n309), .Q(n76) );
  AO22X1 U65 ( .IN1(n311), .IN2(single_in_r[8]), .IN3(\mat_r[3][0][8] ), .IN4(
        n309), .Q(n77) );
  AO22X1 U66 ( .IN1(n311), .IN2(single_in_r[9]), .IN3(\mat_r[3][0][9] ), .IN4(
        n309), .Q(n78) );
  AO22X1 U67 ( .IN1(n311), .IN2(single_in_r[10]), .IN3(\mat_r[3][0][10] ), 
        .IN4(n309), .Q(n79) );
  AO22X1 U68 ( .IN1(n311), .IN2(single_in_r[11]), .IN3(\mat_r[3][0][11] ), 
        .IN4(n309), .Q(n80) );
  AO22X1 U69 ( .IN1(n326), .IN2(single_in_r[0]), .IN3(\mat_r[2][2][0] ), .IN4(
        n22), .Q(n81) );
  AO22X1 U70 ( .IN1(n326), .IN2(single_in_r[1]), .IN3(\mat_r[2][2][1] ), .IN4(
        n22), .Q(n82) );
  AO22X1 U71 ( .IN1(n326), .IN2(single_in_r[2]), .IN3(\mat_r[2][2][2] ), .IN4(
        n22), .Q(n83) );
  AO22X1 U72 ( .IN1(n326), .IN2(single_in_r[3]), .IN3(\mat_r[2][2][3] ), .IN4(
        n22), .Q(n84) );
  AO22X1 U73 ( .IN1(n326), .IN2(single_in_r[4]), .IN3(\mat_r[2][2][4] ), .IN4(
        n22), .Q(n85) );
  AO22X1 U74 ( .IN1(n326), .IN2(single_in_r[5]), .IN3(\mat_r[2][2][5] ), .IN4(
        n22), .Q(n86) );
  AO22X1 U75 ( .IN1(n326), .IN2(single_in_r[6]), .IN3(\mat_r[2][2][6] ), .IN4(
        n22), .Q(n87) );
  AO22X1 U76 ( .IN1(n326), .IN2(single_in_r[7]), .IN3(\mat_r[2][2][7] ), .IN4(
        n22), .Q(n88) );
  AO22X1 U77 ( .IN1(n326), .IN2(single_in_r[8]), .IN3(\mat_r[2][2][8] ), .IN4(
        n22), .Q(n89) );
  AO22X1 U78 ( .IN1(n326), .IN2(single_in_r[9]), .IN3(\mat_r[2][2][9] ), .IN4(
        n22), .Q(n90) );
  AO22X1 U79 ( .IN1(n326), .IN2(single_in_r[10]), .IN3(\mat_r[2][2][10] ), 
        .IN4(n22), .Q(n91) );
  AO22X1 U80 ( .IN1(n326), .IN2(single_in_r[11]), .IN3(\mat_r[2][2][11] ), 
        .IN4(n22), .Q(n92) );
  AO22X1 U81 ( .IN1(n305), .IN2(single_in_r[0]), .IN3(\mat_r[2][1][0] ), .IN4(
        n304), .Q(n93) );
  AO22X1 U82 ( .IN1(n305), .IN2(single_in_r[1]), .IN3(\mat_r[2][1][1] ), .IN4(
        n304), .Q(n94) );
  AO22X1 U83 ( .IN1(n305), .IN2(single_in_r[2]), .IN3(\mat_r[2][1][2] ), .IN4(
        n304), .Q(n95) );
  AO22X1 U84 ( .IN1(n305), .IN2(single_in_r[3]), .IN3(\mat_r[2][1][3] ), .IN4(
        n304), .Q(n96) );
  AO22X1 U85 ( .IN1(n305), .IN2(single_in_r[4]), .IN3(\mat_r[2][1][4] ), .IN4(
        n304), .Q(n97) );
  AO22X1 U86 ( .IN1(n306), .IN2(single_in_r[5]), .IN3(\mat_r[2][1][5] ), .IN4(
        n304), .Q(n98) );
  AO22X1 U87 ( .IN1(n306), .IN2(single_in_r[6]), .IN3(\mat_r[2][1][6] ), .IN4(
        n304), .Q(n99) );
  AO22X1 U88 ( .IN1(n306), .IN2(single_in_r[7]), .IN3(\mat_r[2][1][7] ), .IN4(
        n304), .Q(n100) );
  AO22X1 U89 ( .IN1(n306), .IN2(single_in_r[8]), .IN3(\mat_r[2][1][8] ), .IN4(
        n304), .Q(n101) );
  AO22X1 U90 ( .IN1(n306), .IN2(single_in_r[9]), .IN3(\mat_r[2][1][9] ), .IN4(
        n304), .Q(n102) );
  AO22X1 U91 ( .IN1(n306), .IN2(single_in_r[10]), .IN3(\mat_r[2][1][10] ), 
        .IN4(n304), .Q(n103) );
  AO22X1 U92 ( .IN1(n306), .IN2(single_in_r[11]), .IN3(\mat_r[2][1][11] ), 
        .IN4(n304), .Q(n104) );
  AO22X1 U93 ( .IN1(n300), .IN2(single_in_r[0]), .IN3(\mat_r[2][0][0] ), .IN4(
        n299), .Q(n105) );
  AO22X1 U94 ( .IN1(n300), .IN2(single_in_r[1]), .IN3(\mat_r[2][0][1] ), .IN4(
        n299), .Q(n106) );
  AO22X1 U95 ( .IN1(n300), .IN2(single_in_r[2]), .IN3(\mat_r[2][0][2] ), .IN4(
        n299), .Q(n107) );
  AO22X1 U96 ( .IN1(n300), .IN2(single_in_r[3]), .IN3(\mat_r[2][0][3] ), .IN4(
        n299), .Q(n108) );
  AO22X1 U97 ( .IN1(n300), .IN2(single_in_r[4]), .IN3(\mat_r[2][0][4] ), .IN4(
        n299), .Q(n109) );
  AO22X1 U98 ( .IN1(n301), .IN2(single_in_r[5]), .IN3(\mat_r[2][0][5] ), .IN4(
        n299), .Q(n110) );
  AO22X1 U99 ( .IN1(n301), .IN2(single_in_r[6]), .IN3(\mat_r[2][0][6] ), .IN4(
        n299), .Q(n111) );
  AO22X1 U100 ( .IN1(n301), .IN2(single_in_r[7]), .IN3(\mat_r[2][0][7] ), 
        .IN4(n299), .Q(n112) );
  AO22X1 U101 ( .IN1(n301), .IN2(single_in_r[8]), .IN3(\mat_r[2][0][8] ), 
        .IN4(n299), .Q(n113) );
  AO22X1 U102 ( .IN1(n301), .IN2(single_in_r[9]), .IN3(\mat_r[2][0][9] ), 
        .IN4(n299), .Q(n114) );
  AO22X1 U103 ( .IN1(n301), .IN2(single_in_r[10]), .IN3(\mat_r[2][0][10] ), 
        .IN4(n299), .Q(n115) );
  AO22X1 U104 ( .IN1(n301), .IN2(single_in_r[11]), .IN3(\mat_r[2][0][11] ), 
        .IN4(n299), .Q(n116) );
  AO22X1 U105 ( .IN1(n327), .IN2(single_in_r[0]), .IN3(\mat_r[1][1][0] ), 
        .IN4(n25), .Q(n117) );
  AO22X1 U106 ( .IN1(n327), .IN2(single_in_r[1]), .IN3(\mat_r[1][1][1] ), 
        .IN4(n25), .Q(n118) );
  AO22X1 U107 ( .IN1(n327), .IN2(single_in_r[2]), .IN3(\mat_r[1][1][2] ), 
        .IN4(n25), .Q(n119) );
  AO22X1 U108 ( .IN1(n327), .IN2(single_in_r[3]), .IN3(\mat_r[1][1][3] ), 
        .IN4(n25), .Q(n120) );
  AO22X1 U109 ( .IN1(n327), .IN2(single_in_r[4]), .IN3(\mat_r[1][1][4] ), 
        .IN4(n25), .Q(n121) );
  AO22X1 U110 ( .IN1(n327), .IN2(single_in_r[5]), .IN3(\mat_r[1][1][5] ), 
        .IN4(n25), .Q(n122) );
  AO22X1 U111 ( .IN1(n327), .IN2(single_in_r[6]), .IN3(\mat_r[1][1][6] ), 
        .IN4(n25), .Q(n123) );
  AO22X1 U112 ( .IN1(n327), .IN2(single_in_r[7]), .IN3(\mat_r[1][1][7] ), 
        .IN4(n25), .Q(n124) );
  AO22X1 U113 ( .IN1(n327), .IN2(single_in_r[8]), .IN3(\mat_r[1][1][8] ), 
        .IN4(n25), .Q(n125) );
  AO22X1 U114 ( .IN1(n327), .IN2(single_in_r[9]), .IN3(\mat_r[1][1][9] ), 
        .IN4(n25), .Q(n126) );
  AO22X1 U115 ( .IN1(n327), .IN2(single_in_r[10]), .IN3(\mat_r[1][1][10] ), 
        .IN4(n25), .Q(n127) );
  AO22X1 U116 ( .IN1(n327), .IN2(single_in_r[11]), .IN3(\mat_r[1][1][11] ), 
        .IN4(n25), .Q(n128) );
  AO22X1 U118 ( .IN1(n295), .IN2(single_in_r[0]), .IN3(\mat_r[1][0][0] ), 
        .IN4(n294), .Q(n129) );
  AO22X1 U119 ( .IN1(n295), .IN2(single_in_r[1]), .IN3(\mat_r[1][0][1] ), 
        .IN4(n294), .Q(n130) );
  AO22X1 U120 ( .IN1(n295), .IN2(single_in_r[2]), .IN3(\mat_r[1][0][2] ), 
        .IN4(n294), .Q(n131) );
  AO22X1 U121 ( .IN1(n295), .IN2(single_in_r[3]), .IN3(\mat_r[1][0][3] ), 
        .IN4(n294), .Q(n132) );
  AO22X1 U122 ( .IN1(n295), .IN2(single_in_r[4]), .IN3(\mat_r[1][0][4] ), 
        .IN4(n294), .Q(n133) );
  AO22X1 U123 ( .IN1(n296), .IN2(single_in_r[5]), .IN3(\mat_r[1][0][5] ), 
        .IN4(n294), .Q(n134) );
  AO22X1 U124 ( .IN1(n296), .IN2(single_in_r[6]), .IN3(\mat_r[1][0][6] ), 
        .IN4(n294), .Q(n135) );
  AO22X1 U125 ( .IN1(n296), .IN2(single_in_r[7]), .IN3(\mat_r[1][0][7] ), 
        .IN4(n294), .Q(n136) );
  AO22X1 U126 ( .IN1(n296), .IN2(single_in_r[8]), .IN3(\mat_r[1][0][8] ), 
        .IN4(n294), .Q(n137) );
  AO22X1 U127 ( .IN1(n296), .IN2(single_in_r[9]), .IN3(\mat_r[1][0][9] ), 
        .IN4(n294), .Q(n138) );
  AO22X1 U128 ( .IN1(n296), .IN2(single_in_r[10]), .IN3(\mat_r[1][0][10] ), 
        .IN4(n294), .Q(n139) );
  AO22X1 U129 ( .IN1(n296), .IN2(single_in_r[11]), .IN3(\mat_r[1][0][11] ), 
        .IN4(n294), .Q(n140) );
  AO22X1 U130 ( .IN1(n325), .IN2(single_in_r[0]), .IN3(\mat_r[0][0][0] ), 
        .IN4(n28), .Q(n141) );
  AO22X1 U131 ( .IN1(n325), .IN2(single_in_r[1]), .IN3(\mat_r[0][0][1] ), 
        .IN4(n28), .Q(n142) );
  AO22X1 U132 ( .IN1(n325), .IN2(single_in_r[2]), .IN3(\mat_r[0][0][2] ), 
        .IN4(n28), .Q(n143) );
  AO22X1 U133 ( .IN1(n325), .IN2(single_in_r[3]), .IN3(\mat_r[0][0][3] ), 
        .IN4(n28), .Q(n144) );
  AO22X1 U134 ( .IN1(n325), .IN2(single_in_r[4]), .IN3(\mat_r[0][0][4] ), 
        .IN4(n28), .Q(n145) );
  AO22X1 U135 ( .IN1(n325), .IN2(single_in_r[5]), .IN3(\mat_r[0][0][5] ), 
        .IN4(n28), .Q(n146) );
  AO22X1 U136 ( .IN1(n325), .IN2(single_in_r[6]), .IN3(\mat_r[0][0][6] ), 
        .IN4(n28), .Q(n147) );
  AO22X1 U137 ( .IN1(n325), .IN2(single_in_r[7]), .IN3(\mat_r[0][0][7] ), 
        .IN4(n28), .Q(n148) );
  AO22X1 U138 ( .IN1(n325), .IN2(single_in_r[8]), .IN3(\mat_r[0][0][8] ), 
        .IN4(n28), .Q(n149) );
  AO22X1 U139 ( .IN1(n325), .IN2(single_in_r[9]), .IN3(\mat_r[0][0][9] ), 
        .IN4(n28), .Q(n150) );
  AO22X1 U140 ( .IN1(n325), .IN2(single_in_r[10]), .IN3(\mat_r[0][0][10] ), 
        .IN4(n28), .Q(n151) );
  AO22X1 U141 ( .IN1(n325), .IN2(single_in_r[11]), .IN3(\mat_r[0][0][11] ), 
        .IN4(n28), .Q(n152) );
  AO22X1 U143 ( .IN1(single_in_i[0]), .IN2(n322), .IN3(\mat_i[3][2][0] ), 
        .IN4(n318), .Q(n153) );
  AO22X1 U144 ( .IN1(single_in_i[1]), .IN2(n322), .IN3(\mat_i[3][2][1] ), 
        .IN4(n318), .Q(n154) );
  AO22X1 U145 ( .IN1(single_in_i[2]), .IN2(n322), .IN3(\mat_i[3][2][2] ), 
        .IN4(n318), .Q(n155) );
  AO22X1 U146 ( .IN1(single_in_i[3]), .IN2(n322), .IN3(\mat_i[3][2][3] ), 
        .IN4(n318), .Q(n156) );
  AO22X1 U147 ( .IN1(single_in_i[4]), .IN2(n322), .IN3(\mat_i[3][2][4] ), 
        .IN4(n318), .Q(n157) );
  AO22X1 U148 ( .IN1(single_in_i[5]), .IN2(n322), .IN3(\mat_i[3][2][5] ), 
        .IN4(n318), .Q(n158) );
  AO22X1 U149 ( .IN1(single_in_i[6]), .IN2(n322), .IN3(\mat_i[3][2][6] ), 
        .IN4(n318), .Q(n159) );
  AO22X1 U150 ( .IN1(single_in_i[7]), .IN2(n322), .IN3(\mat_i[3][2][7] ), 
        .IN4(n318), .Q(n160) );
  AO22X1 U151 ( .IN1(single_in_i[8]), .IN2(n321), .IN3(\mat_i[3][2][8] ), 
        .IN4(n318), .Q(n161) );
  AO22X1 U152 ( .IN1(single_in_i[9]), .IN2(n322), .IN3(\mat_i[3][2][9] ), 
        .IN4(n318), .Q(n162) );
  AO22X1 U153 ( .IN1(single_in_i[10]), .IN2(n322), .IN3(\mat_i[3][2][10] ), 
        .IN4(n318), .Q(n163) );
  AO22X1 U154 ( .IN1(single_in_i[11]), .IN2(n321), .IN3(\mat_i[3][2][11] ), 
        .IN4(n318), .Q(n164) );
  NAND3X0 U155 ( .IN1(n18), .IN2(n329), .IN3(N11), .QN(n19) );
  AND3X1 U156 ( .IN1(n30), .IN2(row_sel[1]), .IN3(wr_enable), .Q(n18) );
  AO22X1 U157 ( .IN1(single_in_i[0]), .IN2(n317), .IN3(\mat_i[3][1][0] ), 
        .IN4(n313), .Q(n165) );
  AO22X1 U158 ( .IN1(single_in_i[1]), .IN2(n317), .IN3(\mat_i[3][1][1] ), 
        .IN4(n313), .Q(n166) );
  AO22X1 U159 ( .IN1(single_in_i[2]), .IN2(n317), .IN3(\mat_i[3][1][2] ), 
        .IN4(n313), .Q(n167) );
  AO22X1 U160 ( .IN1(single_in_i[3]), .IN2(n317), .IN3(\mat_i[3][1][3] ), 
        .IN4(n313), .Q(n168) );
  AO22X1 U161 ( .IN1(single_in_i[4]), .IN2(n317), .IN3(\mat_i[3][1][4] ), 
        .IN4(n313), .Q(n169) );
  AO22X1 U162 ( .IN1(single_in_i[5]), .IN2(n317), .IN3(\mat_i[3][1][5] ), 
        .IN4(n313), .Q(n170) );
  AO22X1 U163 ( .IN1(single_in_i[6]), .IN2(n317), .IN3(\mat_i[3][1][6] ), 
        .IN4(n313), .Q(n171) );
  AO22X1 U164 ( .IN1(single_in_i[7]), .IN2(n317), .IN3(\mat_i[3][1][7] ), 
        .IN4(n313), .Q(n172) );
  AO22X1 U165 ( .IN1(single_in_i[8]), .IN2(n316), .IN3(\mat_i[3][1][8] ), 
        .IN4(n313), .Q(n173) );
  AO22X1 U166 ( .IN1(single_in_i[9]), .IN2(n317), .IN3(\mat_i[3][1][9] ), 
        .IN4(n313), .Q(n174) );
  AO22X1 U167 ( .IN1(single_in_i[10]), .IN2(n317), .IN3(\mat_i[3][1][10] ), 
        .IN4(n313), .Q(n175) );
  AO22X1 U168 ( .IN1(single_in_i[11]), .IN2(n316), .IN3(\mat_i[3][1][11] ), 
        .IN4(n313), .Q(n176) );
  AO22X1 U169 ( .IN1(single_in_i[0]), .IN2(n312), .IN3(\mat_i[3][0][0] ), 
        .IN4(n308), .Q(n177) );
  AO22X1 U170 ( .IN1(single_in_i[1]), .IN2(n312), .IN3(\mat_i[3][0][1] ), 
        .IN4(n308), .Q(n178) );
  AO22X1 U171 ( .IN1(single_in_i[2]), .IN2(n312), .IN3(\mat_i[3][0][2] ), 
        .IN4(n308), .Q(n179) );
  AO22X1 U172 ( .IN1(single_in_i[3]), .IN2(n312), .IN3(\mat_i[3][0][3] ), 
        .IN4(n308), .Q(n180) );
  AO22X1 U173 ( .IN1(single_in_i[4]), .IN2(n312), .IN3(\mat_i[3][0][4] ), 
        .IN4(n308), .Q(n181) );
  AO22X1 U174 ( .IN1(single_in_i[5]), .IN2(n312), .IN3(\mat_i[3][0][5] ), 
        .IN4(n308), .Q(n182) );
  AO22X1 U175 ( .IN1(single_in_i[6]), .IN2(n312), .IN3(\mat_i[3][0][6] ), 
        .IN4(n308), .Q(n183) );
  AO22X1 U176 ( .IN1(single_in_i[7]), .IN2(n312), .IN3(\mat_i[3][0][7] ), 
        .IN4(n308), .Q(n184) );
  AO22X1 U177 ( .IN1(single_in_i[8]), .IN2(n311), .IN3(\mat_i[3][0][8] ), 
        .IN4(n308), .Q(n185) );
  AO22X1 U178 ( .IN1(single_in_i[9]), .IN2(n312), .IN3(\mat_i[3][0][9] ), 
        .IN4(n308), .Q(n186) );
  AO22X1 U179 ( .IN1(single_in_i[10]), .IN2(n312), .IN3(\mat_i[3][0][10] ), 
        .IN4(n308), .Q(n187) );
  AO22X1 U180 ( .IN1(single_in_i[11]), .IN2(n311), .IN3(\mat_i[3][0][11] ), 
        .IN4(n308), .Q(n188) );
  NAND3X0 U181 ( .IN1(N11), .IN2(N12), .IN3(n29), .QN(n21) );
  AO22X1 U182 ( .IN1(single_in_i[0]), .IN2(n307), .IN3(\mat_i[2][1][0] ), 
        .IN4(n303), .Q(n189) );
  AO22X1 U183 ( .IN1(single_in_i[1]), .IN2(n307), .IN3(\mat_i[2][1][1] ), 
        .IN4(n303), .Q(n190) );
  AO22X1 U184 ( .IN1(single_in_i[2]), .IN2(n307), .IN3(\mat_i[2][1][2] ), 
        .IN4(n303), .Q(n191) );
  AO22X1 U185 ( .IN1(single_in_i[3]), .IN2(n307), .IN3(\mat_i[2][1][3] ), 
        .IN4(n303), .Q(n192) );
  AO22X1 U186 ( .IN1(single_in_i[4]), .IN2(n307), .IN3(\mat_i[2][1][4] ), 
        .IN4(n303), .Q(n193) );
  AO22X1 U187 ( .IN1(single_in_i[5]), .IN2(n307), .IN3(\mat_i[2][1][5] ), 
        .IN4(n303), .Q(n194) );
  AO22X1 U188 ( .IN1(single_in_i[6]), .IN2(n307), .IN3(\mat_i[2][1][6] ), 
        .IN4(n303), .Q(n195) );
  AO22X1 U189 ( .IN1(single_in_i[7]), .IN2(n307), .IN3(\mat_i[2][1][7] ), 
        .IN4(n303), .Q(n196) );
  AO22X1 U190 ( .IN1(single_in_i[8]), .IN2(n306), .IN3(\mat_i[2][1][8] ), 
        .IN4(n303), .Q(n197) );
  AO22X1 U191 ( .IN1(single_in_i[9]), .IN2(n307), .IN3(\mat_i[2][1][9] ), 
        .IN4(n303), .Q(n198) );
  AO22X1 U192 ( .IN1(single_in_i[10]), .IN2(n307), .IN3(\mat_i[2][1][10] ), 
        .IN4(n303), .Q(n199) );
  AO22X1 U193 ( .IN1(single_in_i[11]), .IN2(n306), .IN3(\mat_i[2][1][11] ), 
        .IN4(n303), .Q(n200) );
  AND3X1 U194 ( .IN1(row_sel[0]), .IN2(N12), .IN3(n26), .Q(n31) );
  AO22X1 U195 ( .IN1(single_in_i[0]), .IN2(n302), .IN3(\mat_i[2][0][0] ), 
        .IN4(n298), .Q(n201) );
  AO22X1 U196 ( .IN1(single_in_i[1]), .IN2(n302), .IN3(\mat_i[2][0][1] ), 
        .IN4(n298), .Q(n202) );
  AO22X1 U197 ( .IN1(single_in_i[2]), .IN2(n302), .IN3(\mat_i[2][0][2] ), 
        .IN4(n298), .Q(n203) );
  AO22X1 U198 ( .IN1(single_in_i[3]), .IN2(n302), .IN3(\mat_i[2][0][3] ), 
        .IN4(n298), .Q(n204) );
  AO22X1 U199 ( .IN1(single_in_i[4]), .IN2(n302), .IN3(\mat_i[2][0][4] ), 
        .IN4(n298), .Q(n205) );
  AO22X1 U200 ( .IN1(single_in_i[5]), .IN2(n302), .IN3(\mat_i[2][0][5] ), 
        .IN4(n298), .Q(n206) );
  AO22X1 U201 ( .IN1(single_in_i[6]), .IN2(n302), .IN3(\mat_i[2][0][6] ), 
        .IN4(n298), .Q(n207) );
  AO22X1 U202 ( .IN1(single_in_i[7]), .IN2(n302), .IN3(\mat_i[2][0][7] ), 
        .IN4(n298), .Q(n208) );
  AO22X1 U203 ( .IN1(single_in_i[8]), .IN2(n301), .IN3(\mat_i[2][0][8] ), 
        .IN4(n298), .Q(n209) );
  AO22X1 U204 ( .IN1(single_in_i[9]), .IN2(n302), .IN3(\mat_i[2][0][9] ), 
        .IN4(n298), .Q(n210) );
  AO22X1 U205 ( .IN1(single_in_i[10]), .IN2(n302), .IN3(\mat_i[2][0][10] ), 
        .IN4(n298), .Q(n211) );
  AO22X1 U206 ( .IN1(single_in_i[11]), .IN2(n301), .IN3(\mat_i[2][0][11] ), 
        .IN4(n298), .Q(n212) );
  NAND3X0 U207 ( .IN1(N12), .IN2(n323), .IN3(n29), .QN(n24) );
  AO22X1 U208 ( .IN1(single_in_i[0]), .IN2(n297), .IN3(\mat_i[1][0][0] ), 
        .IN4(n293), .Q(n213) );
  AO22X1 U209 ( .IN1(single_in_i[1]), .IN2(n297), .IN3(\mat_i[1][0][1] ), 
        .IN4(n293), .Q(n214) );
  AO22X1 U210 ( .IN1(single_in_i[2]), .IN2(n297), .IN3(\mat_i[1][0][2] ), 
        .IN4(n293), .Q(n215) );
  AO22X1 U211 ( .IN1(single_in_i[3]), .IN2(n297), .IN3(\mat_i[1][0][3] ), 
        .IN4(n293), .Q(n216) );
  AO22X1 U212 ( .IN1(single_in_i[4]), .IN2(n297), .IN3(\mat_i[1][0][4] ), 
        .IN4(n293), .Q(n217) );
  AO22X1 U213 ( .IN1(single_in_i[5]), .IN2(n297), .IN3(\mat_i[1][0][5] ), 
        .IN4(n293), .Q(n218) );
  AO22X1 U214 ( .IN1(single_in_i[6]), .IN2(n297), .IN3(\mat_i[1][0][6] ), 
        .IN4(n293), .Q(n219) );
  AO22X1 U215 ( .IN1(single_in_i[7]), .IN2(n297), .IN3(\mat_i[1][0][7] ), 
        .IN4(n293), .Q(n220) );
  AO22X1 U216 ( .IN1(single_in_i[8]), .IN2(n296), .IN3(\mat_i[1][0][8] ), 
        .IN4(n293), .Q(n221) );
  AO22X1 U217 ( .IN1(single_in_i[9]), .IN2(n297), .IN3(\mat_i[1][0][9] ), 
        .IN4(n293), .Q(n222) );
  AO22X1 U218 ( .IN1(single_in_i[10]), .IN2(n297), .IN3(\mat_i[1][0][10] ), 
        .IN4(n293), .Q(n223) );
  AO22X1 U219 ( .IN1(single_in_i[11]), .IN2(n296), .IN3(\mat_i[1][0][11] ), 
        .IN4(n293), .Q(n224) );
  NAND3X0 U220 ( .IN1(N11), .IN2(n324), .IN3(n29), .QN(n27) );
  AND2X1 U221 ( .IN1(n26), .IN2(n329), .Q(n29) );
  AND3X1 U222 ( .IN1(n30), .IN2(n330), .IN3(wr_enable), .Q(n26) );
  AOI22X1 U223 ( .IN1(n32), .IN2(row_sel[0]), .IN3(row_sel[1]), .IN4(n324), 
        .QN(n30) );
  NAND2X0 U2 ( .IN1(n31), .IN2(n323), .QN(n23) );
  INVX0 U3 ( .INP(n28), .ZN(n325) );
  NBUFFX2 U4 ( .INP(n1), .Z(n292) );
  NBUFFX2 U5 ( .INP(n1), .Z(n291) );
  INVX0 U6 ( .INP(n20), .ZN(n315) );
  INVX0 U7 ( .INP(n20), .ZN(n317) );
  INVX0 U8 ( .INP(n20), .ZN(n316) );
  NAND3X0 U9 ( .IN1(n323), .IN2(n324), .IN3(n29), .QN(n28) );
  INVX0 U10 ( .INP(n22), .ZN(n326) );
  INVX0 U11 ( .INP(n24), .ZN(n300) );
  INVX0 U12 ( .INP(n21), .ZN(n310) );
  INVX0 U13 ( .INP(n27), .ZN(n295) );
  INVX0 U14 ( .INP(n24), .ZN(n302) );
  INVX0 U15 ( .INP(n24), .ZN(n301) );
  INVX0 U16 ( .INP(n19), .ZN(n320) );
  INVX0 U17 ( .INP(n21), .ZN(n312) );
  INVX0 U18 ( .INP(n27), .ZN(n297) );
  INVX0 U19 ( .INP(n21), .ZN(n311) );
  INVX0 U20 ( .INP(n27), .ZN(n296) );
  INVX0 U117 ( .INP(n19), .ZN(n322) );
  INVX0 U142 ( .INP(n19), .ZN(n321) );
  INVX0 U225 ( .INP(n23), .ZN(n305) );
  INVX0 U226 ( .INP(n23), .ZN(n307) );
  INVX0 U227 ( .INP(n23), .ZN(n306) );
  INVX0 U228 ( .INP(n323), .ZN(n289) );
  INVX0 U229 ( .INP(n323), .ZN(n288) );
  INVX0 U230 ( .INP(n323), .ZN(n290) );
  INVX0 U231 ( .INP(n323), .ZN(n287) );
  INVX0 U232 ( .INP(n324), .ZN(n283) );
  INVX0 U233 ( .INP(n324), .ZN(n285) );
  INVX0 U234 ( .INP(n324), .ZN(n284) );
  NOR2X0 U235 ( .IN1(n324), .IN2(n323), .QN(n1) );
  NAND2X0 U236 ( .IN1(n31), .IN2(N11), .QN(n20) );
  NAND2X1 U237 ( .IN1(n18), .IN2(n323), .QN(n22) );
  INVX0 U238 ( .INP(n17), .ZN(n328) );
  INVX0 U239 ( .INP(n25), .ZN(n327) );
  NAND2X1 U240 ( .IN1(n18), .IN2(row_sel[0]), .QN(n17) );
  NAND3X0 U241 ( .IN1(row_sel[0]), .IN2(n324), .IN3(n26), .QN(n25) );
  INVX0 U242 ( .INP(row_sel[1]), .ZN(n330) );
  OA21X1 U243 ( .IN1(row_sel[1]), .IN2(n324), .IN3(n323), .Q(n32) );
  INVX0 U244 ( .INP(row_sel[0]), .ZN(n329) );
  AND2X1 U245 ( .IN1(\mat_i[3][2][0] ), .IN2(n292), .Q(\vector_out_i[2][0] )
         );
  AND2X1 U246 ( .IN1(\mat_i[3][2][1] ), .IN2(n292), .Q(\vector_out_i[2][1] )
         );
  AND2X1 U247 ( .IN1(\mat_i[3][2][2] ), .IN2(n292), .Q(\vector_out_i[2][2] )
         );
  AND2X1 U248 ( .IN1(\mat_i[3][2][3] ), .IN2(n292), .Q(\vector_out_i[2][3] )
         );
  AND2X1 U249 ( .IN1(\mat_i[3][2][4] ), .IN2(n292), .Q(\vector_out_i[2][4] )
         );
  AND2X1 U250 ( .IN1(\mat_i[3][2][5] ), .IN2(n292), .Q(\vector_out_i[2][5] )
         );
  AND2X1 U251 ( .IN1(\mat_i[3][2][6] ), .IN2(n292), .Q(\vector_out_i[2][6] )
         );
  AND2X1 U252 ( .IN1(\mat_i[3][2][7] ), .IN2(n292), .Q(\vector_out_i[2][7] )
         );
  AND2X1 U253 ( .IN1(\mat_i[3][2][8] ), .IN2(n292), .Q(\vector_out_i[2][8] )
         );
  AND2X1 U254 ( .IN1(\mat_i[3][2][9] ), .IN2(n292), .Q(\vector_out_i[2][9] )
         );
  AND2X1 U255 ( .IN1(\mat_i[3][2][10] ), .IN2(n292), .Q(\vector_out_i[2][10] )
         );
  AND2X1 U256 ( .IN1(\mat_i[3][2][11] ), .IN2(n292), .Q(\vector_out_i[2][11] )
         );
  AND2X1 U257 ( .IN1(n2), .IN2(n282), .Q(\vector_out_i[1][0] ) );
  AND2X1 U258 ( .IN1(n3), .IN2(n282), .Q(\vector_out_i[1][1] ) );
  AND2X1 U259 ( .IN1(n4), .IN2(n282), .Q(\vector_out_i[1][2] ) );
  AND2X1 U260 ( .IN1(n5), .IN2(n282), .Q(\vector_out_i[1][3] ) );
  AND2X1 U261 ( .IN1(n6), .IN2(n282), .Q(\vector_out_i[1][4] ) );
  AND2X1 U262 ( .IN1(n7), .IN2(n282), .Q(\vector_out_i[1][5] ) );
  AND2X1 U263 ( .IN1(n8), .IN2(n282), .Q(\vector_out_i[1][6] ) );
  AND2X1 U264 ( .IN1(n9), .IN2(n282), .Q(\vector_out_i[1][7] ) );
  AND2X1 U265 ( .IN1(n10), .IN2(n282), .Q(\vector_out_i[1][8] ) );
  AND2X1 U266 ( .IN1(n11), .IN2(n282), .Q(\vector_out_i[1][9] ) );
  AND2X1 U267 ( .IN1(n12), .IN2(n282), .Q(\vector_out_i[1][10] ) );
  AND2X1 U268 ( .IN1(n13), .IN2(n282), .Q(\vector_out_i[1][11] ) );
  AND2X1 U269 ( .IN1(\mat_r[3][3][0] ), .IN2(n291), .Q(\vector_out_r[3][0] )
         );
  AND2X1 U270 ( .IN1(\mat_r[3][3][1] ), .IN2(n291), .Q(\vector_out_r[3][1] )
         );
  AND2X1 U271 ( .IN1(\mat_r[3][3][2] ), .IN2(n291), .Q(\vector_out_r[3][2] )
         );
  AND2X1 U272 ( .IN1(\mat_r[3][3][3] ), .IN2(n291), .Q(\vector_out_r[3][3] )
         );
  AND2X1 U273 ( .IN1(\mat_r[3][3][4] ), .IN2(n291), .Q(\vector_out_r[3][4] )
         );
  AND2X1 U274 ( .IN1(\mat_r[3][3][5] ), .IN2(n291), .Q(\vector_out_r[3][5] )
         );
  AND2X1 U275 ( .IN1(\mat_r[3][3][6] ), .IN2(n291), .Q(\vector_out_r[3][6] )
         );
  AND2X1 U276 ( .IN1(\mat_r[3][3][7] ), .IN2(n291), .Q(\vector_out_r[3][7] )
         );
  AND2X1 U277 ( .IN1(\mat_r[3][3][8] ), .IN2(n291), .Q(\vector_out_r[3][8] )
         );
  AND2X1 U278 ( .IN1(\mat_r[3][3][9] ), .IN2(n291), .Q(\vector_out_r[3][9] )
         );
  AND2X1 U279 ( .IN1(\mat_r[3][3][10] ), .IN2(n291), .Q(\vector_out_r[3][10] )
         );
  AND2X1 U280 ( .IN1(\mat_r[3][3][11] ), .IN2(n291), .Q(\vector_out_r[3][11] )
         );
  AND2X1 U281 ( .IN1(n14), .IN2(n282), .Q(\vector_out_r[2][0] ) );
  AND2X1 U282 ( .IN1(n15), .IN2(n282), .Q(\vector_out_r[2][1] ) );
  AND2X1 U283 ( .IN1(n16), .IN2(n282), .Q(\vector_out_r[2][2] ) );
  AND2X1 U284 ( .IN1(n225), .IN2(n282), .Q(\vector_out_r[2][3] ) );
  AND2X1 U285 ( .IN1(n226), .IN2(n282), .Q(\vector_out_r[2][4] ) );
  AND2X1 U286 ( .IN1(n227), .IN2(n282), .Q(\vector_out_r[2][5] ) );
  AND2X1 U287 ( .IN1(n228), .IN2(n282), .Q(\vector_out_r[2][6] ) );
  AND2X1 U288 ( .IN1(n229), .IN2(n283), .Q(\vector_out_r[2][7] ) );
  AND2X1 U289 ( .IN1(n230), .IN2(n283), .Q(\vector_out_r[2][8] ) );
  AND2X1 U290 ( .IN1(n231), .IN2(n283), .Q(\vector_out_r[2][9] ) );
  AND2X1 U291 ( .IN1(n232), .IN2(n283), .Q(\vector_out_r[2][10] ) );
  AND2X1 U292 ( .IN1(n233), .IN2(n283), .Q(\vector_out_r[2][11] ) );
  MUX21X1 U293 ( .IN1(\mat_i[2][0][0] ), .IN2(\mat_i[3][0][0] ), .S(n288), .Q(
        n234) );
  AND2X1 U294 ( .IN1(\mat_i[1][0][0] ), .IN2(n286), .Q(n235) );
  MUX21X1 U295 ( .IN1(n235), .IN2(n234), .S(n285), .Q(\vector_out_i[0][0] ) );
  MUX21X1 U296 ( .IN1(\mat_i[2][0][1] ), .IN2(\mat_i[3][0][1] ), .S(n289), .Q(
        n236) );
  AND2X1 U297 ( .IN1(\mat_i[1][0][1] ), .IN2(n286), .Q(n237) );
  MUX21X1 U298 ( .IN1(n237), .IN2(n236), .S(n285), .Q(\vector_out_i[0][1] ) );
  MUX21X1 U299 ( .IN1(\mat_i[2][0][2] ), .IN2(\mat_i[3][0][2] ), .S(n289), .Q(
        n238) );
  AND2X1 U300 ( .IN1(\mat_i[1][0][2] ), .IN2(n286), .Q(n239) );
  MUX21X1 U301 ( .IN1(n239), .IN2(n238), .S(n285), .Q(\vector_out_i[0][2] ) );
  MUX21X1 U302 ( .IN1(\mat_i[2][0][3] ), .IN2(\mat_i[3][0][3] ), .S(n289), .Q(
        n240) );
  AND2X1 U303 ( .IN1(\mat_i[1][0][3] ), .IN2(n286), .Q(n241) );
  MUX21X1 U304 ( .IN1(n241), .IN2(n240), .S(n285), .Q(\vector_out_i[0][3] ) );
  MUX21X1 U305 ( .IN1(\mat_i[2][0][4] ), .IN2(\mat_i[3][0][4] ), .S(n289), .Q(
        n242) );
  AND2X1 U306 ( .IN1(\mat_i[1][0][4] ), .IN2(n286), .Q(n243) );
  MUX21X1 U307 ( .IN1(n243), .IN2(n242), .S(n285), .Q(\vector_out_i[0][4] ) );
  MUX21X1 U308 ( .IN1(\mat_i[2][0][5] ), .IN2(\mat_i[3][0][5] ), .S(n289), .Q(
        n244) );
  AND2X1 U309 ( .IN1(\mat_i[1][0][5] ), .IN2(n286), .Q(n245) );
  MUX21X1 U310 ( .IN1(n245), .IN2(n244), .S(n285), .Q(\vector_out_i[0][5] ) );
  MUX21X1 U311 ( .IN1(\mat_i[2][0][6] ), .IN2(\mat_i[3][0][6] ), .S(n289), .Q(
        n246) );
  AND2X1 U312 ( .IN1(\mat_i[1][0][6] ), .IN2(n286), .Q(n247) );
  MUX21X1 U313 ( .IN1(n247), .IN2(n246), .S(n285), .Q(\vector_out_i[0][6] ) );
  MUX21X1 U314 ( .IN1(\mat_i[2][0][7] ), .IN2(\mat_i[3][0][7] ), .S(n289), .Q(
        n248) );
  AND2X1 U315 ( .IN1(\mat_i[1][0][7] ), .IN2(n286), .Q(n249) );
  MUX21X1 U316 ( .IN1(n249), .IN2(n248), .S(n285), .Q(\vector_out_i[0][7] ) );
  MUX21X1 U317 ( .IN1(\mat_i[2][0][8] ), .IN2(\mat_i[3][0][8] ), .S(n289), .Q(
        n250) );
  AND2X1 U318 ( .IN1(\mat_i[1][0][8] ), .IN2(n286), .Q(n251) );
  MUX21X1 U319 ( .IN1(n251), .IN2(n250), .S(n285), .Q(\vector_out_i[0][8] ) );
  MUX21X1 U320 ( .IN1(\mat_i[2][0][9] ), .IN2(\mat_i[3][0][9] ), .S(n289), .Q(
        n252) );
  AND2X1 U321 ( .IN1(\mat_i[1][0][9] ), .IN2(n286), .Q(n253) );
  MUX21X1 U322 ( .IN1(n253), .IN2(n252), .S(n285), .Q(\vector_out_i[0][9] ) );
  MUX21X1 U323 ( .IN1(\mat_i[2][0][10] ), .IN2(\mat_i[3][0][10] ), .S(n289), 
        .Q(n254) );
  AND2X1 U324 ( .IN1(\mat_i[1][0][10] ), .IN2(n286), .Q(n255) );
  MUX21X1 U325 ( .IN1(n255), .IN2(n254), .S(n285), .Q(\vector_out_i[0][10] )
         );
  MUX21X1 U326 ( .IN1(\mat_i[2][0][11] ), .IN2(\mat_i[3][0][11] ), .S(n288), 
        .Q(n256) );
  AND2X1 U327 ( .IN1(\mat_i[1][0][11] ), .IN2(n287), .Q(n257) );
  MUX21X1 U328 ( .IN1(n257), .IN2(n256), .S(n285), .Q(\vector_out_i[0][11] )
         );
  MUX21X1 U329 ( .IN1(\mat_r[2][1][0] ), .IN2(\mat_r[3][1][0] ), .S(n289), .Q(
        n258) );
  AND2X1 U330 ( .IN1(\mat_r[1][1][0] ), .IN2(n287), .Q(n259) );
  MUX21X1 U331 ( .IN1(n259), .IN2(n258), .S(n284), .Q(\vector_out_r[1][0] ) );
  MUX21X1 U332 ( .IN1(\mat_r[2][1][1] ), .IN2(\mat_r[3][1][1] ), .S(n289), .Q(
        n260) );
  AND2X1 U333 ( .IN1(\mat_r[1][1][1] ), .IN2(n286), .Q(n261) );
  MUX21X1 U334 ( .IN1(n261), .IN2(n260), .S(n284), .Q(\vector_out_r[1][1] ) );
  MUX21X1 U335 ( .IN1(\mat_r[2][1][2] ), .IN2(\mat_r[3][1][2] ), .S(n289), .Q(
        n262) );
  AND2X1 U336 ( .IN1(\mat_r[1][1][2] ), .IN2(n287), .Q(n263) );
  MUX21X1 U337 ( .IN1(n263), .IN2(n262), .S(n284), .Q(\vector_out_r[1][2] ) );
  MUX21X1 U338 ( .IN1(\mat_r[2][1][3] ), .IN2(\mat_r[3][1][3] ), .S(n289), .Q(
        n264) );
  AND2X1 U339 ( .IN1(\mat_r[1][1][3] ), .IN2(n287), .Q(n265) );
  MUX21X1 U340 ( .IN1(n265), .IN2(n264), .S(n284), .Q(\vector_out_r[1][3] ) );
  MUX21X1 U341 ( .IN1(\mat_r[2][1][4] ), .IN2(\mat_r[3][1][4] ), .S(n289), .Q(
        n266) );
  AND2X1 U342 ( .IN1(\mat_r[1][1][4] ), .IN2(n287), .Q(n267) );
  MUX21X1 U343 ( .IN1(n267), .IN2(n266), .S(n284), .Q(\vector_out_r[1][4] ) );
  MUX21X1 U344 ( .IN1(\mat_r[2][1][5] ), .IN2(\mat_r[3][1][5] ), .S(n288), .Q(
        n268) );
  AND2X1 U345 ( .IN1(\mat_r[1][1][5] ), .IN2(n287), .Q(n269) );
  MUX21X1 U346 ( .IN1(n269), .IN2(n268), .S(n284), .Q(\vector_out_r[1][5] ) );
  MUX21X1 U347 ( .IN1(\mat_r[2][1][6] ), .IN2(\mat_r[3][1][6] ), .S(n289), .Q(
        n270) );
  AND2X1 U348 ( .IN1(\mat_r[1][1][6] ), .IN2(n287), .Q(n271) );
  MUX21X1 U349 ( .IN1(n271), .IN2(n270), .S(n284), .Q(\vector_out_r[1][6] ) );
  MUX21X1 U350 ( .IN1(\mat_r[2][1][7] ), .IN2(\mat_r[3][1][7] ), .S(n288), .Q(
        n272) );
  AND2X1 U351 ( .IN1(\mat_r[1][1][7] ), .IN2(n287), .Q(n273) );
  MUX21X1 U352 ( .IN1(n273), .IN2(n272), .S(n284), .Q(\vector_out_r[1][7] ) );
  MUX21X1 U353 ( .IN1(\mat_r[2][1][8] ), .IN2(\mat_r[3][1][8] ), .S(n288), .Q(
        n274) );
  AND2X1 U354 ( .IN1(\mat_r[1][1][8] ), .IN2(n287), .Q(n275) );
  MUX21X1 U355 ( .IN1(n275), .IN2(n274), .S(n284), .Q(\vector_out_r[1][8] ) );
  MUX21X1 U356 ( .IN1(\mat_r[2][1][9] ), .IN2(\mat_r[3][1][9] ), .S(n288), .Q(
        n276) );
  AND2X1 U357 ( .IN1(\mat_r[1][1][9] ), .IN2(n287), .Q(n277) );
  MUX21X1 U358 ( .IN1(n277), .IN2(n276), .S(n284), .Q(\vector_out_r[1][9] ) );
  MUX21X1 U359 ( .IN1(\mat_r[2][1][10] ), .IN2(\mat_r[3][1][10] ), .S(n289), 
        .Q(n278) );
  AND2X1 U360 ( .IN1(\mat_r[1][1][10] ), .IN2(n287), .Q(n279) );
  MUX21X1 U361 ( .IN1(n279), .IN2(n278), .S(n284), .Q(\vector_out_r[1][10] )
         );
  MUX21X1 U362 ( .IN1(\mat_r[2][1][11] ), .IN2(\mat_r[3][1][11] ), .S(n288), 
        .Q(n280) );
  AND2X1 U363 ( .IN1(\mat_r[1][1][11] ), .IN2(n287), .Q(n281) );
  MUX21X1 U364 ( .IN1(n281), .IN2(n280), .S(n284), .Q(\vector_out_r[1][11] )
         );
  MUX41X1 U365 ( .IN1(\mat_r[0][0][0] ), .IN3(\mat_r[2][0][0] ), .IN2(
        \mat_r[1][0][0] ), .IN4(\mat_r[3][0][0] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][0] ) );
  MUX41X1 U366 ( .IN1(\mat_r[0][0][1] ), .IN3(\mat_r[2][0][1] ), .IN2(
        \mat_r[1][0][1] ), .IN4(\mat_r[3][0][1] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][1] ) );
  MUX41X1 U367 ( .IN1(\mat_r[0][0][2] ), .IN3(\mat_r[2][0][2] ), .IN2(
        \mat_r[1][0][2] ), .IN4(\mat_r[3][0][2] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][2] ) );
  MUX41X1 U368 ( .IN1(\mat_r[0][0][3] ), .IN3(\mat_r[2][0][3] ), .IN2(
        \mat_r[1][0][3] ), .IN4(\mat_r[3][0][3] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][3] ) );
  MUX41X1 U369 ( .IN1(\mat_r[0][0][4] ), .IN3(\mat_r[2][0][4] ), .IN2(
        \mat_r[1][0][4] ), .IN4(\mat_r[3][0][4] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][4] ) );
  MUX41X1 U370 ( .IN1(\mat_r[0][0][5] ), .IN3(\mat_r[2][0][5] ), .IN2(
        \mat_r[1][0][5] ), .IN4(\mat_r[3][0][5] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][5] ) );
  MUX41X1 U371 ( .IN1(\mat_r[0][0][6] ), .IN3(\mat_r[2][0][6] ), .IN2(
        \mat_r[1][0][6] ), .IN4(\mat_r[3][0][6] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][6] ) );
  MUX41X1 U372 ( .IN1(\mat_r[0][0][7] ), .IN3(\mat_r[2][0][7] ), .IN2(
        \mat_r[1][0][7] ), .IN4(\mat_r[3][0][7] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][7] ) );
  MUX41X1 U373 ( .IN1(\mat_r[0][0][8] ), .IN3(\mat_r[2][0][8] ), .IN2(
        \mat_r[1][0][8] ), .IN4(\mat_r[3][0][8] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][8] ) );
  MUX41X1 U374 ( .IN1(\mat_r[0][0][9] ), .IN3(\mat_r[2][0][9] ), .IN2(
        \mat_r[1][0][9] ), .IN4(\mat_r[3][0][9] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][9] ) );
  MUX41X1 U375 ( .IN1(\mat_r[0][0][10] ), .IN3(\mat_r[2][0][10] ), .IN2(
        \mat_r[1][0][10] ), .IN4(\mat_r[3][0][10] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][10] ) );
  MUX41X1 U376 ( .IN1(\mat_r[0][0][11] ), .IN3(\mat_r[2][0][11] ), .IN2(
        \mat_r[1][0][11] ), .IN4(\mat_r[3][0][11] ), .S0(n283), .S1(n290), .Q(
        \vector_out_r[0][11] ) );
  MUX21X1 U377 ( .IN1(\mat_i[2][1][0] ), .IN2(\mat_i[3][1][0] ), .S(n288), .Q(
        n2) );
  MUX21X1 U378 ( .IN1(\mat_i[2][1][1] ), .IN2(\mat_i[3][1][1] ), .S(n288), .Q(
        n3) );
  MUX21X1 U379 ( .IN1(\mat_i[2][1][2] ), .IN2(\mat_i[3][1][2] ), .S(n288), .Q(
        n4) );
  MUX21X1 U380 ( .IN1(\mat_i[2][1][3] ), .IN2(\mat_i[3][1][3] ), .S(n288), .Q(
        n5) );
  MUX21X1 U381 ( .IN1(\mat_i[2][1][4] ), .IN2(\mat_i[3][1][4] ), .S(n288), .Q(
        n6) );
  MUX21X1 U382 ( .IN1(\mat_i[2][1][5] ), .IN2(\mat_i[3][1][5] ), .S(n288), .Q(
        n7) );
  MUX21X1 U383 ( .IN1(\mat_i[2][1][6] ), .IN2(\mat_i[3][1][6] ), .S(n288), .Q(
        n8) );
  MUX21X1 U384 ( .IN1(\mat_i[2][1][7] ), .IN2(\mat_i[3][1][7] ), .S(n288), .Q(
        n9) );
  MUX21X1 U385 ( .IN1(\mat_i[2][1][8] ), .IN2(\mat_i[3][1][8] ), .S(n288), .Q(
        n10) );
  MUX21X1 U386 ( .IN1(\mat_i[2][1][9] ), .IN2(\mat_i[3][1][9] ), .S(n288), .Q(
        n11) );
  MUX21X1 U387 ( .IN1(\mat_i[2][1][10] ), .IN2(\mat_i[3][1][10] ), .S(n287), 
        .Q(n12) );
  MUX21X1 U388 ( .IN1(\mat_i[2][1][11] ), .IN2(\mat_i[3][1][11] ), .S(n287), 
        .Q(n13) );
  MUX21X1 U389 ( .IN1(\mat_r[2][2][0] ), .IN2(\mat_r[3][2][0] ), .S(n287), .Q(
        n14) );
  MUX21X1 U390 ( .IN1(\mat_r[2][2][1] ), .IN2(\mat_r[3][2][1] ), .S(n288), .Q(
        n15) );
  MUX21X1 U391 ( .IN1(\mat_r[2][2][2] ), .IN2(\mat_r[3][2][2] ), .S(n287), .Q(
        n16) );
  MUX21X1 U392 ( .IN1(\mat_r[2][2][3] ), .IN2(\mat_r[3][2][3] ), .S(n287), .Q(
        n225) );
  MUX21X1 U393 ( .IN1(\mat_r[2][2][4] ), .IN2(\mat_r[3][2][4] ), .S(n287), .Q(
        n226) );
  MUX21X1 U394 ( .IN1(\mat_r[2][2][5] ), .IN2(\mat_r[3][2][5] ), .S(n287), .Q(
        n227) );
  MUX21X1 U395 ( .IN1(\mat_r[2][2][6] ), .IN2(\mat_r[3][2][6] ), .S(n287), .Q(
        n228) );
  MUX21X1 U396 ( .IN1(\mat_r[2][2][7] ), .IN2(\mat_r[3][2][7] ), .S(n287), .Q(
        n229) );
  MUX21X1 U397 ( .IN1(\mat_r[2][2][8] ), .IN2(\mat_r[3][2][8] ), .S(n287), .Q(
        n230) );
  MUX21X1 U398 ( .IN1(\mat_r[2][2][9] ), .IN2(\mat_r[3][2][9] ), .S(n287), .Q(
        n231) );
  MUX21X1 U399 ( .IN1(\mat_r[2][2][10] ), .IN2(\mat_r[3][2][10] ), .S(n287), 
        .Q(n232) );
  MUX21X1 U400 ( .IN1(\mat_r[2][2][11] ), .IN2(\mat_r[3][2][11] ), .S(n289), 
        .Q(n233) );
  INVX0 U401 ( .INP(n324), .ZN(n282) );
  INVX0 U402 ( .INP(n323), .ZN(n286) );
  INVX0 U403 ( .INP(n295), .ZN(n293) );
  INVX0 U404 ( .INP(n295), .ZN(n294) );
  INVX0 U405 ( .INP(n300), .ZN(n298) );
  INVX0 U406 ( .INP(n300), .ZN(n299) );
  INVX0 U407 ( .INP(n305), .ZN(n303) );
  INVX0 U408 ( .INP(n305), .ZN(n304) );
  INVX0 U409 ( .INP(n310), .ZN(n308) );
  INVX0 U410 ( .INP(n310), .ZN(n309) );
  INVX0 U411 ( .INP(n315), .ZN(n313) );
  INVX0 U412 ( .INP(n315), .ZN(n314) );
  INVX0 U413 ( .INP(n320), .ZN(n318) );
  INVX0 U414 ( .INP(n320), .ZN(n319) );
  INVX0 U415 ( .INP(N11), .ZN(n323) );
  INVX0 U416 ( .INP(N12), .ZN(n324) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_19_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n422), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U6 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U20 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n424), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n426), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n428), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n430), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(n25), .ZN(n422) );
  INVX0 U312 ( .INP(n3), .ZN(product[23]) );
  INVX0 U313 ( .INP(n55), .ZN(n428) );
  NBUFFX2 U314 ( .INP(a[1]), .Z(n409) );
  INVX0 U315 ( .INP(n463), .ZN(n431) );
  AND2X1 U316 ( .IN1(n409), .IN2(n411), .Q(n438) );
  INVX0 U317 ( .INP(n408), .ZN(n432) );
  INVX0 U318 ( .INP(n473), .ZN(n429) );
  INVX0 U319 ( .INP(n484), .ZN(n427) );
  INVX0 U320 ( .INP(n73), .ZN(n430) );
  INVX0 U321 ( .INP(n495), .ZN(n425) );
  INVX0 U322 ( .INP(n506), .ZN(n423) );
  INVX0 U323 ( .INP(n31), .ZN(n424) );
  INVX0 U324 ( .INP(n41), .ZN(n426) );
  AND2X1 U325 ( .IN1(n463), .IN2(n518), .Q(n436) );
  NBUFFX2 U326 ( .INP(a[3]), .Z(n413) );
  NBUFFX2 U327 ( .INP(b[0]), .Z(n408) );
  NBUFFX2 U328 ( .INP(a[5]), .Z(n415) );
  NBUFFX2 U329 ( .INP(a[3]), .Z(n412) );
  NBUFFX2 U330 ( .INP(a[5]), .Z(n414) );
  NBUFFX2 U331 ( .INP(a[7]), .Z(n416) );
  AND2X1 U332 ( .IN1(n484), .IN2(n522), .Q(n445) );
  AND2X1 U333 ( .IN1(n473), .IN2(n520), .Q(n442) );
  NBUFFX2 U334 ( .INP(a[9]), .Z(n418) );
  NBUFFX2 U335 ( .INP(a[11]), .Z(n420) );
  AND2X1 U336 ( .IN1(n495), .IN2(n524), .Q(n448) );
  AND2X1 U337 ( .IN1(n506), .IN2(n526), .Q(n451) );
  NBUFFX2 U338 ( .INP(a[7]), .Z(n417) );
  NBUFFX2 U339 ( .INP(a[9]), .Z(n419) );
  INVX0 U340 ( .INP(n411), .ZN(n410) );
  INVX0 U341 ( .INP(a[0]), .ZN(n411) );
  NOR2X0 U342 ( .IN1(n411), .IN2(n432), .QN(product[0]) );
  XNOR2X1 U343 ( .IN1(n433), .IN2(n434), .Q(n84) );
  NAND2X0 U344 ( .IN1(n434), .IN2(n433), .QN(n83) );
  AOI22X1 U345 ( .IN1(n435), .IN2(n431), .IN3(n436), .IN4(n437), .QN(n433) );
  OA21X1 U346 ( .IN1(n438), .IN2(n410), .IN3(n439), .Q(n434) );
  AO22X1 U347 ( .IN1(n440), .IN2(n431), .IN3(n436), .IN4(n435), .Q(n73) );
  XOR2X1 U348 ( .IN1(b[10]), .IN2(n412), .Q(n435) );
  AO22X1 U349 ( .IN1(n441), .IN2(n429), .IN3(n442), .IN4(n443), .Q(n55) );
  AO22X1 U350 ( .IN1(n444), .IN2(n427), .IN3(n445), .IN4(n446), .Q(n41) );
  AO22X1 U351 ( .IN1(n447), .IN2(n425), .IN3(n448), .IN4(n449), .Q(n31) );
  AO22X1 U352 ( .IN1(n450), .IN2(n423), .IN3(n451), .IN4(n452), .Q(n25) );
  AO22X1 U353 ( .IN1(n410), .IN2(n453), .IN3(n438), .IN4(n432), .Q(n224) );
  AO22X1 U354 ( .IN1(n410), .IN2(n454), .IN3(n438), .IN4(n453), .Q(n223) );
  XOR2X1 U355 ( .IN1(b[1]), .IN2(n409), .Q(n453) );
  AO22X1 U356 ( .IN1(n410), .IN2(n455), .IN3(n438), .IN4(n454), .Q(n222) );
  XOR2X1 U357 ( .IN1(b[2]), .IN2(n409), .Q(n454) );
  AO22X1 U358 ( .IN1(n410), .IN2(n456), .IN3(n438), .IN4(n455), .Q(n221) );
  XOR2X1 U359 ( .IN1(b[3]), .IN2(n409), .Q(n455) );
  AO22X1 U360 ( .IN1(n410), .IN2(n457), .IN3(n438), .IN4(n456), .Q(n220) );
  XOR2X1 U361 ( .IN1(b[4]), .IN2(n409), .Q(n456) );
  AO22X1 U362 ( .IN1(n410), .IN2(n458), .IN3(n438), .IN4(n457), .Q(n219) );
  XOR2X1 U363 ( .IN1(b[5]), .IN2(n409), .Q(n457) );
  AO22X1 U364 ( .IN1(n410), .IN2(n459), .IN3(n438), .IN4(n458), .Q(n218) );
  XOR2X1 U365 ( .IN1(b[6]), .IN2(n409), .Q(n458) );
  AO22X1 U366 ( .IN1(n410), .IN2(n460), .IN3(n438), .IN4(n459), .Q(n217) );
  XOR2X1 U367 ( .IN1(b[7]), .IN2(n409), .Q(n459) );
  AO22X1 U368 ( .IN1(n410), .IN2(n461), .IN3(n438), .IN4(n460), .Q(n216) );
  XOR2X1 U369 ( .IN1(b[8]), .IN2(n409), .Q(n460) );
  AO22X1 U370 ( .IN1(n410), .IN2(n462), .IN3(n438), .IN4(n461), .Q(n215) );
  XOR2X1 U371 ( .IN1(b[9]), .IN2(n409), .Q(n461) );
  AO22X1 U372 ( .IN1(n410), .IN2(n439), .IN3(n438), .IN4(n462), .Q(n214) );
  XOR2X1 U373 ( .IN1(b[10]), .IN2(n409), .Q(n462) );
  XOR2X1 U374 ( .IN1(b[11]), .IN2(n409), .Q(n439) );
  NOR2X0 U375 ( .IN1(n463), .IN2(n432), .QN(n212) );
  AO22X1 U376 ( .IN1(n464), .IN2(n431), .IN3(n436), .IN4(n465), .Q(n211) );
  XOR2X1 U377 ( .IN1(n408), .IN2(n412), .Q(n465) );
  AO22X1 U378 ( .IN1(n466), .IN2(n431), .IN3(n436), .IN4(n464), .Q(n210) );
  XOR2X1 U379 ( .IN1(b[1]), .IN2(n412), .Q(n464) );
  AO22X1 U380 ( .IN1(n467), .IN2(n431), .IN3(n436), .IN4(n466), .Q(n209) );
  XOR2X1 U381 ( .IN1(b[2]), .IN2(n412), .Q(n466) );
  AO22X1 U382 ( .IN1(n468), .IN2(n431), .IN3(n436), .IN4(n467), .Q(n208) );
  XOR2X1 U383 ( .IN1(b[3]), .IN2(n412), .Q(n467) );
  AO22X1 U384 ( .IN1(n469), .IN2(n431), .IN3(n436), .IN4(n468), .Q(n207) );
  XOR2X1 U385 ( .IN1(b[4]), .IN2(n412), .Q(n468) );
  AO22X1 U386 ( .IN1(n470), .IN2(n431), .IN3(n436), .IN4(n469), .Q(n206) );
  XOR2X1 U387 ( .IN1(b[5]), .IN2(n412), .Q(n469) );
  AO22X1 U388 ( .IN1(n471), .IN2(n431), .IN3(n436), .IN4(n470), .Q(n205) );
  XOR2X1 U389 ( .IN1(b[6]), .IN2(n412), .Q(n470) );
  AO22X1 U390 ( .IN1(n472), .IN2(n431), .IN3(n436), .IN4(n471), .Q(n204) );
  XOR2X1 U391 ( .IN1(b[7]), .IN2(n412), .Q(n471) );
  AO22X1 U392 ( .IN1(n437), .IN2(n431), .IN3(n436), .IN4(n472), .Q(n203) );
  XOR2X1 U393 ( .IN1(b[8]), .IN2(n412), .Q(n472) );
  XOR2X1 U394 ( .IN1(b[9]), .IN2(n412), .Q(n437) );
  OAI21X1 U395 ( .IN1(n431), .IN2(n436), .IN3(n440), .QN(n201) );
  XOR2X1 U396 ( .IN1(b[11]), .IN2(n412), .Q(n440) );
  NOR2X0 U397 ( .IN1(n473), .IN2(n432), .QN(n200) );
  AO22X1 U398 ( .IN1(n474), .IN2(n429), .IN3(n442), .IN4(n475), .Q(n199) );
  XOR2X1 U399 ( .IN1(n408), .IN2(n414), .Q(n475) );
  AO22X1 U400 ( .IN1(n476), .IN2(n429), .IN3(n442), .IN4(n474), .Q(n198) );
  XOR2X1 U401 ( .IN1(b[1]), .IN2(n414), .Q(n474) );
  AO22X1 U402 ( .IN1(n477), .IN2(n429), .IN3(n442), .IN4(n476), .Q(n197) );
  XOR2X1 U403 ( .IN1(b[2]), .IN2(n414), .Q(n476) );
  AO22X1 U404 ( .IN1(n478), .IN2(n429), .IN3(n442), .IN4(n477), .Q(n196) );
  XOR2X1 U405 ( .IN1(b[3]), .IN2(n414), .Q(n477) );
  AO22X1 U406 ( .IN1(n479), .IN2(n429), .IN3(n442), .IN4(n478), .Q(n195) );
  XOR2X1 U407 ( .IN1(b[4]), .IN2(n414), .Q(n478) );
  AO22X1 U408 ( .IN1(n480), .IN2(n429), .IN3(n442), .IN4(n479), .Q(n194) );
  XOR2X1 U409 ( .IN1(b[5]), .IN2(n414), .Q(n479) );
  AO22X1 U410 ( .IN1(n481), .IN2(n429), .IN3(n442), .IN4(n480), .Q(n193) );
  XOR2X1 U411 ( .IN1(b[6]), .IN2(n414), .Q(n480) );
  AO22X1 U412 ( .IN1(n482), .IN2(n429), .IN3(n442), .IN4(n481), .Q(n192) );
  XOR2X1 U413 ( .IN1(b[7]), .IN2(n414), .Q(n481) );
  AO22X1 U414 ( .IN1(n483), .IN2(n429), .IN3(n442), .IN4(n482), .Q(n191) );
  XOR2X1 U415 ( .IN1(b[8]), .IN2(n414), .Q(n482) );
  AO22X1 U416 ( .IN1(n443), .IN2(n429), .IN3(n442), .IN4(n483), .Q(n190) );
  XOR2X1 U417 ( .IN1(b[9]), .IN2(n414), .Q(n483) );
  XOR2X1 U418 ( .IN1(b[10]), .IN2(n414), .Q(n443) );
  OAI21X1 U419 ( .IN1(n429), .IN2(n442), .IN3(n441), .QN(n189) );
  XOR2X1 U420 ( .IN1(b[11]), .IN2(n414), .Q(n441) );
  NOR2X0 U421 ( .IN1(n484), .IN2(n432), .QN(n188) );
  AO22X1 U422 ( .IN1(n485), .IN2(n427), .IN3(n445), .IN4(n486), .Q(n187) );
  XOR2X1 U423 ( .IN1(n408), .IN2(n416), .Q(n486) );
  AO22X1 U424 ( .IN1(n487), .IN2(n427), .IN3(n445), .IN4(n485), .Q(n186) );
  XOR2X1 U425 ( .IN1(b[1]), .IN2(n416), .Q(n485) );
  AO22X1 U426 ( .IN1(n488), .IN2(n427), .IN3(n445), .IN4(n487), .Q(n185) );
  XOR2X1 U427 ( .IN1(b[2]), .IN2(n416), .Q(n487) );
  AO22X1 U428 ( .IN1(n489), .IN2(n427), .IN3(n445), .IN4(n488), .Q(n184) );
  XOR2X1 U429 ( .IN1(b[3]), .IN2(n416), .Q(n488) );
  AO22X1 U430 ( .IN1(n490), .IN2(n427), .IN3(n445), .IN4(n489), .Q(n183) );
  XOR2X1 U431 ( .IN1(b[4]), .IN2(n416), .Q(n489) );
  AO22X1 U432 ( .IN1(n491), .IN2(n427), .IN3(n445), .IN4(n490), .Q(n182) );
  XOR2X1 U433 ( .IN1(b[5]), .IN2(n416), .Q(n490) );
  AO22X1 U434 ( .IN1(n492), .IN2(n427), .IN3(n445), .IN4(n491), .Q(n181) );
  XOR2X1 U435 ( .IN1(b[6]), .IN2(n416), .Q(n491) );
  AO22X1 U436 ( .IN1(n493), .IN2(n427), .IN3(n445), .IN4(n492), .Q(n180) );
  XOR2X1 U437 ( .IN1(b[7]), .IN2(n416), .Q(n492) );
  AO22X1 U438 ( .IN1(n494), .IN2(n427), .IN3(n445), .IN4(n493), .Q(n179) );
  XOR2X1 U439 ( .IN1(b[8]), .IN2(n416), .Q(n493) );
  AO22X1 U440 ( .IN1(n446), .IN2(n427), .IN3(n445), .IN4(n494), .Q(n178) );
  XOR2X1 U441 ( .IN1(b[9]), .IN2(n416), .Q(n494) );
  XOR2X1 U442 ( .IN1(b[10]), .IN2(n416), .Q(n446) );
  OAI21X1 U443 ( .IN1(n427), .IN2(n445), .IN3(n444), .QN(n177) );
  XOR2X1 U444 ( .IN1(b[11]), .IN2(n416), .Q(n444) );
  NOR2X0 U445 ( .IN1(n495), .IN2(n432), .QN(n176) );
  AO22X1 U446 ( .IN1(n496), .IN2(n425), .IN3(n448), .IN4(n497), .Q(n175) );
  XOR2X1 U447 ( .IN1(n408), .IN2(n418), .Q(n497) );
  AO22X1 U448 ( .IN1(n498), .IN2(n425), .IN3(n448), .IN4(n496), .Q(n174) );
  XOR2X1 U449 ( .IN1(b[1]), .IN2(n418), .Q(n496) );
  AO22X1 U450 ( .IN1(n499), .IN2(n425), .IN3(n448), .IN4(n498), .Q(n173) );
  XOR2X1 U451 ( .IN1(b[2]), .IN2(n418), .Q(n498) );
  AO22X1 U452 ( .IN1(n500), .IN2(n425), .IN3(n448), .IN4(n499), .Q(n172) );
  XOR2X1 U453 ( .IN1(b[3]), .IN2(n418), .Q(n499) );
  AO22X1 U454 ( .IN1(n501), .IN2(n425), .IN3(n448), .IN4(n500), .Q(n171) );
  XOR2X1 U455 ( .IN1(b[4]), .IN2(n418), .Q(n500) );
  AO22X1 U456 ( .IN1(n502), .IN2(n425), .IN3(n448), .IN4(n501), .Q(n170) );
  XOR2X1 U457 ( .IN1(b[5]), .IN2(n418), .Q(n501) );
  AO22X1 U458 ( .IN1(n503), .IN2(n425), .IN3(n448), .IN4(n502), .Q(n169) );
  XOR2X1 U459 ( .IN1(b[6]), .IN2(n418), .Q(n502) );
  AO22X1 U460 ( .IN1(n504), .IN2(n425), .IN3(n448), .IN4(n503), .Q(n168) );
  XOR2X1 U461 ( .IN1(b[7]), .IN2(n418), .Q(n503) );
  AO22X1 U462 ( .IN1(n505), .IN2(n425), .IN3(n448), .IN4(n504), .Q(n167) );
  XOR2X1 U463 ( .IN1(b[8]), .IN2(n418), .Q(n504) );
  AO22X1 U464 ( .IN1(n449), .IN2(n425), .IN3(n448), .IN4(n505), .Q(n166) );
  XOR2X1 U465 ( .IN1(b[9]), .IN2(n418), .Q(n505) );
  XOR2X1 U466 ( .IN1(b[10]), .IN2(n418), .Q(n449) );
  OAI21X1 U467 ( .IN1(n425), .IN2(n448), .IN3(n447), .QN(n165) );
  XOR2X1 U468 ( .IN1(b[11]), .IN2(n418), .Q(n447) );
  NOR2X0 U469 ( .IN1(n506), .IN2(n432), .QN(n164) );
  AO22X1 U470 ( .IN1(n507), .IN2(n423), .IN3(n451), .IN4(n508), .Q(n163) );
  XOR2X1 U471 ( .IN1(n408), .IN2(n420), .Q(n508) );
  AO22X1 U472 ( .IN1(n509), .IN2(n423), .IN3(n451), .IN4(n507), .Q(n162) );
  XOR2X1 U473 ( .IN1(b[1]), .IN2(n420), .Q(n507) );
  AO22X1 U474 ( .IN1(n510), .IN2(n423), .IN3(n451), .IN4(n509), .Q(n161) );
  XOR2X1 U475 ( .IN1(b[2]), .IN2(n420), .Q(n509) );
  AO22X1 U476 ( .IN1(n511), .IN2(n423), .IN3(n451), .IN4(n510), .Q(n160) );
  XOR2X1 U477 ( .IN1(b[3]), .IN2(n420), .Q(n510) );
  AO22X1 U478 ( .IN1(n512), .IN2(n423), .IN3(n451), .IN4(n511), .Q(n159) );
  XOR2X1 U479 ( .IN1(b[4]), .IN2(n420), .Q(n511) );
  AO22X1 U480 ( .IN1(n513), .IN2(n423), .IN3(n451), .IN4(n512), .Q(n158) );
  XOR2X1 U481 ( .IN1(b[5]), .IN2(n420), .Q(n512) );
  AO22X1 U482 ( .IN1(n514), .IN2(n423), .IN3(n451), .IN4(n513), .Q(n157) );
  XOR2X1 U483 ( .IN1(b[6]), .IN2(n420), .Q(n513) );
  AO22X1 U484 ( .IN1(n515), .IN2(n423), .IN3(n451), .IN4(n514), .Q(n156) );
  XOR2X1 U485 ( .IN1(b[7]), .IN2(n420), .Q(n514) );
  AO22X1 U486 ( .IN1(n516), .IN2(n423), .IN3(n451), .IN4(n515), .Q(n155) );
  XOR2X1 U487 ( .IN1(b[8]), .IN2(n420), .Q(n515) );
  AO22X1 U488 ( .IN1(n452), .IN2(n423), .IN3(n451), .IN4(n516), .Q(n154) );
  XOR2X1 U489 ( .IN1(b[9]), .IN2(n420), .Q(n516) );
  XOR2X1 U490 ( .IN1(b[10]), .IN2(n420), .Q(n452) );
  OAI21X1 U491 ( .IN1(n423), .IN2(n451), .IN3(n450), .QN(n153) );
  XOR2X1 U492 ( .IN1(b[11]), .IN2(n420), .Q(n450) );
  AO21X1 U493 ( .IN1(n409), .IN2(n432), .IN3(n438), .Q(n152) );
  AO22X1 U494 ( .IN1(n517), .IN2(n413), .IN3(n436), .IN4(n413), .Q(n151) );
  XOR2X1 U495 ( .IN1(n412), .IN2(a[2]), .Q(n518) );
  NOR2X0 U496 ( .IN1(n408), .IN2(n463), .QN(n517) );
  XNOR2X1 U497 ( .IN1(a[2]), .IN2(n409), .Q(n463) );
  AO22X1 U498 ( .IN1(n519), .IN2(n415), .IN3(n442), .IN4(n415), .Q(n150) );
  XOR2X1 U499 ( .IN1(n414), .IN2(a[4]), .Q(n520) );
  NOR2X0 U500 ( .IN1(n408), .IN2(n473), .QN(n519) );
  XNOR2X1 U501 ( .IN1(a[4]), .IN2(n412), .Q(n473) );
  AO22X1 U502 ( .IN1(n521), .IN2(n417), .IN3(n445), .IN4(n417), .Q(n149) );
  XOR2X1 U503 ( .IN1(n416), .IN2(a[6]), .Q(n522) );
  NOR2X0 U504 ( .IN1(n408), .IN2(n484), .QN(n521) );
  XNOR2X1 U505 ( .IN1(a[6]), .IN2(n414), .Q(n484) );
  AO22X1 U506 ( .IN1(n523), .IN2(n419), .IN3(n448), .IN4(n419), .Q(n148) );
  XOR2X1 U507 ( .IN1(n418), .IN2(a[8]), .Q(n524) );
  NOR2X0 U508 ( .IN1(n408), .IN2(n495), .QN(n523) );
  XNOR2X1 U509 ( .IN1(a[8]), .IN2(n416), .Q(n495) );
  AO22X1 U510 ( .IN1(n525), .IN2(a[11]), .IN3(n451), .IN4(n420), .Q(n147) );
  XOR2X1 U511 ( .IN1(n420), .IN2(a[10]), .Q(n526) );
  NOR2X0 U512 ( .IN1(n408), .IN2(n506), .QN(n525) );
  XNOR2X1 U513 ( .IN1(a[10]), .IN2(n418), .Q(n506) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_19 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_19_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_18_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n425), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U6 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U20 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n424), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n423), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n422), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n421), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(n25), .ZN(n425) );
  INVX0 U312 ( .INP(n3), .ZN(product[23]) );
  INVX0 U313 ( .INP(n55), .ZN(n422) );
  INVX0 U314 ( .INP(n462), .ZN(n431) );
  INVX0 U315 ( .INP(n408), .ZN(n426) );
  AND2X1 U316 ( .IN1(a[1]), .IN2(n410), .Q(n437) );
  INVX0 U317 ( .INP(n472), .ZN(n430) );
  INVX0 U318 ( .INP(n483), .ZN(n429) );
  INVX0 U319 ( .INP(n494), .ZN(n428) );
  INVX0 U320 ( .INP(n505), .ZN(n427) );
  INVX0 U321 ( .INP(n73), .ZN(n421) );
  INVX0 U322 ( .INP(n31), .ZN(n424) );
  INVX0 U323 ( .INP(n41), .ZN(n423) );
  NBUFFX2 U324 ( .INP(b[0]), .Z(n408) );
  AND2X1 U325 ( .IN1(n462), .IN2(n517), .Q(n435) );
  NBUFFX2 U326 ( .INP(a[3]), .Z(n412) );
  NBUFFX2 U327 ( .INP(a[3]), .Z(n411) );
  NBUFFX2 U328 ( .INP(a[5]), .Z(n413) );
  NBUFFX2 U329 ( .INP(a[7]), .Z(n415) );
  AND2X1 U330 ( .IN1(n483), .IN2(n521), .Q(n444) );
  AND2X1 U331 ( .IN1(n472), .IN2(n519), .Q(n441) );
  NBUFFX2 U332 ( .INP(a[5]), .Z(n414) );
  NBUFFX2 U333 ( .INP(a[9]), .Z(n417) );
  NBUFFX2 U334 ( .INP(a[11]), .Z(n419) );
  AND2X1 U335 ( .IN1(n494), .IN2(n523), .Q(n447) );
  AND2X1 U336 ( .IN1(n505), .IN2(n525), .Q(n450) );
  NBUFFX2 U337 ( .INP(a[7]), .Z(n416) );
  NBUFFX2 U338 ( .INP(a[9]), .Z(n418) );
  INVX0 U339 ( .INP(n410), .ZN(n409) );
  INVX0 U340 ( .INP(a[0]), .ZN(n410) );
  NOR2X0 U341 ( .IN1(n410), .IN2(n426), .QN(product[0]) );
  XNOR2X1 U342 ( .IN1(n432), .IN2(n433), .Q(n84) );
  NAND2X0 U343 ( .IN1(n433), .IN2(n432), .QN(n83) );
  AOI22X1 U344 ( .IN1(n434), .IN2(n431), .IN3(n435), .IN4(n436), .QN(n432) );
  OA21X1 U345 ( .IN1(n437), .IN2(n409), .IN3(n438), .Q(n433) );
  AO22X1 U346 ( .IN1(n439), .IN2(n431), .IN3(n435), .IN4(n434), .Q(n73) );
  XOR2X1 U347 ( .IN1(b[10]), .IN2(n411), .Q(n434) );
  AO22X1 U348 ( .IN1(n440), .IN2(n430), .IN3(n441), .IN4(n442), .Q(n55) );
  AO22X1 U349 ( .IN1(n443), .IN2(n429), .IN3(n444), .IN4(n445), .Q(n41) );
  AO22X1 U350 ( .IN1(n446), .IN2(n428), .IN3(n447), .IN4(n448), .Q(n31) );
  AO22X1 U351 ( .IN1(n449), .IN2(n427), .IN3(n450), .IN4(n451), .Q(n25) );
  AO22X1 U352 ( .IN1(n409), .IN2(n452), .IN3(n437), .IN4(n426), .Q(n224) );
  AO22X1 U353 ( .IN1(n409), .IN2(n453), .IN3(n437), .IN4(n452), .Q(n223) );
  XOR2X1 U354 ( .IN1(b[1]), .IN2(a[1]), .Q(n452) );
  AO22X1 U355 ( .IN1(n409), .IN2(n454), .IN3(n437), .IN4(n453), .Q(n222) );
  XOR2X1 U356 ( .IN1(b[2]), .IN2(a[1]), .Q(n453) );
  AO22X1 U357 ( .IN1(n409), .IN2(n455), .IN3(n437), .IN4(n454), .Q(n221) );
  XOR2X1 U358 ( .IN1(b[3]), .IN2(a[1]), .Q(n454) );
  AO22X1 U359 ( .IN1(n409), .IN2(n456), .IN3(n437), .IN4(n455), .Q(n220) );
  XOR2X1 U360 ( .IN1(b[4]), .IN2(a[1]), .Q(n455) );
  AO22X1 U361 ( .IN1(n409), .IN2(n457), .IN3(n437), .IN4(n456), .Q(n219) );
  XOR2X1 U362 ( .IN1(b[5]), .IN2(a[1]), .Q(n456) );
  AO22X1 U363 ( .IN1(n409), .IN2(n458), .IN3(n437), .IN4(n457), .Q(n218) );
  XOR2X1 U364 ( .IN1(b[6]), .IN2(a[1]), .Q(n457) );
  AO22X1 U365 ( .IN1(n409), .IN2(n459), .IN3(n437), .IN4(n458), .Q(n217) );
  XOR2X1 U366 ( .IN1(b[7]), .IN2(a[1]), .Q(n458) );
  AO22X1 U367 ( .IN1(n409), .IN2(n460), .IN3(n437), .IN4(n459), .Q(n216) );
  XOR2X1 U368 ( .IN1(b[8]), .IN2(a[1]), .Q(n459) );
  AO22X1 U369 ( .IN1(n409), .IN2(n461), .IN3(n437), .IN4(n460), .Q(n215) );
  XOR2X1 U370 ( .IN1(b[9]), .IN2(a[1]), .Q(n460) );
  AO22X1 U371 ( .IN1(n409), .IN2(n438), .IN3(n437), .IN4(n461), .Q(n214) );
  XOR2X1 U372 ( .IN1(b[10]), .IN2(a[1]), .Q(n461) );
  XOR2X1 U373 ( .IN1(b[11]), .IN2(a[1]), .Q(n438) );
  NOR2X0 U374 ( .IN1(n462), .IN2(n426), .QN(n212) );
  AO22X1 U375 ( .IN1(n463), .IN2(n431), .IN3(n435), .IN4(n464), .Q(n211) );
  XOR2X1 U376 ( .IN1(n408), .IN2(n411), .Q(n464) );
  AO22X1 U377 ( .IN1(n465), .IN2(n431), .IN3(n435), .IN4(n463), .Q(n210) );
  XOR2X1 U378 ( .IN1(b[1]), .IN2(n411), .Q(n463) );
  AO22X1 U379 ( .IN1(n466), .IN2(n431), .IN3(n435), .IN4(n465), .Q(n209) );
  XOR2X1 U380 ( .IN1(b[2]), .IN2(n411), .Q(n465) );
  AO22X1 U381 ( .IN1(n467), .IN2(n431), .IN3(n435), .IN4(n466), .Q(n208) );
  XOR2X1 U382 ( .IN1(b[3]), .IN2(n411), .Q(n466) );
  AO22X1 U383 ( .IN1(n468), .IN2(n431), .IN3(n435), .IN4(n467), .Q(n207) );
  XOR2X1 U384 ( .IN1(b[4]), .IN2(n411), .Q(n467) );
  AO22X1 U385 ( .IN1(n469), .IN2(n431), .IN3(n435), .IN4(n468), .Q(n206) );
  XOR2X1 U386 ( .IN1(b[5]), .IN2(n411), .Q(n468) );
  AO22X1 U387 ( .IN1(n470), .IN2(n431), .IN3(n435), .IN4(n469), .Q(n205) );
  XOR2X1 U388 ( .IN1(b[6]), .IN2(n411), .Q(n469) );
  AO22X1 U389 ( .IN1(n471), .IN2(n431), .IN3(n435), .IN4(n470), .Q(n204) );
  XOR2X1 U390 ( .IN1(b[7]), .IN2(n411), .Q(n470) );
  AO22X1 U391 ( .IN1(n436), .IN2(n431), .IN3(n435), .IN4(n471), .Q(n203) );
  XOR2X1 U392 ( .IN1(b[8]), .IN2(n411), .Q(n471) );
  XOR2X1 U393 ( .IN1(b[9]), .IN2(n411), .Q(n436) );
  OAI21X1 U394 ( .IN1(n431), .IN2(n435), .IN3(n439), .QN(n201) );
  XOR2X1 U395 ( .IN1(b[11]), .IN2(n411), .Q(n439) );
  NOR2X0 U396 ( .IN1(n472), .IN2(n426), .QN(n200) );
  AO22X1 U397 ( .IN1(n473), .IN2(n430), .IN3(n441), .IN4(n474), .Q(n199) );
  XOR2X1 U398 ( .IN1(n408), .IN2(n413), .Q(n474) );
  AO22X1 U399 ( .IN1(n475), .IN2(n430), .IN3(n441), .IN4(n473), .Q(n198) );
  XOR2X1 U400 ( .IN1(b[1]), .IN2(n413), .Q(n473) );
  AO22X1 U401 ( .IN1(n476), .IN2(n430), .IN3(n441), .IN4(n475), .Q(n197) );
  XOR2X1 U402 ( .IN1(b[2]), .IN2(n413), .Q(n475) );
  AO22X1 U403 ( .IN1(n477), .IN2(n430), .IN3(n441), .IN4(n476), .Q(n196) );
  XOR2X1 U404 ( .IN1(b[3]), .IN2(n413), .Q(n476) );
  AO22X1 U405 ( .IN1(n478), .IN2(n430), .IN3(n441), .IN4(n477), .Q(n195) );
  XOR2X1 U406 ( .IN1(b[4]), .IN2(n413), .Q(n477) );
  AO22X1 U407 ( .IN1(n479), .IN2(n430), .IN3(n441), .IN4(n478), .Q(n194) );
  XOR2X1 U408 ( .IN1(b[5]), .IN2(n413), .Q(n478) );
  AO22X1 U409 ( .IN1(n480), .IN2(n430), .IN3(n441), .IN4(n479), .Q(n193) );
  XOR2X1 U410 ( .IN1(b[6]), .IN2(n413), .Q(n479) );
  AO22X1 U411 ( .IN1(n481), .IN2(n430), .IN3(n441), .IN4(n480), .Q(n192) );
  XOR2X1 U412 ( .IN1(b[7]), .IN2(n413), .Q(n480) );
  AO22X1 U413 ( .IN1(n482), .IN2(n430), .IN3(n441), .IN4(n481), .Q(n191) );
  XOR2X1 U414 ( .IN1(b[8]), .IN2(n413), .Q(n481) );
  AO22X1 U415 ( .IN1(n442), .IN2(n430), .IN3(n441), .IN4(n482), .Q(n190) );
  XOR2X1 U416 ( .IN1(b[9]), .IN2(n413), .Q(n482) );
  XOR2X1 U417 ( .IN1(b[10]), .IN2(n413), .Q(n442) );
  OAI21X1 U418 ( .IN1(n430), .IN2(n441), .IN3(n440), .QN(n189) );
  XOR2X1 U419 ( .IN1(b[11]), .IN2(n413), .Q(n440) );
  NOR2X0 U420 ( .IN1(n483), .IN2(n426), .QN(n188) );
  AO22X1 U421 ( .IN1(n484), .IN2(n429), .IN3(n444), .IN4(n485), .Q(n187) );
  XOR2X1 U422 ( .IN1(n408), .IN2(n415), .Q(n485) );
  AO22X1 U423 ( .IN1(n486), .IN2(n429), .IN3(n444), .IN4(n484), .Q(n186) );
  XOR2X1 U424 ( .IN1(b[1]), .IN2(n415), .Q(n484) );
  AO22X1 U425 ( .IN1(n487), .IN2(n429), .IN3(n444), .IN4(n486), .Q(n185) );
  XOR2X1 U426 ( .IN1(b[2]), .IN2(n415), .Q(n486) );
  AO22X1 U427 ( .IN1(n488), .IN2(n429), .IN3(n444), .IN4(n487), .Q(n184) );
  XOR2X1 U428 ( .IN1(b[3]), .IN2(n415), .Q(n487) );
  AO22X1 U429 ( .IN1(n489), .IN2(n429), .IN3(n444), .IN4(n488), .Q(n183) );
  XOR2X1 U430 ( .IN1(b[4]), .IN2(n415), .Q(n488) );
  AO22X1 U431 ( .IN1(n490), .IN2(n429), .IN3(n444), .IN4(n489), .Q(n182) );
  XOR2X1 U432 ( .IN1(b[5]), .IN2(n415), .Q(n489) );
  AO22X1 U433 ( .IN1(n491), .IN2(n429), .IN3(n444), .IN4(n490), .Q(n181) );
  XOR2X1 U434 ( .IN1(b[6]), .IN2(n415), .Q(n490) );
  AO22X1 U435 ( .IN1(n492), .IN2(n429), .IN3(n444), .IN4(n491), .Q(n180) );
  XOR2X1 U436 ( .IN1(b[7]), .IN2(n415), .Q(n491) );
  AO22X1 U437 ( .IN1(n493), .IN2(n429), .IN3(n444), .IN4(n492), .Q(n179) );
  XOR2X1 U438 ( .IN1(b[8]), .IN2(n415), .Q(n492) );
  AO22X1 U439 ( .IN1(n445), .IN2(n429), .IN3(n444), .IN4(n493), .Q(n178) );
  XOR2X1 U440 ( .IN1(b[9]), .IN2(n415), .Q(n493) );
  XOR2X1 U441 ( .IN1(b[10]), .IN2(n415), .Q(n445) );
  OAI21X1 U442 ( .IN1(n429), .IN2(n444), .IN3(n443), .QN(n177) );
  XOR2X1 U443 ( .IN1(b[11]), .IN2(n415), .Q(n443) );
  NOR2X0 U444 ( .IN1(n494), .IN2(n426), .QN(n176) );
  AO22X1 U445 ( .IN1(n495), .IN2(n428), .IN3(n447), .IN4(n496), .Q(n175) );
  XOR2X1 U446 ( .IN1(n408), .IN2(n417), .Q(n496) );
  AO22X1 U447 ( .IN1(n497), .IN2(n428), .IN3(n447), .IN4(n495), .Q(n174) );
  XOR2X1 U448 ( .IN1(b[1]), .IN2(n417), .Q(n495) );
  AO22X1 U449 ( .IN1(n498), .IN2(n428), .IN3(n447), .IN4(n497), .Q(n173) );
  XOR2X1 U450 ( .IN1(b[2]), .IN2(n417), .Q(n497) );
  AO22X1 U451 ( .IN1(n499), .IN2(n428), .IN3(n447), .IN4(n498), .Q(n172) );
  XOR2X1 U452 ( .IN1(b[3]), .IN2(n417), .Q(n498) );
  AO22X1 U453 ( .IN1(n500), .IN2(n428), .IN3(n447), .IN4(n499), .Q(n171) );
  XOR2X1 U454 ( .IN1(b[4]), .IN2(n417), .Q(n499) );
  AO22X1 U455 ( .IN1(n501), .IN2(n428), .IN3(n447), .IN4(n500), .Q(n170) );
  XOR2X1 U456 ( .IN1(b[5]), .IN2(n417), .Q(n500) );
  AO22X1 U457 ( .IN1(n502), .IN2(n428), .IN3(n447), .IN4(n501), .Q(n169) );
  XOR2X1 U458 ( .IN1(b[6]), .IN2(n417), .Q(n501) );
  AO22X1 U459 ( .IN1(n503), .IN2(n428), .IN3(n447), .IN4(n502), .Q(n168) );
  XOR2X1 U460 ( .IN1(b[7]), .IN2(n417), .Q(n502) );
  AO22X1 U461 ( .IN1(n504), .IN2(n428), .IN3(n447), .IN4(n503), .Q(n167) );
  XOR2X1 U462 ( .IN1(b[8]), .IN2(n417), .Q(n503) );
  AO22X1 U463 ( .IN1(n448), .IN2(n428), .IN3(n447), .IN4(n504), .Q(n166) );
  XOR2X1 U464 ( .IN1(b[9]), .IN2(n417), .Q(n504) );
  XOR2X1 U465 ( .IN1(b[10]), .IN2(n417), .Q(n448) );
  OAI21X1 U466 ( .IN1(n428), .IN2(n447), .IN3(n446), .QN(n165) );
  XOR2X1 U467 ( .IN1(b[11]), .IN2(n417), .Q(n446) );
  NOR2X0 U468 ( .IN1(n505), .IN2(n426), .QN(n164) );
  AO22X1 U469 ( .IN1(n506), .IN2(n427), .IN3(n450), .IN4(n507), .Q(n163) );
  XOR2X1 U470 ( .IN1(n408), .IN2(n419), .Q(n507) );
  AO22X1 U471 ( .IN1(n508), .IN2(n427), .IN3(n450), .IN4(n506), .Q(n162) );
  XOR2X1 U472 ( .IN1(b[1]), .IN2(n419), .Q(n506) );
  AO22X1 U473 ( .IN1(n509), .IN2(n427), .IN3(n450), .IN4(n508), .Q(n161) );
  XOR2X1 U474 ( .IN1(b[2]), .IN2(n419), .Q(n508) );
  AO22X1 U475 ( .IN1(n510), .IN2(n427), .IN3(n450), .IN4(n509), .Q(n160) );
  XOR2X1 U476 ( .IN1(b[3]), .IN2(n419), .Q(n509) );
  AO22X1 U477 ( .IN1(n511), .IN2(n427), .IN3(n450), .IN4(n510), .Q(n159) );
  XOR2X1 U478 ( .IN1(b[4]), .IN2(n419), .Q(n510) );
  AO22X1 U479 ( .IN1(n512), .IN2(n427), .IN3(n450), .IN4(n511), .Q(n158) );
  XOR2X1 U480 ( .IN1(b[5]), .IN2(n419), .Q(n511) );
  AO22X1 U481 ( .IN1(n513), .IN2(n427), .IN3(n450), .IN4(n512), .Q(n157) );
  XOR2X1 U482 ( .IN1(b[6]), .IN2(n419), .Q(n512) );
  AO22X1 U483 ( .IN1(n514), .IN2(n427), .IN3(n450), .IN4(n513), .Q(n156) );
  XOR2X1 U484 ( .IN1(b[7]), .IN2(n419), .Q(n513) );
  AO22X1 U485 ( .IN1(n515), .IN2(n427), .IN3(n450), .IN4(n514), .Q(n155) );
  XOR2X1 U486 ( .IN1(b[8]), .IN2(n419), .Q(n514) );
  AO22X1 U487 ( .IN1(n451), .IN2(n427), .IN3(n450), .IN4(n515), .Q(n154) );
  XOR2X1 U488 ( .IN1(b[9]), .IN2(n419), .Q(n515) );
  XOR2X1 U489 ( .IN1(b[10]), .IN2(n419), .Q(n451) );
  OAI21X1 U490 ( .IN1(n427), .IN2(n450), .IN3(n449), .QN(n153) );
  XOR2X1 U491 ( .IN1(b[11]), .IN2(n419), .Q(n449) );
  AO21X1 U492 ( .IN1(a[1]), .IN2(n426), .IN3(n437), .Q(n152) );
  AO22X1 U493 ( .IN1(n516), .IN2(n412), .IN3(n435), .IN4(n412), .Q(n151) );
  XOR2X1 U494 ( .IN1(n411), .IN2(a[2]), .Q(n517) );
  NOR2X0 U495 ( .IN1(n408), .IN2(n462), .QN(n516) );
  XNOR2X1 U496 ( .IN1(a[2]), .IN2(a[1]), .Q(n462) );
  AO22X1 U497 ( .IN1(n518), .IN2(n414), .IN3(n441), .IN4(n414), .Q(n150) );
  XOR2X1 U498 ( .IN1(n413), .IN2(a[4]), .Q(n519) );
  NOR2X0 U499 ( .IN1(n408), .IN2(n472), .QN(n518) );
  XNOR2X1 U500 ( .IN1(a[4]), .IN2(n411), .Q(n472) );
  AO22X1 U501 ( .IN1(n520), .IN2(n416), .IN3(n444), .IN4(n416), .Q(n149) );
  XOR2X1 U502 ( .IN1(n415), .IN2(a[6]), .Q(n521) );
  NOR2X0 U503 ( .IN1(n408), .IN2(n483), .QN(n520) );
  XNOR2X1 U504 ( .IN1(a[6]), .IN2(n413), .Q(n483) );
  AO22X1 U505 ( .IN1(n522), .IN2(n418), .IN3(n447), .IN4(n418), .Q(n148) );
  XOR2X1 U506 ( .IN1(n417), .IN2(a[8]), .Q(n523) );
  NOR2X0 U507 ( .IN1(n408), .IN2(n494), .QN(n522) );
  XNOR2X1 U508 ( .IN1(a[8]), .IN2(n415), .Q(n494) );
  AO22X1 U509 ( .IN1(n524), .IN2(a[11]), .IN3(n450), .IN4(n419), .Q(n147) );
  XOR2X1 U510 ( .IN1(n419), .IN2(a[10]), .Q(n525) );
  NOR2X0 U511 ( .IN1(n408), .IN2(n505), .QN(n524) );
  XNOR2X1 U512 ( .IN1(a[10]), .IN2(n417), .Q(n505) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_18 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_18_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_17_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n425), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U6 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U20 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n424), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n423), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n422), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n421), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(n25), .ZN(n425) );
  INVX0 U312 ( .INP(n3), .ZN(product[23]) );
  INVX0 U313 ( .INP(n55), .ZN(n422) );
  INVX0 U314 ( .INP(n462), .ZN(n431) );
  INVX0 U315 ( .INP(n408), .ZN(n426) );
  AND2X1 U316 ( .IN1(a[1]), .IN2(n410), .Q(n437) );
  INVX0 U317 ( .INP(n472), .ZN(n430) );
  INVX0 U318 ( .INP(n483), .ZN(n429) );
  INVX0 U319 ( .INP(n494), .ZN(n428) );
  INVX0 U320 ( .INP(n505), .ZN(n427) );
  INVX0 U321 ( .INP(n73), .ZN(n421) );
  INVX0 U322 ( .INP(n31), .ZN(n424) );
  INVX0 U323 ( .INP(n41), .ZN(n423) );
  NBUFFX2 U324 ( .INP(b[0]), .Z(n408) );
  AND2X1 U325 ( .IN1(n462), .IN2(n517), .Q(n435) );
  NBUFFX2 U326 ( .INP(a[3]), .Z(n412) );
  NBUFFX2 U327 ( .INP(a[3]), .Z(n411) );
  NBUFFX2 U328 ( .INP(a[5]), .Z(n413) );
  NBUFFX2 U329 ( .INP(a[7]), .Z(n415) );
  AND2X1 U330 ( .IN1(n483), .IN2(n521), .Q(n444) );
  AND2X1 U331 ( .IN1(n472), .IN2(n519), .Q(n441) );
  NBUFFX2 U332 ( .INP(a[5]), .Z(n414) );
  NBUFFX2 U333 ( .INP(a[9]), .Z(n417) );
  NBUFFX2 U334 ( .INP(a[11]), .Z(n419) );
  AND2X1 U335 ( .IN1(n494), .IN2(n523), .Q(n447) );
  AND2X1 U336 ( .IN1(n505), .IN2(n525), .Q(n450) );
  NBUFFX2 U337 ( .INP(a[7]), .Z(n416) );
  NBUFFX2 U338 ( .INP(a[9]), .Z(n418) );
  INVX0 U339 ( .INP(n410), .ZN(n409) );
  INVX0 U340 ( .INP(a[0]), .ZN(n410) );
  NOR2X0 U341 ( .IN1(n410), .IN2(n426), .QN(product[0]) );
  XNOR2X1 U342 ( .IN1(n432), .IN2(n433), .Q(n84) );
  NAND2X0 U343 ( .IN1(n433), .IN2(n432), .QN(n83) );
  AOI22X1 U344 ( .IN1(n434), .IN2(n431), .IN3(n435), .IN4(n436), .QN(n432) );
  OA21X1 U345 ( .IN1(n437), .IN2(n409), .IN3(n438), .Q(n433) );
  AO22X1 U346 ( .IN1(n439), .IN2(n431), .IN3(n435), .IN4(n434), .Q(n73) );
  XOR2X1 U347 ( .IN1(b[10]), .IN2(n411), .Q(n434) );
  AO22X1 U348 ( .IN1(n440), .IN2(n430), .IN3(n441), .IN4(n442), .Q(n55) );
  AO22X1 U349 ( .IN1(n443), .IN2(n429), .IN3(n444), .IN4(n445), .Q(n41) );
  AO22X1 U350 ( .IN1(n446), .IN2(n428), .IN3(n447), .IN4(n448), .Q(n31) );
  AO22X1 U351 ( .IN1(n449), .IN2(n427), .IN3(n450), .IN4(n451), .Q(n25) );
  AO22X1 U352 ( .IN1(n409), .IN2(n452), .IN3(n437), .IN4(n426), .Q(n224) );
  AO22X1 U353 ( .IN1(n409), .IN2(n453), .IN3(n437), .IN4(n452), .Q(n223) );
  XOR2X1 U354 ( .IN1(b[1]), .IN2(a[1]), .Q(n452) );
  AO22X1 U355 ( .IN1(n409), .IN2(n454), .IN3(n437), .IN4(n453), .Q(n222) );
  XOR2X1 U356 ( .IN1(b[2]), .IN2(a[1]), .Q(n453) );
  AO22X1 U357 ( .IN1(n409), .IN2(n455), .IN3(n437), .IN4(n454), .Q(n221) );
  XOR2X1 U358 ( .IN1(b[3]), .IN2(a[1]), .Q(n454) );
  AO22X1 U359 ( .IN1(n409), .IN2(n456), .IN3(n437), .IN4(n455), .Q(n220) );
  XOR2X1 U360 ( .IN1(b[4]), .IN2(a[1]), .Q(n455) );
  AO22X1 U361 ( .IN1(n409), .IN2(n457), .IN3(n437), .IN4(n456), .Q(n219) );
  XOR2X1 U362 ( .IN1(b[5]), .IN2(a[1]), .Q(n456) );
  AO22X1 U363 ( .IN1(n409), .IN2(n458), .IN3(n437), .IN4(n457), .Q(n218) );
  XOR2X1 U364 ( .IN1(b[6]), .IN2(a[1]), .Q(n457) );
  AO22X1 U365 ( .IN1(n409), .IN2(n459), .IN3(n437), .IN4(n458), .Q(n217) );
  XOR2X1 U366 ( .IN1(b[7]), .IN2(a[1]), .Q(n458) );
  AO22X1 U367 ( .IN1(n409), .IN2(n460), .IN3(n437), .IN4(n459), .Q(n216) );
  XOR2X1 U368 ( .IN1(b[8]), .IN2(a[1]), .Q(n459) );
  AO22X1 U369 ( .IN1(n409), .IN2(n461), .IN3(n437), .IN4(n460), .Q(n215) );
  XOR2X1 U370 ( .IN1(b[9]), .IN2(a[1]), .Q(n460) );
  AO22X1 U371 ( .IN1(n409), .IN2(n438), .IN3(n437), .IN4(n461), .Q(n214) );
  XOR2X1 U372 ( .IN1(b[10]), .IN2(a[1]), .Q(n461) );
  XOR2X1 U373 ( .IN1(b[11]), .IN2(a[1]), .Q(n438) );
  NOR2X0 U374 ( .IN1(n462), .IN2(n426), .QN(n212) );
  AO22X1 U375 ( .IN1(n463), .IN2(n431), .IN3(n435), .IN4(n464), .Q(n211) );
  XOR2X1 U376 ( .IN1(n408), .IN2(n411), .Q(n464) );
  AO22X1 U377 ( .IN1(n465), .IN2(n431), .IN3(n435), .IN4(n463), .Q(n210) );
  XOR2X1 U378 ( .IN1(b[1]), .IN2(n411), .Q(n463) );
  AO22X1 U379 ( .IN1(n466), .IN2(n431), .IN3(n435), .IN4(n465), .Q(n209) );
  XOR2X1 U380 ( .IN1(b[2]), .IN2(n411), .Q(n465) );
  AO22X1 U381 ( .IN1(n467), .IN2(n431), .IN3(n435), .IN4(n466), .Q(n208) );
  XOR2X1 U382 ( .IN1(b[3]), .IN2(n411), .Q(n466) );
  AO22X1 U383 ( .IN1(n468), .IN2(n431), .IN3(n435), .IN4(n467), .Q(n207) );
  XOR2X1 U384 ( .IN1(b[4]), .IN2(n411), .Q(n467) );
  AO22X1 U385 ( .IN1(n469), .IN2(n431), .IN3(n435), .IN4(n468), .Q(n206) );
  XOR2X1 U386 ( .IN1(b[5]), .IN2(n411), .Q(n468) );
  AO22X1 U387 ( .IN1(n470), .IN2(n431), .IN3(n435), .IN4(n469), .Q(n205) );
  XOR2X1 U388 ( .IN1(b[6]), .IN2(n411), .Q(n469) );
  AO22X1 U389 ( .IN1(n471), .IN2(n431), .IN3(n435), .IN4(n470), .Q(n204) );
  XOR2X1 U390 ( .IN1(b[7]), .IN2(n411), .Q(n470) );
  AO22X1 U391 ( .IN1(n436), .IN2(n431), .IN3(n435), .IN4(n471), .Q(n203) );
  XOR2X1 U392 ( .IN1(b[8]), .IN2(n411), .Q(n471) );
  XOR2X1 U393 ( .IN1(b[9]), .IN2(n411), .Q(n436) );
  OAI21X1 U394 ( .IN1(n431), .IN2(n435), .IN3(n439), .QN(n201) );
  XOR2X1 U395 ( .IN1(b[11]), .IN2(n411), .Q(n439) );
  NOR2X0 U396 ( .IN1(n472), .IN2(n426), .QN(n200) );
  AO22X1 U397 ( .IN1(n473), .IN2(n430), .IN3(n441), .IN4(n474), .Q(n199) );
  XOR2X1 U398 ( .IN1(n408), .IN2(n413), .Q(n474) );
  AO22X1 U399 ( .IN1(n475), .IN2(n430), .IN3(n441), .IN4(n473), .Q(n198) );
  XOR2X1 U400 ( .IN1(b[1]), .IN2(n413), .Q(n473) );
  AO22X1 U401 ( .IN1(n476), .IN2(n430), .IN3(n441), .IN4(n475), .Q(n197) );
  XOR2X1 U402 ( .IN1(b[2]), .IN2(n413), .Q(n475) );
  AO22X1 U403 ( .IN1(n477), .IN2(n430), .IN3(n441), .IN4(n476), .Q(n196) );
  XOR2X1 U404 ( .IN1(b[3]), .IN2(n413), .Q(n476) );
  AO22X1 U405 ( .IN1(n478), .IN2(n430), .IN3(n441), .IN4(n477), .Q(n195) );
  XOR2X1 U406 ( .IN1(b[4]), .IN2(n413), .Q(n477) );
  AO22X1 U407 ( .IN1(n479), .IN2(n430), .IN3(n441), .IN4(n478), .Q(n194) );
  XOR2X1 U408 ( .IN1(b[5]), .IN2(n413), .Q(n478) );
  AO22X1 U409 ( .IN1(n480), .IN2(n430), .IN3(n441), .IN4(n479), .Q(n193) );
  XOR2X1 U410 ( .IN1(b[6]), .IN2(n413), .Q(n479) );
  AO22X1 U411 ( .IN1(n481), .IN2(n430), .IN3(n441), .IN4(n480), .Q(n192) );
  XOR2X1 U412 ( .IN1(b[7]), .IN2(n413), .Q(n480) );
  AO22X1 U413 ( .IN1(n482), .IN2(n430), .IN3(n441), .IN4(n481), .Q(n191) );
  XOR2X1 U414 ( .IN1(b[8]), .IN2(n413), .Q(n481) );
  AO22X1 U415 ( .IN1(n442), .IN2(n430), .IN3(n441), .IN4(n482), .Q(n190) );
  XOR2X1 U416 ( .IN1(b[9]), .IN2(n413), .Q(n482) );
  XOR2X1 U417 ( .IN1(b[10]), .IN2(n413), .Q(n442) );
  OAI21X1 U418 ( .IN1(n430), .IN2(n441), .IN3(n440), .QN(n189) );
  XOR2X1 U419 ( .IN1(b[11]), .IN2(n413), .Q(n440) );
  NOR2X0 U420 ( .IN1(n483), .IN2(n426), .QN(n188) );
  AO22X1 U421 ( .IN1(n484), .IN2(n429), .IN3(n444), .IN4(n485), .Q(n187) );
  XOR2X1 U422 ( .IN1(n408), .IN2(n415), .Q(n485) );
  AO22X1 U423 ( .IN1(n486), .IN2(n429), .IN3(n444), .IN4(n484), .Q(n186) );
  XOR2X1 U424 ( .IN1(b[1]), .IN2(n415), .Q(n484) );
  AO22X1 U425 ( .IN1(n487), .IN2(n429), .IN3(n444), .IN4(n486), .Q(n185) );
  XOR2X1 U426 ( .IN1(b[2]), .IN2(n415), .Q(n486) );
  AO22X1 U427 ( .IN1(n488), .IN2(n429), .IN3(n444), .IN4(n487), .Q(n184) );
  XOR2X1 U428 ( .IN1(b[3]), .IN2(n415), .Q(n487) );
  AO22X1 U429 ( .IN1(n489), .IN2(n429), .IN3(n444), .IN4(n488), .Q(n183) );
  XOR2X1 U430 ( .IN1(b[4]), .IN2(n415), .Q(n488) );
  AO22X1 U431 ( .IN1(n490), .IN2(n429), .IN3(n444), .IN4(n489), .Q(n182) );
  XOR2X1 U432 ( .IN1(b[5]), .IN2(n415), .Q(n489) );
  AO22X1 U433 ( .IN1(n491), .IN2(n429), .IN3(n444), .IN4(n490), .Q(n181) );
  XOR2X1 U434 ( .IN1(b[6]), .IN2(n415), .Q(n490) );
  AO22X1 U435 ( .IN1(n492), .IN2(n429), .IN3(n444), .IN4(n491), .Q(n180) );
  XOR2X1 U436 ( .IN1(b[7]), .IN2(n415), .Q(n491) );
  AO22X1 U437 ( .IN1(n493), .IN2(n429), .IN3(n444), .IN4(n492), .Q(n179) );
  XOR2X1 U438 ( .IN1(b[8]), .IN2(n415), .Q(n492) );
  AO22X1 U439 ( .IN1(n445), .IN2(n429), .IN3(n444), .IN4(n493), .Q(n178) );
  XOR2X1 U440 ( .IN1(b[9]), .IN2(n415), .Q(n493) );
  XOR2X1 U441 ( .IN1(b[10]), .IN2(n415), .Q(n445) );
  OAI21X1 U442 ( .IN1(n429), .IN2(n444), .IN3(n443), .QN(n177) );
  XOR2X1 U443 ( .IN1(b[11]), .IN2(n415), .Q(n443) );
  NOR2X0 U444 ( .IN1(n494), .IN2(n426), .QN(n176) );
  AO22X1 U445 ( .IN1(n495), .IN2(n428), .IN3(n447), .IN4(n496), .Q(n175) );
  XOR2X1 U446 ( .IN1(n408), .IN2(n417), .Q(n496) );
  AO22X1 U447 ( .IN1(n497), .IN2(n428), .IN3(n447), .IN4(n495), .Q(n174) );
  XOR2X1 U448 ( .IN1(b[1]), .IN2(n417), .Q(n495) );
  AO22X1 U449 ( .IN1(n498), .IN2(n428), .IN3(n447), .IN4(n497), .Q(n173) );
  XOR2X1 U450 ( .IN1(b[2]), .IN2(n417), .Q(n497) );
  AO22X1 U451 ( .IN1(n499), .IN2(n428), .IN3(n447), .IN4(n498), .Q(n172) );
  XOR2X1 U452 ( .IN1(b[3]), .IN2(n417), .Q(n498) );
  AO22X1 U453 ( .IN1(n500), .IN2(n428), .IN3(n447), .IN4(n499), .Q(n171) );
  XOR2X1 U454 ( .IN1(b[4]), .IN2(n417), .Q(n499) );
  AO22X1 U455 ( .IN1(n501), .IN2(n428), .IN3(n447), .IN4(n500), .Q(n170) );
  XOR2X1 U456 ( .IN1(b[5]), .IN2(n417), .Q(n500) );
  AO22X1 U457 ( .IN1(n502), .IN2(n428), .IN3(n447), .IN4(n501), .Q(n169) );
  XOR2X1 U458 ( .IN1(b[6]), .IN2(n417), .Q(n501) );
  AO22X1 U459 ( .IN1(n503), .IN2(n428), .IN3(n447), .IN4(n502), .Q(n168) );
  XOR2X1 U460 ( .IN1(b[7]), .IN2(n417), .Q(n502) );
  AO22X1 U461 ( .IN1(n504), .IN2(n428), .IN3(n447), .IN4(n503), .Q(n167) );
  XOR2X1 U462 ( .IN1(b[8]), .IN2(n417), .Q(n503) );
  AO22X1 U463 ( .IN1(n448), .IN2(n428), .IN3(n447), .IN4(n504), .Q(n166) );
  XOR2X1 U464 ( .IN1(b[9]), .IN2(n417), .Q(n504) );
  XOR2X1 U465 ( .IN1(b[10]), .IN2(n417), .Q(n448) );
  OAI21X1 U466 ( .IN1(n428), .IN2(n447), .IN3(n446), .QN(n165) );
  XOR2X1 U467 ( .IN1(b[11]), .IN2(n417), .Q(n446) );
  NOR2X0 U468 ( .IN1(n505), .IN2(n426), .QN(n164) );
  AO22X1 U469 ( .IN1(n506), .IN2(n427), .IN3(n450), .IN4(n507), .Q(n163) );
  XOR2X1 U470 ( .IN1(n408), .IN2(n419), .Q(n507) );
  AO22X1 U471 ( .IN1(n508), .IN2(n427), .IN3(n450), .IN4(n506), .Q(n162) );
  XOR2X1 U472 ( .IN1(b[1]), .IN2(n419), .Q(n506) );
  AO22X1 U473 ( .IN1(n509), .IN2(n427), .IN3(n450), .IN4(n508), .Q(n161) );
  XOR2X1 U474 ( .IN1(b[2]), .IN2(n419), .Q(n508) );
  AO22X1 U475 ( .IN1(n510), .IN2(n427), .IN3(n450), .IN4(n509), .Q(n160) );
  XOR2X1 U476 ( .IN1(b[3]), .IN2(n419), .Q(n509) );
  AO22X1 U477 ( .IN1(n511), .IN2(n427), .IN3(n450), .IN4(n510), .Q(n159) );
  XOR2X1 U478 ( .IN1(b[4]), .IN2(n419), .Q(n510) );
  AO22X1 U479 ( .IN1(n512), .IN2(n427), .IN3(n450), .IN4(n511), .Q(n158) );
  XOR2X1 U480 ( .IN1(b[5]), .IN2(n419), .Q(n511) );
  AO22X1 U481 ( .IN1(n513), .IN2(n427), .IN3(n450), .IN4(n512), .Q(n157) );
  XOR2X1 U482 ( .IN1(b[6]), .IN2(n419), .Q(n512) );
  AO22X1 U483 ( .IN1(n514), .IN2(n427), .IN3(n450), .IN4(n513), .Q(n156) );
  XOR2X1 U484 ( .IN1(b[7]), .IN2(n419), .Q(n513) );
  AO22X1 U485 ( .IN1(n515), .IN2(n427), .IN3(n450), .IN4(n514), .Q(n155) );
  XOR2X1 U486 ( .IN1(b[8]), .IN2(n419), .Q(n514) );
  AO22X1 U487 ( .IN1(n451), .IN2(n427), .IN3(n450), .IN4(n515), .Q(n154) );
  XOR2X1 U488 ( .IN1(b[9]), .IN2(n419), .Q(n515) );
  XOR2X1 U489 ( .IN1(b[10]), .IN2(n419), .Q(n451) );
  OAI21X1 U490 ( .IN1(n427), .IN2(n450), .IN3(n449), .QN(n153) );
  XOR2X1 U491 ( .IN1(b[11]), .IN2(n419), .Q(n449) );
  AO21X1 U492 ( .IN1(a[1]), .IN2(n426), .IN3(n437), .Q(n152) );
  AO22X1 U493 ( .IN1(n516), .IN2(n412), .IN3(n435), .IN4(n412), .Q(n151) );
  XOR2X1 U494 ( .IN1(n411), .IN2(a[2]), .Q(n517) );
  NOR2X0 U495 ( .IN1(n408), .IN2(n462), .QN(n516) );
  XNOR2X1 U496 ( .IN1(a[2]), .IN2(a[1]), .Q(n462) );
  AO22X1 U497 ( .IN1(n518), .IN2(n414), .IN3(n441), .IN4(n414), .Q(n150) );
  XOR2X1 U498 ( .IN1(n413), .IN2(a[4]), .Q(n519) );
  NOR2X0 U499 ( .IN1(n408), .IN2(n472), .QN(n518) );
  XNOR2X1 U500 ( .IN1(a[4]), .IN2(n411), .Q(n472) );
  AO22X1 U501 ( .IN1(n520), .IN2(n416), .IN3(n444), .IN4(n416), .Q(n149) );
  XOR2X1 U502 ( .IN1(n415), .IN2(a[6]), .Q(n521) );
  NOR2X0 U503 ( .IN1(n408), .IN2(n483), .QN(n520) );
  XNOR2X1 U504 ( .IN1(a[6]), .IN2(n413), .Q(n483) );
  AO22X1 U505 ( .IN1(n522), .IN2(n418), .IN3(n447), .IN4(n418), .Q(n148) );
  XOR2X1 U506 ( .IN1(n417), .IN2(a[8]), .Q(n523) );
  NOR2X0 U507 ( .IN1(n408), .IN2(n494), .QN(n522) );
  XNOR2X1 U508 ( .IN1(a[8]), .IN2(n415), .Q(n494) );
  AO22X1 U509 ( .IN1(n524), .IN2(a[11]), .IN3(n450), .IN4(n419), .Q(n147) );
  XOR2X1 U510 ( .IN1(n419), .IN2(a[10]), .Q(n525) );
  NOR2X0 U511 ( .IN1(n408), .IN2(n505), .QN(n524) );
  XNOR2X1 U512 ( .IN1(a[10]), .IN2(n417), .Q(n505) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_17 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_17_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_16_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n422), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U6 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U20 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n424), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n426), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n428), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n430), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(n25), .ZN(n422) );
  INVX0 U312 ( .INP(n3), .ZN(product[23]) );
  INVX0 U313 ( .INP(n55), .ZN(n428) );
  NBUFFX2 U314 ( .INP(a[1]), .Z(n409) );
  INVX0 U315 ( .INP(n463), .ZN(n431) );
  AND2X1 U316 ( .IN1(n409), .IN2(n411), .Q(n438) );
  INVX0 U317 ( .INP(n408), .ZN(n432) );
  INVX0 U318 ( .INP(n473), .ZN(n429) );
  INVX0 U319 ( .INP(n484), .ZN(n427) );
  INVX0 U320 ( .INP(n73), .ZN(n430) );
  INVX0 U321 ( .INP(n495), .ZN(n425) );
  INVX0 U322 ( .INP(n506), .ZN(n423) );
  INVX0 U323 ( .INP(n31), .ZN(n424) );
  INVX0 U324 ( .INP(n41), .ZN(n426) );
  AND2X1 U325 ( .IN1(n463), .IN2(n518), .Q(n436) );
  NBUFFX2 U326 ( .INP(a[3]), .Z(n413) );
  NBUFFX2 U327 ( .INP(b[0]), .Z(n408) );
  NBUFFX2 U328 ( .INP(a[5]), .Z(n415) );
  NBUFFX2 U329 ( .INP(a[3]), .Z(n412) );
  NBUFFX2 U330 ( .INP(a[5]), .Z(n414) );
  NBUFFX2 U331 ( .INP(a[7]), .Z(n416) );
  AND2X1 U332 ( .IN1(n484), .IN2(n522), .Q(n445) );
  AND2X1 U333 ( .IN1(n473), .IN2(n520), .Q(n442) );
  NBUFFX2 U334 ( .INP(a[9]), .Z(n418) );
  NBUFFX2 U335 ( .INP(a[11]), .Z(n420) );
  AND2X1 U336 ( .IN1(n495), .IN2(n524), .Q(n448) );
  AND2X1 U337 ( .IN1(n506), .IN2(n526), .Q(n451) );
  NBUFFX2 U338 ( .INP(a[7]), .Z(n417) );
  NBUFFX2 U339 ( .INP(a[9]), .Z(n419) );
  INVX0 U340 ( .INP(n411), .ZN(n410) );
  INVX0 U341 ( .INP(a[0]), .ZN(n411) );
  NOR2X0 U342 ( .IN1(n411), .IN2(n432), .QN(product[0]) );
  XNOR2X1 U343 ( .IN1(n433), .IN2(n434), .Q(n84) );
  NAND2X0 U344 ( .IN1(n434), .IN2(n433), .QN(n83) );
  AOI22X1 U345 ( .IN1(n435), .IN2(n431), .IN3(n436), .IN4(n437), .QN(n433) );
  OA21X1 U346 ( .IN1(n438), .IN2(n410), .IN3(n439), .Q(n434) );
  AO22X1 U347 ( .IN1(n440), .IN2(n431), .IN3(n436), .IN4(n435), .Q(n73) );
  XOR2X1 U348 ( .IN1(b[10]), .IN2(n412), .Q(n435) );
  AO22X1 U349 ( .IN1(n441), .IN2(n429), .IN3(n442), .IN4(n443), .Q(n55) );
  AO22X1 U350 ( .IN1(n444), .IN2(n427), .IN3(n445), .IN4(n446), .Q(n41) );
  AO22X1 U351 ( .IN1(n447), .IN2(n425), .IN3(n448), .IN4(n449), .Q(n31) );
  AO22X1 U352 ( .IN1(n450), .IN2(n423), .IN3(n451), .IN4(n452), .Q(n25) );
  AO22X1 U353 ( .IN1(n410), .IN2(n453), .IN3(n438), .IN4(n432), .Q(n224) );
  AO22X1 U354 ( .IN1(n410), .IN2(n454), .IN3(n438), .IN4(n453), .Q(n223) );
  XOR2X1 U355 ( .IN1(b[1]), .IN2(n409), .Q(n453) );
  AO22X1 U356 ( .IN1(n410), .IN2(n455), .IN3(n438), .IN4(n454), .Q(n222) );
  XOR2X1 U357 ( .IN1(b[2]), .IN2(n409), .Q(n454) );
  AO22X1 U358 ( .IN1(n410), .IN2(n456), .IN3(n438), .IN4(n455), .Q(n221) );
  XOR2X1 U359 ( .IN1(b[3]), .IN2(n409), .Q(n455) );
  AO22X1 U360 ( .IN1(n410), .IN2(n457), .IN3(n438), .IN4(n456), .Q(n220) );
  XOR2X1 U361 ( .IN1(b[4]), .IN2(n409), .Q(n456) );
  AO22X1 U362 ( .IN1(n410), .IN2(n458), .IN3(n438), .IN4(n457), .Q(n219) );
  XOR2X1 U363 ( .IN1(b[5]), .IN2(n409), .Q(n457) );
  AO22X1 U364 ( .IN1(n410), .IN2(n459), .IN3(n438), .IN4(n458), .Q(n218) );
  XOR2X1 U365 ( .IN1(b[6]), .IN2(n409), .Q(n458) );
  AO22X1 U366 ( .IN1(n410), .IN2(n460), .IN3(n438), .IN4(n459), .Q(n217) );
  XOR2X1 U367 ( .IN1(b[7]), .IN2(n409), .Q(n459) );
  AO22X1 U368 ( .IN1(n410), .IN2(n461), .IN3(n438), .IN4(n460), .Q(n216) );
  XOR2X1 U369 ( .IN1(b[8]), .IN2(n409), .Q(n460) );
  AO22X1 U370 ( .IN1(n410), .IN2(n462), .IN3(n438), .IN4(n461), .Q(n215) );
  XOR2X1 U371 ( .IN1(b[9]), .IN2(n409), .Q(n461) );
  AO22X1 U372 ( .IN1(n410), .IN2(n439), .IN3(n438), .IN4(n462), .Q(n214) );
  XOR2X1 U373 ( .IN1(b[10]), .IN2(n409), .Q(n462) );
  XOR2X1 U374 ( .IN1(b[11]), .IN2(n409), .Q(n439) );
  NOR2X0 U375 ( .IN1(n463), .IN2(n432), .QN(n212) );
  AO22X1 U376 ( .IN1(n464), .IN2(n431), .IN3(n436), .IN4(n465), .Q(n211) );
  XOR2X1 U377 ( .IN1(n408), .IN2(n412), .Q(n465) );
  AO22X1 U378 ( .IN1(n466), .IN2(n431), .IN3(n436), .IN4(n464), .Q(n210) );
  XOR2X1 U379 ( .IN1(b[1]), .IN2(n412), .Q(n464) );
  AO22X1 U380 ( .IN1(n467), .IN2(n431), .IN3(n436), .IN4(n466), .Q(n209) );
  XOR2X1 U381 ( .IN1(b[2]), .IN2(n412), .Q(n466) );
  AO22X1 U382 ( .IN1(n468), .IN2(n431), .IN3(n436), .IN4(n467), .Q(n208) );
  XOR2X1 U383 ( .IN1(b[3]), .IN2(n412), .Q(n467) );
  AO22X1 U384 ( .IN1(n469), .IN2(n431), .IN3(n436), .IN4(n468), .Q(n207) );
  XOR2X1 U385 ( .IN1(b[4]), .IN2(n412), .Q(n468) );
  AO22X1 U386 ( .IN1(n470), .IN2(n431), .IN3(n436), .IN4(n469), .Q(n206) );
  XOR2X1 U387 ( .IN1(b[5]), .IN2(n412), .Q(n469) );
  AO22X1 U388 ( .IN1(n471), .IN2(n431), .IN3(n436), .IN4(n470), .Q(n205) );
  XOR2X1 U389 ( .IN1(b[6]), .IN2(n412), .Q(n470) );
  AO22X1 U390 ( .IN1(n472), .IN2(n431), .IN3(n436), .IN4(n471), .Q(n204) );
  XOR2X1 U391 ( .IN1(b[7]), .IN2(n412), .Q(n471) );
  AO22X1 U392 ( .IN1(n437), .IN2(n431), .IN3(n436), .IN4(n472), .Q(n203) );
  XOR2X1 U393 ( .IN1(b[8]), .IN2(n412), .Q(n472) );
  XOR2X1 U394 ( .IN1(b[9]), .IN2(n412), .Q(n437) );
  OAI21X1 U395 ( .IN1(n431), .IN2(n436), .IN3(n440), .QN(n201) );
  XOR2X1 U396 ( .IN1(b[11]), .IN2(n412), .Q(n440) );
  NOR2X0 U397 ( .IN1(n473), .IN2(n432), .QN(n200) );
  AO22X1 U398 ( .IN1(n474), .IN2(n429), .IN3(n442), .IN4(n475), .Q(n199) );
  XOR2X1 U399 ( .IN1(n408), .IN2(n414), .Q(n475) );
  AO22X1 U400 ( .IN1(n476), .IN2(n429), .IN3(n442), .IN4(n474), .Q(n198) );
  XOR2X1 U401 ( .IN1(b[1]), .IN2(n414), .Q(n474) );
  AO22X1 U402 ( .IN1(n477), .IN2(n429), .IN3(n442), .IN4(n476), .Q(n197) );
  XOR2X1 U403 ( .IN1(b[2]), .IN2(n414), .Q(n476) );
  AO22X1 U404 ( .IN1(n478), .IN2(n429), .IN3(n442), .IN4(n477), .Q(n196) );
  XOR2X1 U405 ( .IN1(b[3]), .IN2(n414), .Q(n477) );
  AO22X1 U406 ( .IN1(n479), .IN2(n429), .IN3(n442), .IN4(n478), .Q(n195) );
  XOR2X1 U407 ( .IN1(b[4]), .IN2(n414), .Q(n478) );
  AO22X1 U408 ( .IN1(n480), .IN2(n429), .IN3(n442), .IN4(n479), .Q(n194) );
  XOR2X1 U409 ( .IN1(b[5]), .IN2(n414), .Q(n479) );
  AO22X1 U410 ( .IN1(n481), .IN2(n429), .IN3(n442), .IN4(n480), .Q(n193) );
  XOR2X1 U411 ( .IN1(b[6]), .IN2(n414), .Q(n480) );
  AO22X1 U412 ( .IN1(n482), .IN2(n429), .IN3(n442), .IN4(n481), .Q(n192) );
  XOR2X1 U413 ( .IN1(b[7]), .IN2(n414), .Q(n481) );
  AO22X1 U414 ( .IN1(n483), .IN2(n429), .IN3(n442), .IN4(n482), .Q(n191) );
  XOR2X1 U415 ( .IN1(b[8]), .IN2(n414), .Q(n482) );
  AO22X1 U416 ( .IN1(n443), .IN2(n429), .IN3(n442), .IN4(n483), .Q(n190) );
  XOR2X1 U417 ( .IN1(b[9]), .IN2(n414), .Q(n483) );
  XOR2X1 U418 ( .IN1(b[10]), .IN2(n414), .Q(n443) );
  OAI21X1 U419 ( .IN1(n429), .IN2(n442), .IN3(n441), .QN(n189) );
  XOR2X1 U420 ( .IN1(b[11]), .IN2(n414), .Q(n441) );
  NOR2X0 U421 ( .IN1(n484), .IN2(n432), .QN(n188) );
  AO22X1 U422 ( .IN1(n485), .IN2(n427), .IN3(n445), .IN4(n486), .Q(n187) );
  XOR2X1 U423 ( .IN1(n408), .IN2(n416), .Q(n486) );
  AO22X1 U424 ( .IN1(n487), .IN2(n427), .IN3(n445), .IN4(n485), .Q(n186) );
  XOR2X1 U425 ( .IN1(b[1]), .IN2(n416), .Q(n485) );
  AO22X1 U426 ( .IN1(n488), .IN2(n427), .IN3(n445), .IN4(n487), .Q(n185) );
  XOR2X1 U427 ( .IN1(b[2]), .IN2(n416), .Q(n487) );
  AO22X1 U428 ( .IN1(n489), .IN2(n427), .IN3(n445), .IN4(n488), .Q(n184) );
  XOR2X1 U429 ( .IN1(b[3]), .IN2(n416), .Q(n488) );
  AO22X1 U430 ( .IN1(n490), .IN2(n427), .IN3(n445), .IN4(n489), .Q(n183) );
  XOR2X1 U431 ( .IN1(b[4]), .IN2(n416), .Q(n489) );
  AO22X1 U432 ( .IN1(n491), .IN2(n427), .IN3(n445), .IN4(n490), .Q(n182) );
  XOR2X1 U433 ( .IN1(b[5]), .IN2(n416), .Q(n490) );
  AO22X1 U434 ( .IN1(n492), .IN2(n427), .IN3(n445), .IN4(n491), .Q(n181) );
  XOR2X1 U435 ( .IN1(b[6]), .IN2(n416), .Q(n491) );
  AO22X1 U436 ( .IN1(n493), .IN2(n427), .IN3(n445), .IN4(n492), .Q(n180) );
  XOR2X1 U437 ( .IN1(b[7]), .IN2(n416), .Q(n492) );
  AO22X1 U438 ( .IN1(n494), .IN2(n427), .IN3(n445), .IN4(n493), .Q(n179) );
  XOR2X1 U439 ( .IN1(b[8]), .IN2(n416), .Q(n493) );
  AO22X1 U440 ( .IN1(n446), .IN2(n427), .IN3(n445), .IN4(n494), .Q(n178) );
  XOR2X1 U441 ( .IN1(b[9]), .IN2(n416), .Q(n494) );
  XOR2X1 U442 ( .IN1(b[10]), .IN2(n416), .Q(n446) );
  OAI21X1 U443 ( .IN1(n427), .IN2(n445), .IN3(n444), .QN(n177) );
  XOR2X1 U444 ( .IN1(b[11]), .IN2(n416), .Q(n444) );
  NOR2X0 U445 ( .IN1(n495), .IN2(n432), .QN(n176) );
  AO22X1 U446 ( .IN1(n496), .IN2(n425), .IN3(n448), .IN4(n497), .Q(n175) );
  XOR2X1 U447 ( .IN1(n408), .IN2(n418), .Q(n497) );
  AO22X1 U448 ( .IN1(n498), .IN2(n425), .IN3(n448), .IN4(n496), .Q(n174) );
  XOR2X1 U449 ( .IN1(b[1]), .IN2(n418), .Q(n496) );
  AO22X1 U450 ( .IN1(n499), .IN2(n425), .IN3(n448), .IN4(n498), .Q(n173) );
  XOR2X1 U451 ( .IN1(b[2]), .IN2(n418), .Q(n498) );
  AO22X1 U452 ( .IN1(n500), .IN2(n425), .IN3(n448), .IN4(n499), .Q(n172) );
  XOR2X1 U453 ( .IN1(b[3]), .IN2(n418), .Q(n499) );
  AO22X1 U454 ( .IN1(n501), .IN2(n425), .IN3(n448), .IN4(n500), .Q(n171) );
  XOR2X1 U455 ( .IN1(b[4]), .IN2(n418), .Q(n500) );
  AO22X1 U456 ( .IN1(n502), .IN2(n425), .IN3(n448), .IN4(n501), .Q(n170) );
  XOR2X1 U457 ( .IN1(b[5]), .IN2(n418), .Q(n501) );
  AO22X1 U458 ( .IN1(n503), .IN2(n425), .IN3(n448), .IN4(n502), .Q(n169) );
  XOR2X1 U459 ( .IN1(b[6]), .IN2(n418), .Q(n502) );
  AO22X1 U460 ( .IN1(n504), .IN2(n425), .IN3(n448), .IN4(n503), .Q(n168) );
  XOR2X1 U461 ( .IN1(b[7]), .IN2(n418), .Q(n503) );
  AO22X1 U462 ( .IN1(n505), .IN2(n425), .IN3(n448), .IN4(n504), .Q(n167) );
  XOR2X1 U463 ( .IN1(b[8]), .IN2(n418), .Q(n504) );
  AO22X1 U464 ( .IN1(n449), .IN2(n425), .IN3(n448), .IN4(n505), .Q(n166) );
  XOR2X1 U465 ( .IN1(b[9]), .IN2(n418), .Q(n505) );
  XOR2X1 U466 ( .IN1(b[10]), .IN2(n418), .Q(n449) );
  OAI21X1 U467 ( .IN1(n425), .IN2(n448), .IN3(n447), .QN(n165) );
  XOR2X1 U468 ( .IN1(b[11]), .IN2(n418), .Q(n447) );
  NOR2X0 U469 ( .IN1(n506), .IN2(n432), .QN(n164) );
  AO22X1 U470 ( .IN1(n507), .IN2(n423), .IN3(n451), .IN4(n508), .Q(n163) );
  XOR2X1 U471 ( .IN1(n408), .IN2(n420), .Q(n508) );
  AO22X1 U472 ( .IN1(n509), .IN2(n423), .IN3(n451), .IN4(n507), .Q(n162) );
  XOR2X1 U473 ( .IN1(b[1]), .IN2(n420), .Q(n507) );
  AO22X1 U474 ( .IN1(n510), .IN2(n423), .IN3(n451), .IN4(n509), .Q(n161) );
  XOR2X1 U475 ( .IN1(b[2]), .IN2(n420), .Q(n509) );
  AO22X1 U476 ( .IN1(n511), .IN2(n423), .IN3(n451), .IN4(n510), .Q(n160) );
  XOR2X1 U477 ( .IN1(b[3]), .IN2(n420), .Q(n510) );
  AO22X1 U478 ( .IN1(n512), .IN2(n423), .IN3(n451), .IN4(n511), .Q(n159) );
  XOR2X1 U479 ( .IN1(b[4]), .IN2(n420), .Q(n511) );
  AO22X1 U480 ( .IN1(n513), .IN2(n423), .IN3(n451), .IN4(n512), .Q(n158) );
  XOR2X1 U481 ( .IN1(b[5]), .IN2(n420), .Q(n512) );
  AO22X1 U482 ( .IN1(n514), .IN2(n423), .IN3(n451), .IN4(n513), .Q(n157) );
  XOR2X1 U483 ( .IN1(b[6]), .IN2(n420), .Q(n513) );
  AO22X1 U484 ( .IN1(n515), .IN2(n423), .IN3(n451), .IN4(n514), .Q(n156) );
  XOR2X1 U485 ( .IN1(b[7]), .IN2(n420), .Q(n514) );
  AO22X1 U486 ( .IN1(n516), .IN2(n423), .IN3(n451), .IN4(n515), .Q(n155) );
  XOR2X1 U487 ( .IN1(b[8]), .IN2(n420), .Q(n515) );
  AO22X1 U488 ( .IN1(n452), .IN2(n423), .IN3(n451), .IN4(n516), .Q(n154) );
  XOR2X1 U489 ( .IN1(b[9]), .IN2(n420), .Q(n516) );
  XOR2X1 U490 ( .IN1(b[10]), .IN2(n420), .Q(n452) );
  OAI21X1 U491 ( .IN1(n423), .IN2(n451), .IN3(n450), .QN(n153) );
  XOR2X1 U492 ( .IN1(b[11]), .IN2(n420), .Q(n450) );
  AO21X1 U493 ( .IN1(n409), .IN2(n432), .IN3(n438), .Q(n152) );
  AO22X1 U494 ( .IN1(n517), .IN2(n413), .IN3(n436), .IN4(n413), .Q(n151) );
  XOR2X1 U495 ( .IN1(n412), .IN2(a[2]), .Q(n518) );
  NOR2X0 U496 ( .IN1(n408), .IN2(n463), .QN(n517) );
  XNOR2X1 U497 ( .IN1(a[2]), .IN2(n409), .Q(n463) );
  AO22X1 U498 ( .IN1(n519), .IN2(n415), .IN3(n442), .IN4(n415), .Q(n150) );
  XOR2X1 U499 ( .IN1(n414), .IN2(a[4]), .Q(n520) );
  NOR2X0 U500 ( .IN1(n408), .IN2(n473), .QN(n519) );
  XNOR2X1 U501 ( .IN1(a[4]), .IN2(n412), .Q(n473) );
  AO22X1 U502 ( .IN1(n521), .IN2(n417), .IN3(n445), .IN4(n417), .Q(n149) );
  XOR2X1 U503 ( .IN1(n416), .IN2(a[6]), .Q(n522) );
  NOR2X0 U504 ( .IN1(n408), .IN2(n484), .QN(n521) );
  XNOR2X1 U505 ( .IN1(a[6]), .IN2(n414), .Q(n484) );
  AO22X1 U506 ( .IN1(n523), .IN2(n419), .IN3(n448), .IN4(n419), .Q(n148) );
  XOR2X1 U507 ( .IN1(n418), .IN2(a[8]), .Q(n524) );
  NOR2X0 U508 ( .IN1(n408), .IN2(n495), .QN(n523) );
  XNOR2X1 U509 ( .IN1(a[8]), .IN2(n416), .Q(n495) );
  AO22X1 U510 ( .IN1(n525), .IN2(a[11]), .IN3(n451), .IN4(n420), .Q(n147) );
  XOR2X1 U511 ( .IN1(n420), .IN2(a[10]), .Q(n526) );
  NOR2X0 U512 ( .IN1(n408), .IN2(n506), .QN(n525) );
  XNOR2X1 U513 ( .IN1(a[10]), .IN2(n418), .Q(n506) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_16 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_16_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_4_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AO22X1 U1 ( .IN1(A[6]), .IN2(n1), .IN3(B[6]), .IN4(n2), .Q(carry[7]) );
  OR2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AO22X1 U3 ( .IN1(A[5]), .IN2(n3), .IN3(B[5]), .IN4(n4), .Q(n1) );
  OR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AO22X1 U5 ( .IN1(A[4]), .IN2(n5), .IN3(B[4]), .IN4(n6), .Q(n3) );
  OR2X1 U6 ( .IN1(n5), .IN2(A[4]), .Q(n6) );
  AO22X1 U7 ( .IN1(A[3]), .IN2(n7), .IN3(B[3]), .IN4(n8), .Q(n5) );
  OR2X1 U8 ( .IN1(n7), .IN2(A[3]), .Q(n8) );
  AO22X1 U9 ( .IN1(A[2]), .IN2(n9), .IN3(B[2]), .IN4(n10), .Q(n7) );
  OR2X1 U10 ( .IN1(n9), .IN2(A[2]), .Q(n10) );
  AO22X1 U11 ( .IN1(B[1]), .IN2(A[1]), .IN3(n11), .IN4(B[0]), .Q(n9) );
  OA21X1 U12 ( .IN1(A[1]), .IN2(B[1]), .IN3(A[0]), .Q(n11) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_4 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_4_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(\output ) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_4_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [24:0] carry;

  FADDX1 U2_22 ( .A(A[22]), .B(n7), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n8), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n9), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n10), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n11), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n12), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n13), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n18), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n21), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n22), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XNOR3X1 U1 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(DIFF[23]) );
  INVX0 U2 ( .INP(B[21]), .ZN(n8) );
  INVX0 U3 ( .INP(B[20]), .ZN(n9) );
  INVX0 U4 ( .INP(B[22]), .ZN(n7) );
  INVX0 U5 ( .INP(B[19]), .ZN(n10) );
  INVX0 U6 ( .INP(B[18]), .ZN(n11) );
  INVX0 U7 ( .INP(B[17]), .ZN(n12) );
  INVX0 U8 ( .INP(B[16]), .ZN(n13) );
  INVX0 U9 ( .INP(B[15]), .ZN(n14) );
  INVX0 U10 ( .INP(B[14]), .ZN(n15) );
  INVX0 U11 ( .INP(B[13]), .ZN(n16) );
  INVX0 U12 ( .INP(B[12]), .ZN(n17) );
  INVX0 U13 ( .INP(B[11]), .ZN(n18) );
  INVX0 U14 ( .INP(B[10]), .ZN(n19) );
  INVX0 U15 ( .INP(B[9]), .ZN(n20) );
  INVX0 U16 ( .INP(B[8]), .ZN(n21) );
  INVX0 U17 ( .INP(B[7]), .ZN(n22) );
  INVX0 U18 ( .INP(A[3]), .ZN(n4) );
  INVX0 U19 ( .INP(A[1]), .ZN(n6) );
  INVX0 U20 ( .INP(A[5]), .ZN(n2) );
  INVX0 U21 ( .INP(A[2]), .ZN(n5) );
  INVX0 U22 ( .INP(B[0]), .ZN(n23) );
  INVX0 U23 ( .INP(A[4]), .ZN(n3) );
  INVX0 U24 ( .INP(A[6]), .ZN(n1) );
  OAI22X1 U25 ( .IN1(n24), .IN2(n1), .IN3(B[6]), .IN4(n25), .QN(carry[7]) );
  AND2X1 U26 ( .IN1(n1), .IN2(n24), .Q(n25) );
  OA22X1 U27 ( .IN1(n26), .IN2(n2), .IN3(B[5]), .IN4(n27), .Q(n24) );
  AND2X1 U28 ( .IN1(n2), .IN2(n26), .Q(n27) );
  OA22X1 U29 ( .IN1(n28), .IN2(n3), .IN3(B[4]), .IN4(n29), .Q(n26) );
  AND2X1 U30 ( .IN1(n3), .IN2(n28), .Q(n29) );
  OA22X1 U31 ( .IN1(n30), .IN2(n4), .IN3(B[3]), .IN4(n31), .Q(n28) );
  AND2X1 U32 ( .IN1(n4), .IN2(n30), .Q(n31) );
  OA22X1 U33 ( .IN1(n32), .IN2(n5), .IN3(B[2]), .IN4(n33), .Q(n30) );
  AND2X1 U34 ( .IN1(n5), .IN2(n32), .Q(n33) );
  OA22X1 U35 ( .IN1(n34), .IN2(n6), .IN3(B[1]), .IN4(n35), .Q(n32) );
  AND2X1 U36 ( .IN1(n6), .IN2(n34), .Q(n35) );
  NOR2X0 U37 ( .IN1(n23), .IN2(A[0]), .QN(n34) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_4 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_4_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(\output ) );
endmodule


module complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12 ( a_r, a_i, b_r, b_i, 
        out_r, out_i, clk );
  input [11:0] a_r;
  input [11:0] a_i;
  input [11:0] b_r;
  input [11:0] b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk;
  wire   N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36;
  wire   [23:0] mult1_out;
  wire   [23:0] mult2_out;
  wire   [23:0] mult3_out;
  wire   [23:0] mult4_out;
  wire   [23:7] pre_out_r;
  wire   [23:7] pre_out_i;
  wire   [11:0] pos_out_r;
  wire   [11:0] pos_out_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFFX1 \out_r_reg_reg[11]  ( .D(pos_out_r[11]), .CLK(clk), .Q(out_r[11]) );
  DFFX1 \out_r_reg_reg[10]  ( .D(pos_out_r[10]), .CLK(clk), .Q(out_r[10]) );
  DFFX1 \out_r_reg_reg[9]  ( .D(pos_out_r[9]), .CLK(clk), .Q(out_r[9]) );
  DFFX1 \out_r_reg_reg[8]  ( .D(pos_out_r[8]), .CLK(clk), .Q(out_r[8]) );
  DFFX1 \out_r_reg_reg[7]  ( .D(pos_out_r[7]), .CLK(clk), .Q(out_r[7]) );
  DFFX1 \out_r_reg_reg[6]  ( .D(pos_out_r[6]), .CLK(clk), .Q(out_r[6]) );
  DFFX1 \out_r_reg_reg[5]  ( .D(pos_out_r[5]), .CLK(clk), .Q(out_r[5]) );
  DFFX1 \out_r_reg_reg[4]  ( .D(pos_out_r[4]), .CLK(clk), .Q(out_r[4]) );
  DFFX1 \out_r_reg_reg[3]  ( .D(pos_out_r[3]), .CLK(clk), .Q(out_r[3]) );
  DFFX1 \out_r_reg_reg[2]  ( .D(pos_out_r[2]), .CLK(clk), .Q(out_r[2]) );
  DFFX1 \out_r_reg_reg[1]  ( .D(pos_out_r[1]), .CLK(clk), .Q(out_r[1]) );
  DFFX1 \out_r_reg_reg[0]  ( .D(pos_out_r[0]), .CLK(clk), .Q(out_r[0]) );
  DFFX1 \out_i_reg_reg[11]  ( .D(pos_out_i[11]), .CLK(clk), .Q(out_i[11]) );
  DFFX1 \out_i_reg_reg[10]  ( .D(pos_out_i[10]), .CLK(clk), .Q(out_i[10]) );
  DFFX1 \out_i_reg_reg[9]  ( .D(pos_out_i[9]), .CLK(clk), .Q(out_i[9]) );
  DFFX1 \out_i_reg_reg[8]  ( .D(pos_out_i[8]), .CLK(clk), .Q(out_i[8]) );
  DFFX1 \out_i_reg_reg[7]  ( .D(pos_out_i[7]), .CLK(clk), .Q(out_i[7]) );
  DFFX1 \out_i_reg_reg[6]  ( .D(pos_out_i[6]), .CLK(clk), .Q(out_i[6]) );
  DFFX1 \out_i_reg_reg[5]  ( .D(pos_out_i[5]), .CLK(clk), .Q(out_i[5]) );
  DFFX1 \out_i_reg_reg[4]  ( .D(pos_out_i[4]), .CLK(clk), .Q(out_i[4]) );
  DFFX1 \out_i_reg_reg[3]  ( .D(pos_out_i[3]), .CLK(clk), .Q(out_i[3]) );
  DFFX1 \out_i_reg_reg[2]  ( .D(pos_out_i[2]), .CLK(clk), .Q(out_i[2]) );
  DFFX1 \out_i_reg_reg[1]  ( .D(pos_out_i[1]), .CLK(clk), .Q(out_i[1]) );
  DFFX1 \out_i_reg_reg[0]  ( .D(pos_out_i[0]), .CLK(clk), .Q(out_i[0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_19 mult1 ( .in_a({a_r[11:2], n6, a_r[0]}), 
        .in_b(b_r), .clk(clk), .\output (mult1_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_18 mult2 ( .in_a({a_i[11:2], n5, a_i[0]}), 
        .in_b(b_i), .clk(clk), .\output (mult2_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_17 mult3 ( .in_a({a_r[11:2], n6, a_r[0]}), 
        .in_b(b_i), .clk(clk), .\output (mult3_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_16 mult4 ( .in_a({a_i[11:2], n5, a_i[0]}), 
        .in_b(b_r), .clk(clk), .\output (mult4_out) );
  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_4 add ( .a(mult1_out), .b(mult2_out), .\output ({pre_out_r, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_4 sub ( .a(mult3_out), .b(mult4_out), .\output ({pre_out_i, SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_DW01_inc_0 add_155_round ( .A(
        pre_out_i[19:7]), .SUM({N108, N107, N106, N105, N104, N103, N102, N101, 
        N100, N99, N98, N97, SYNOPSYS_UNCONNECTED__14}) );
  complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12_DW01_inc_1 add_141_round ( .A(
        pre_out_r[19:7]), .SUM({N53, N52, N51, N50, N49, N48, N47, N46, N45, 
        N44, N43, N42, SYNOPSYS_UNCONNECTED__15}) );
  INVX0 U3 ( .INP(pre_out_i[23]), .ZN(n14) );
  INVX0 U4 ( .INP(pre_out_r[23]), .ZN(n29) );
  NBUFFX2 U5 ( .INP(a_i[1]), .Z(n5) );
  NBUFFX2 U6 ( .INP(a_r[1]), .Z(n6) );
  INVX0 U7 ( .INP(n15), .ZN(n17) );
  INVX0 U8 ( .INP(n30), .ZN(n32) );
  AND2X1 U9 ( .IN1(n31), .IN2(n33), .Q(n1) );
  AND2X1 U10 ( .IN1(n16), .IN2(n18), .Q(n2) );
  AND2X1 U11 ( .IN1(n32), .IN2(n33), .Q(n3) );
  AND2X1 U12 ( .IN1(n17), .IN2(n18), .Q(n4) );
  NOR2X0 U13 ( .IN1(pre_out_i[21]), .IN2(pre_out_i[22]), .QN(n7) );
  NOR2X0 U14 ( .IN1(pre_out_r[21]), .IN2(pre_out_r[22]), .QN(n22) );
  NAND2X0 U15 ( .IN1(n8), .IN2(n7), .QN(n10) );
  NOR2X0 U16 ( .IN1(pre_out_i[19]), .IN2(pre_out_i[20]), .QN(n8) );
  NAND2X0 U17 ( .IN1(n23), .IN2(n22), .QN(n25) );
  NOR2X0 U18 ( .IN1(pre_out_r[19]), .IN2(pre_out_r[20]), .QN(n23) );
  INVX0 U19 ( .INP(n35), .ZN(n28) );
  INVX0 U20 ( .INP(n33), .ZN(n34) );
  INVX0 U21 ( .INP(n18), .ZN(n19) );
  INVX0 U22 ( .INP(n20), .ZN(n13) );
  XNOR2X1 U23 ( .IN1(mult1_out[23]), .IN2(mult2_out[23]), .Q(n27) );
  NAND2X0 U24 ( .IN1(n12), .IN2(n11), .QN(n20) );
  NAND4X0 U25 ( .IN1(pre_out_i[22]), .IN2(pre_out_i[21]), .IN3(pre_out_i[20]), 
        .IN4(pre_out_i[19]), .QN(n9) );
  MUX21X1 U26 ( .IN1(n10), .IN2(n9), .S(pre_out_i[23]), .Q(n15) );
  XOR2X1 U27 ( .IN1(mult4_out[23]), .IN2(mult3_out[23]), .Q(n12) );
  XOR2X1 U28 ( .IN1(pre_out_i[23]), .IN2(mult3_out[23]), .Q(n11) );
  NAND2X1 U29 ( .IN1(mult3_out[23]), .IN2(n13), .QN(n18) );
  AO21X1 U30 ( .IN1(n15), .IN2(n14), .IN3(n13), .Q(n16) );
  AO21X1 U31 ( .IN1(N97), .IN2(n4), .IN3(n2), .Q(pos_out_i[0]) );
  AO21X1 U32 ( .IN1(N98), .IN2(n4), .IN3(n2), .Q(pos_out_i[1]) );
  AO21X1 U33 ( .IN1(N99), .IN2(n4), .IN3(n2), .Q(pos_out_i[2]) );
  AO21X1 U34 ( .IN1(N100), .IN2(n4), .IN3(n2), .Q(pos_out_i[3]) );
  AO21X1 U35 ( .IN1(N101), .IN2(n4), .IN3(n2), .Q(pos_out_i[4]) );
  AO21X1 U36 ( .IN1(N102), .IN2(n4), .IN3(n2), .Q(pos_out_i[5]) );
  AO21X1 U37 ( .IN1(N103), .IN2(n4), .IN3(n2), .Q(pos_out_i[6]) );
  AO21X1 U38 ( .IN1(N104), .IN2(n4), .IN3(n2), .Q(pos_out_i[7]) );
  AO21X1 U39 ( .IN1(N105), .IN2(n4), .IN3(n2), .Q(pos_out_i[8]) );
  AO21X1 U40 ( .IN1(N106), .IN2(n4), .IN3(n2), .Q(pos_out_i[9]) );
  AO21X1 U41 ( .IN1(N107), .IN2(n4), .IN3(n2), .Q(pos_out_i[10]) );
  MUX21X1 U42 ( .IN1(pre_out_i[23]), .IN2(N108), .S(n17), .Q(n21) );
  AO21X1 U43 ( .IN1(n21), .IN2(n20), .IN3(n19), .Q(pos_out_i[11]) );
  NAND4X0 U44 ( .IN1(pre_out_r[22]), .IN2(pre_out_r[21]), .IN3(pre_out_r[20]), 
        .IN4(pre_out_r[19]), .QN(n24) );
  MUX21X1 U45 ( .IN1(n25), .IN2(n24), .S(pre_out_r[23]), .Q(n30) );
  XOR2X1 U46 ( .IN1(pre_out_r[23]), .IN2(mult1_out[23]), .Q(n26) );
  NAND2X1 U47 ( .IN1(n27), .IN2(n26), .QN(n35) );
  NAND2X1 U48 ( .IN1(mult1_out[23]), .IN2(n28), .QN(n33) );
  AO21X1 U49 ( .IN1(n30), .IN2(n29), .IN3(n28), .Q(n31) );
  AO21X1 U50 ( .IN1(N42), .IN2(n3), .IN3(n1), .Q(pos_out_r[0]) );
  AO21X1 U51 ( .IN1(N43), .IN2(n3), .IN3(n1), .Q(pos_out_r[1]) );
  AO21X1 U52 ( .IN1(N44), .IN2(n3), .IN3(n1), .Q(pos_out_r[2]) );
  AO21X1 U53 ( .IN1(N45), .IN2(n3), .IN3(n1), .Q(pos_out_r[3]) );
  AO21X1 U54 ( .IN1(N46), .IN2(n3), .IN3(n1), .Q(pos_out_r[4]) );
  AO21X1 U55 ( .IN1(N47), .IN2(n3), .IN3(n1), .Q(pos_out_r[5]) );
  AO21X1 U56 ( .IN1(N48), .IN2(n3), .IN3(n1), .Q(pos_out_r[6]) );
  AO21X1 U57 ( .IN1(N49), .IN2(n3), .IN3(n1), .Q(pos_out_r[7]) );
  AO21X1 U58 ( .IN1(N50), .IN2(n3), .IN3(n1), .Q(pos_out_r[8]) );
  AO21X1 U59 ( .IN1(N51), .IN2(n3), .IN3(n1), .Q(pos_out_r[9]) );
  AO21X1 U60 ( .IN1(N52), .IN2(n3), .IN3(n1), .Q(pos_out_r[10]) );
  MUX21X1 U61 ( .IN1(pre_out_r[23]), .IN2(N53), .S(n32), .Q(n36) );
  AO21X1 U62 ( .IN1(n36), .IN2(n35), .IN3(n34), .Q(pos_out_r[11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_1_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [11:1] carry;

  FADDX1 U1_10 ( .A(A[10]), .B(n1), .CI(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(n2), .CI(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n12), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_11 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(SUM[11]) );
  FADDX1 U1_4 ( .A(A[4]), .B(n8), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FADDX1 U1_6 ( .A(A[6]), .B(n4), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FADDX1 U1_8 ( .A(A[8]), .B(n6), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FADDX2 U1_5 ( .A(A[5]), .B(carry[5]), .CI(B[5]), .CO(carry[6]), .S(SUM[5])
         );
  DELLN2X2 U1 ( .INP(B[10]), .Z(n1) );
  DELLN2X2 U2 ( .INP(B[9]), .Z(n2) );
  INVX0 U3 ( .INP(B[6]), .ZN(n3) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U5 ( .INP(B[8]), .ZN(n5) );
  INVX0 U6 ( .INP(n5), .ZN(n6) );
  INVX0 U7 ( .INP(B[4]), .ZN(n7) );
  INVX0 U8 ( .INP(n7), .ZN(n8) );
  XOR3X1 U9 ( .IN1(B[2]), .IN2(A[2]), .IN3(carry[2]), .Q(SUM[2]) );
  NAND2X0 U10 ( .IN1(carry[2]), .IN2(B[2]), .QN(n9) );
  NAND2X0 U11 ( .IN1(A[2]), .IN2(B[2]), .QN(n10) );
  NAND2X1 U12 ( .IN1(A[2]), .IN2(carry[2]), .QN(n11) );
  NAND3X0 U13 ( .IN1(n9), .IN2(n11), .IN3(n10), .QN(carry[3]) );
  AND2X1 U14 ( .IN1(A[0]), .IN2(B[0]), .Q(n12) );
  XOR2X1 U15 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_1 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_1_DW01_add_0 add_37 ( .A(a), .B({
        b[11:3], n6, b[1:0]}), .CI(1'b0), .SUM(pre_out) );
  INVX0 U2 ( .INP(b[11]), .ZN(n12) );
  DELLN1X2 U3 ( .INP(pre_out[11]), .Z(n1) );
  AND2X1 U4 ( .IN1(n11), .IN2(n10), .Q(n2) );
  AND2X1 U5 ( .IN1(n2), .IN2(n12), .Q(n8) );
  NAND2X1 U6 ( .IN1(n11), .IN2(n10), .QN(n4) );
  INVX0 U7 ( .INP(b[2]), .ZN(n5) );
  INVX0 U8 ( .INP(n5), .ZN(n6) );
  AND2X1 U9 ( .IN1(n2), .IN2(n12), .Q(n7) );
  AND2X1 U10 ( .IN1(n2), .IN2(n12), .Q(n9) );
  MUX21X2 U11 ( .IN1(n1), .IN2(b[11]), .S(n2), .Q(\output [11]) );
  XOR2X1 U12 ( .IN1(n12), .IN2(a[11]), .Q(n11) );
  XOR2X1 U13 ( .IN1(a[11]), .IN2(pre_out[11]), .Q(n10) );
  AO21X1 U14 ( .IN1(pre_out[0]), .IN2(n4), .IN3(n8), .Q(\output [0]) );
  AO21X1 U15 ( .IN1(pre_out[1]), .IN2(n4), .IN3(n7), .Q(\output [1]) );
  AO21X1 U16 ( .IN1(pre_out[2]), .IN2(n4), .IN3(n8), .Q(\output [2]) );
  AO21X1 U17 ( .IN1(pre_out[3]), .IN2(n4), .IN3(n7), .Q(\output [3]) );
  AO21X1 U18 ( .IN1(pre_out[4]), .IN2(n4), .IN3(n8), .Q(\output [4]) );
  AO21X1 U19 ( .IN1(pre_out[5]), .IN2(n4), .IN3(n7), .Q(\output [5]) );
  AO21X1 U20 ( .IN1(pre_out[6]), .IN2(n4), .IN3(n9), .Q(\output [6]) );
  AO21X1 U21 ( .IN1(pre_out[7]), .IN2(n4), .IN3(n9), .Q(\output [7]) );
  AO21X1 U22 ( .IN1(pre_out[8]), .IN2(n4), .IN3(n9), .Q(\output [8]) );
  AO21X1 U23 ( .IN1(pre_out[9]), .IN2(n4), .IN3(n7), .Q(\output [9]) );
  AO21X1 U24 ( .IN1(pre_out[10]), .IN2(n4), .IN3(n9), .Q(\output [10]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_0_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [11:1] carry;

  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_11 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(SUM[11]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_0 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n7, n8;
  wire   [11:0] pre_out;

  AO21X1 U6 ( .IN1(pre_out[9]), .IN2(n8), .IN3(n7), .Q(\output [9]) );
  AO21X1 U7 ( .IN1(pre_out[8]), .IN2(n8), .IN3(n7), .Q(\output [8]) );
  AO21X1 U8 ( .IN1(pre_out[7]), .IN2(n8), .IN3(n7), .Q(\output [7]) );
  AO21X1 U9 ( .IN1(pre_out[6]), .IN2(n8), .IN3(n7), .Q(\output [6]) );
  AO21X1 U10 ( .IN1(pre_out[5]), .IN2(n8), .IN3(n7), .Q(\output [5]) );
  AO21X1 U11 ( .IN1(pre_out[4]), .IN2(n8), .IN3(n7), .Q(\output [4]) );
  AO21X1 U12 ( .IN1(pre_out[3]), .IN2(n8), .IN3(n7), .Q(\output [3]) );
  AO21X1 U13 ( .IN1(pre_out[2]), .IN2(n8), .IN3(n7), .Q(\output [2]) );
  AO21X1 U14 ( .IN1(pre_out[1]), .IN2(n8), .IN3(n7), .Q(\output [1]) );
  AO22X1 U15 ( .IN1(n1), .IN2(b[11]), .IN3(pre_out[11]), .IN4(n8), .Q(
        \output [11]) );
  AO21X1 U16 ( .IN1(pre_out[10]), .IN2(n8), .IN3(n7), .Q(\output [10]) );
  AO21X1 U17 ( .IN1(pre_out[0]), .IN2(n8), .IN3(n7), .Q(\output [0]) );
  XOR2X1 U18 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n2) );
  XNOR2X1 U19 ( .IN1(a[11]), .IN2(b[11]), .Q(n4) );
  add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_0_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(pre_out) );
  NOR2X0 U2 ( .IN1(n8), .IN2(b[11]), .QN(n7) );
  NAND2X1 U3 ( .IN1(n4), .IN2(n2), .QN(n8) );
  INVX0 U4 ( .INP(n8), .ZN(n1) );
endmodule


module inner_prod_INT_BITS4_WORD_WIDTH12_N4 ( clk, rst, in_a_r, in_a_i, in_b_r, 
        in_b_i, out_r, out_i, reduced_matrix, start, done );
  input [11:0] in_a_r;
  input [11:0] in_a_i;
  input [11:0] in_b_r;
  input [11:0] in_b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk, rst, reduced_matrix, start;
  output done;
  wire   in_reg_enable_fsm, acc_clear, acc_enable, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, n91, n93, n95, n96, n97, n98, n101, n102, n103, n104, n105, n106,
         n107, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37;
  wire   [2:0] in_counter;
  wire   [1:0] state;
  wire   [2:0] pipe_counter;
  wire   [11:0] in_a_r_reg;
  wire   [11:0] in_a_i_reg;
  wire   [11:0] in_b_r_reg;
  wire   [11:0] in_b_i_reg;
  wire   [11:0] add_r_out;
  wire   [11:0] add_i_out;
  wire   [11:0] mult_out_r;
  wire   [11:0] mult_out_i;

  DFFARX1 \pipe_counter_reg[0]  ( .D(n144), .CLK(clk), .RSTB(n19), .Q(
        pipe_counter[0]) );
  DFFARX1 \pipe_counter_reg[1]  ( .D(n134), .CLK(clk), .RSTB(n19), .Q(
        pipe_counter[1]) );
  DFFARX1 \pipe_counter_reg[2]  ( .D(n143), .CLK(clk), .RSTB(n19), .Q(
        pipe_counter[2]) );
  DFFARX1 \state_reg[0]  ( .D(n141), .CLK(clk), .RSTB(n19), .Q(state[0]) );
  DFFARX1 \state_reg[1]  ( .D(n142), .CLK(clk), .RSTB(n19), .Q(state[1]), .QN(
        n91) );
  DFFARX1 acc_enable_reg ( .D(n133), .CLK(clk), .RSTB(n25), .Q(acc_enable), 
        .QN(n93) );
  DFFARX1 \in_counter_reg[0]  ( .D(n138), .CLK(clk), .RSTB(n19), .Q(
        in_counter[0]) );
  DFFARX1 \in_counter_reg[1]  ( .D(n137), .CLK(clk), .RSTB(n19), .Q(
        in_counter[1]) );
  DFFARX1 \in_counter_reg[2]  ( .D(n136), .CLK(clk), .RSTB(n19), .Q(
        in_counter[2]) );
  DFFARX1 in_reg_enable_fsm_reg ( .D(n135), .CLK(clk), .RSTB(n24), .Q(
        in_reg_enable_fsm) );
  DFFASX1 acc_clear_reg ( .D(n139), .CLK(clk), .SETB(n25), .Q(acc_clear), .QN(
        n1) );
  DFFARX1 done_reg ( .D(n140), .CLK(clk), .RSTB(n19), .Q(done) );
  DFFARX1 \in_b_i_reg_reg[11]  ( .D(N80), .CLK(clk), .RSTB(n23), .Q(
        in_b_i_reg[11]) );
  DFFARX1 \in_b_i_reg_reg[10]  ( .D(N79), .CLK(clk), .RSTB(n23), .Q(
        in_b_i_reg[10]) );
  DFFARX1 \in_b_i_reg_reg[9]  ( .D(N78), .CLK(clk), .RSTB(n23), .Q(
        in_b_i_reg[9]) );
  DFFARX1 \in_b_i_reg_reg[8]  ( .D(N77), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[8]) );
  DFFARX1 \in_b_i_reg_reg[7]  ( .D(N76), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[7]) );
  DFFARX1 \in_b_i_reg_reg[6]  ( .D(N75), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[6]) );
  DFFARX1 \in_b_i_reg_reg[5]  ( .D(N74), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[5]) );
  DFFARX1 \in_b_i_reg_reg[4]  ( .D(N73), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[4]) );
  DFFARX1 \in_b_i_reg_reg[3]  ( .D(N72), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[3]) );
  DFFARX1 \in_b_i_reg_reg[2]  ( .D(N71), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[2]) );
  DFFARX1 \in_b_i_reg_reg[1]  ( .D(N70), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[1]) );
  DFFARX1 \in_b_i_reg_reg[0]  ( .D(N69), .CLK(clk), .RSTB(n24), .Q(
        in_b_i_reg[0]) );
  DFFARX1 \in_a_r_reg_reg[11]  ( .D(N44), .CLK(clk), .RSTB(n20), .Q(
        in_a_r_reg[11]) );
  DFFARX1 \in_a_r_reg_reg[10]  ( .D(N43), .CLK(clk), .RSTB(n20), .Q(
        in_a_r_reg[10]) );
  DFFARX1 \in_a_r_reg_reg[9]  ( .D(N42), .CLK(clk), .RSTB(n20), .Q(
        in_a_r_reg[9]) );
  DFFARX1 \in_a_r_reg_reg[8]  ( .D(N41), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[8]) );
  DFFARX1 \in_a_r_reg_reg[7]  ( .D(N40), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[7]) );
  DFFARX1 \in_a_r_reg_reg[6]  ( .D(N39), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[6]) );
  DFFARX1 \in_a_r_reg_reg[5]  ( .D(N38), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[5]) );
  DFFARX1 \in_a_r_reg_reg[4]  ( .D(N37), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[4]) );
  DFFARX1 \in_a_r_reg_reg[3]  ( .D(N36), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[3]) );
  DFFARX1 \in_a_r_reg_reg[2]  ( .D(N35), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[2]) );
  DFFARX1 \in_a_r_reg_reg[1]  ( .D(N34), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[1]) );
  DFFARX1 \in_a_r_reg_reg[0]  ( .D(N33), .CLK(clk), .RSTB(n21), .Q(
        in_a_r_reg[0]) );
  DFFARX1 \in_a_i_reg_reg[11]  ( .D(N56), .CLK(clk), .RSTB(n21), .Q(
        in_a_i_reg[11]) );
  DFFARX1 \in_a_i_reg_reg[10]  ( .D(N55), .CLK(clk), .RSTB(n21), .Q(
        in_a_i_reg[10]) );
  DFFARX1 \in_a_i_reg_reg[9]  ( .D(N54), .CLK(clk), .RSTB(n21), .Q(
        in_a_i_reg[9]) );
  DFFARX1 \in_a_i_reg_reg[8]  ( .D(N53), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[8]) );
  DFFARX1 \in_a_i_reg_reg[7]  ( .D(N52), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[7]) );
  DFFARX1 \in_a_i_reg_reg[6]  ( .D(N51), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[6]) );
  DFFARX1 \in_a_i_reg_reg[5]  ( .D(N50), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[5]) );
  DFFARX1 \in_a_i_reg_reg[4]  ( .D(N49), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[4]) );
  DFFARX1 \in_a_i_reg_reg[3]  ( .D(N48), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[3]) );
  DFFARX1 \in_a_i_reg_reg[2]  ( .D(N47), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[2]) );
  DFFARX1 \in_a_i_reg_reg[1]  ( .D(N46), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[1]) );
  DFFARX1 \in_a_i_reg_reg[0]  ( .D(N45), .CLK(clk), .RSTB(n22), .Q(
        in_a_i_reg[0]) );
  DFFARX1 \in_b_r_reg_reg[11]  ( .D(N68), .CLK(clk), .RSTB(n22), .Q(
        in_b_r_reg[11]) );
  DFFARX1 \in_b_r_reg_reg[10]  ( .D(N67), .CLK(clk), .RSTB(n22), .Q(
        in_b_r_reg[10]) );
  DFFARX1 \in_b_r_reg_reg[9]  ( .D(N66), .CLK(clk), .RSTB(n22), .Q(
        in_b_r_reg[9]) );
  DFFARX1 \in_b_r_reg_reg[8]  ( .D(N65), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[8]) );
  DFFARX1 \in_b_r_reg_reg[7]  ( .D(N64), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[7]) );
  DFFARX1 \in_b_r_reg_reg[6]  ( .D(N63), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[6]) );
  DFFARX1 \in_b_r_reg_reg[5]  ( .D(N62), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[5]) );
  DFFARX1 \in_b_r_reg_reg[4]  ( .D(N61), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[4]) );
  DFFARX1 \in_b_r_reg_reg[3]  ( .D(N60), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[3]) );
  DFFARX1 \in_b_r_reg_reg[2]  ( .D(N59), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[2]) );
  DFFARX1 \in_b_r_reg_reg[1]  ( .D(N58), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[1]) );
  DFFARX1 \in_b_r_reg_reg[0]  ( .D(N57), .CLK(clk), .RSTB(n23), .Q(
        in_b_r_reg[0]) );
  DFFARX1 \acc_i_reg[0]  ( .D(n132), .CLK(clk), .RSTB(n19), .Q(out_i[0]) );
  DFFARX1 \acc_i_reg[1]  ( .D(n131), .CLK(clk), .RSTB(n19), .Q(out_i[1]) );
  DFFARX1 \acc_i_reg[2]  ( .D(n130), .CLK(clk), .RSTB(n19), .Q(out_i[2]) );
  DFFARX1 \acc_i_reg[3]  ( .D(n129), .CLK(clk), .RSTB(n20), .Q(out_i[3]) );
  DFFARX1 \acc_i_reg[4]  ( .D(n128), .CLK(clk), .RSTB(n20), .Q(out_i[4]) );
  DFFARX1 \acc_i_reg[5]  ( .D(n127), .CLK(clk), .RSTB(n20), .Q(out_i[5]) );
  DFFARX1 \acc_i_reg[6]  ( .D(n126), .CLK(clk), .RSTB(n20), .Q(out_i[6]) );
  DFFARX1 \acc_i_reg[7]  ( .D(n125), .CLK(clk), .RSTB(n20), .Q(out_i[7]) );
  DFFARX1 \acc_i_reg[8]  ( .D(n124), .CLK(clk), .RSTB(n20), .Q(out_i[8]) );
  DFFARX1 \acc_i_reg[9]  ( .D(n123), .CLK(clk), .RSTB(n20), .Q(out_i[9]) );
  DFFARX1 \acc_i_reg[10]  ( .D(n122), .CLK(clk), .RSTB(n20), .Q(out_i[10]) );
  DFFARX1 \acc_i_reg[11]  ( .D(n121), .CLK(clk), .RSTB(n20), .Q(out_i[11]) );
  DFFARX1 \acc_r_reg[0]  ( .D(n120), .CLK(clk), .RSTB(n25), .Q(out_r[0]) );
  DFFARX1 \acc_r_reg[1]  ( .D(n119), .CLK(clk), .RSTB(n25), .Q(out_r[1]), .QN(
        n8) );
  DFFARX1 \acc_r_reg[2]  ( .D(n118), .CLK(clk), .RSTB(n25), .Q(out_r[2]) );
  DFFARX1 \acc_r_reg[3]  ( .D(n117), .CLK(clk), .RSTB(n25), .Q(out_r[3]), .QN(
        n6) );
  DFFARX1 \acc_r_reg[4]  ( .D(n116), .CLK(clk), .RSTB(n25), .Q(out_r[4]) );
  DFFARX1 \acc_r_reg[5]  ( .D(n115), .CLK(clk), .RSTB(n25), .Q(out_r[5]) );
  DFFARX1 \acc_r_reg[6]  ( .D(n114), .CLK(clk), .RSTB(n25), .Q(out_r[6]), .QN(
        n4) );
  DFFARX1 \acc_r_reg[7]  ( .D(n113), .CLK(clk), .RSTB(n25), .Q(out_r[7]), .QN(
        n2) );
  DFFARX1 \acc_r_reg[8]  ( .D(n112), .CLK(clk), .RSTB(n25), .Q(out_r[8]) );
  DFFARX1 \acc_r_reg[9]  ( .D(n111), .CLK(clk), .RSTB(n25), .Q(out_r[9]) );
  DFFARX1 \acc_r_reg[10]  ( .D(n110), .CLK(clk), .RSTB(n24), .Q(out_r[10]) );
  DFFARX1 \acc_r_reg[11]  ( .D(n109), .CLK(clk), .RSTB(n24), .Q(out_r[11]) );
  AO22X1 U105 ( .IN1(done), .IN2(n36), .IN3(pipe_counter[2]), .IN4(n95), .Q(
        n140) );
  AO22X1 U106 ( .IN1(n96), .IN2(n97), .IN3(n30), .IN4(state[0]), .Q(n141) );
  AO22X1 U107 ( .IN1(n37), .IN2(n97), .IN3(n30), .IN4(state[1]), .Q(n142) );
  AO21X1 U108 ( .IN1(pipe_counter[2]), .IN2(n95), .IN3(n31), .Q(n97) );
  AO22X1 U109 ( .IN1(n33), .IN2(pipe_counter[2]), .IN3(pipe_counter[1]), .IN4(
        n95), .Q(n143) );
  AO22X1 U110 ( .IN1(n37), .IN2(n98), .IN3(pipe_counter[0]), .IN4(n33), .Q(
        n144) );
  AO22X1 U123 ( .IN1(out_i[11]), .IN2(n17), .IN3(add_i_out[11]), .IN4(n15), 
        .Q(n121) );
  AO22X1 U124 ( .IN1(out_i[10]), .IN2(n17), .IN3(add_i_out[10]), .IN4(n15), 
        .Q(n122) );
  AO22X1 U125 ( .IN1(out_i[9]), .IN2(n17), .IN3(add_i_out[9]), .IN4(n15), .Q(
        n123) );
  AO22X1 U126 ( .IN1(out_i[8]), .IN2(n17), .IN3(add_i_out[8]), .IN4(n15), .Q(
        n124) );
  AO22X1 U127 ( .IN1(out_i[7]), .IN2(n17), .IN3(add_i_out[7]), .IN4(n15), .Q(
        n125) );
  AO22X1 U128 ( .IN1(out_i[6]), .IN2(n17), .IN3(add_i_out[6]), .IN4(n15), .Q(
        n126) );
  AO22X1 U129 ( .IN1(out_i[5]), .IN2(n17), .IN3(add_i_out[5]), .IN4(n15), .Q(
        n127) );
  AO22X1 U130 ( .IN1(out_i[4]), .IN2(n17), .IN3(add_i_out[4]), .IN4(n15), .Q(
        n128) );
  AO22X1 U131 ( .IN1(out_i[3]), .IN2(n17), .IN3(add_i_out[3]), .IN4(n15), .Q(
        n129) );
  AO22X1 U132 ( .IN1(out_i[2]), .IN2(n17), .IN3(add_i_out[2]), .IN4(n15), .Q(
        n130) );
  AO22X1 U133 ( .IN1(out_i[1]), .IN2(n17), .IN3(add_i_out[1]), .IN4(n15), .Q(
        n131) );
  AO22X1 U134 ( .IN1(out_i[0]), .IN2(n17), .IN3(add_i_out[0]), .IN4(n15), .Q(
        n132) );
  AO21X1 U135 ( .IN1(pipe_counter[2]), .IN2(n95), .IN3(n93), .Q(n102) );
  AO22X1 U136 ( .IN1(n33), .IN2(pipe_counter[1]), .IN3(pipe_counter[0]), .IN4(
        n95), .Q(n134) );
  AO21X1 U137 ( .IN1(n37), .IN2(n103), .IN3(n95), .Q(n98) );
  AO22X1 U139 ( .IN1(in_counter[2]), .IN2(n34), .IN3(reduced_matrix), .IN4(
        in_counter[0]), .Q(n103) );
  AO22X1 U140 ( .IN1(n35), .IN2(in_counter[2]), .IN3(in_counter[1]), .IN4(n37), 
        .Q(n136) );
  AO22X1 U141 ( .IN1(n35), .IN2(in_counter[1]), .IN3(n37), .IN4(in_counter[0]), 
        .Q(n137) );
  AO22X1 U142 ( .IN1(n96), .IN2(n106), .IN3(n35), .IN4(in_counter[0]), .Q(n138) );
  NAND3X0 U143 ( .IN1(n101), .IN2(n36), .IN3(acc_clear), .QN(n107) );
  complex_mult_pipe_prod_INT_BITS4_WORD_WIDTH12 cp_mult ( .a_r(in_a_r_reg), 
        .a_i(in_a_i_reg), .b_r(in_b_r_reg), .b_i(in_b_i_reg), .out_r(
        mult_out_r), .out_i(mult_out_i), .clk(clk) );
  add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_1 add_r ( .a(mult_out_r), .b({
        out_r[11:8], n3, out_r[6:4], n7, out_r[2], n9, out_r[0]}), .\output (
        add_r_out) );
  add_sub_WORD_WIDTH12_OPERATION1_USE_SAT1_0 add_i ( .a(mult_out_i), .b(out_i), 
        .\output (add_i_out) );
  INVX0 U3 ( .INP(n2), .ZN(n3) );
  INVX0 U4 ( .INP(n8), .ZN(n9) );
  INVX0 U5 ( .INP(n4), .ZN(n5) );
  INVX0 U6 ( .INP(n6), .ZN(n7) );
  NBUFFX2 U7 ( .INP(n28), .Z(n18) );
  NBUFFX2 U8 ( .INP(n28), .Z(n17) );
  INVX0 U9 ( .INP(n98), .ZN(n33) );
  INVX0 U10 ( .INP(n106), .ZN(n35) );
  INVX0 U11 ( .INP(n104), .ZN(n31) );
  NBUFFX2 U12 ( .INP(n10), .Z(n16) );
  NBUFFX2 U13 ( .INP(n10), .Z(n15) );
  NBUFFX2 U14 ( .INP(n27), .Z(n13) );
  NBUFFX2 U15 ( .INP(n27), .Z(n12) );
  NBUFFX2 U16 ( .INP(n27), .Z(n11) );
  NBUFFX2 U17 ( .INP(n27), .Z(n14) );
  INVX0 U18 ( .INP(n101), .ZN(n37) );
  OA21X1 U19 ( .IN1(n101), .IN2(n32), .IN3(n105), .Q(n104) );
  INVX0 U20 ( .INP(n103), .ZN(n32) );
  NAND2X1 U21 ( .IN1(n101), .IN2(n105), .QN(n106) );
  INVX0 U22 ( .INP(n96), .ZN(n36) );
  INVX0 U23 ( .INP(n26), .ZN(n28) );
  INVX0 U24 ( .INP(n97), .ZN(n30) );
  NBUFFX2 U25 ( .INP(n29), .Z(n22) );
  NBUFFX2 U26 ( .INP(n29), .Z(n21) );
  NBUFFX2 U27 ( .INP(n29), .Z(n20) );
  NBUFFX2 U28 ( .INP(n29), .Z(n23) );
  NBUFFX2 U29 ( .INP(n29), .Z(n24) );
  NBUFFX2 U30 ( .INP(n29), .Z(n19) );
  NBUFFX2 U31 ( .INP(n29), .Z(n25) );
  NOR2X0 U32 ( .IN1(state[0]), .IN2(state[1]), .QN(n96) );
  OR2X1 U33 ( .IN1(in_reg_enable_fsm), .IN2(start), .Q(n27) );
  NAND2X1 U34 ( .IN1(state[0]), .IN2(n91), .QN(n101) );
  NOR2X0 U35 ( .IN1(n91), .IN2(state[0]), .QN(n95) );
  NAND2X0 U36 ( .IN1(start), .IN2(n96), .QN(n105) );
  INVX0 U37 ( .INP(reduced_matrix), .ZN(n34) );
  NAND2X0 U38 ( .IN1(n105), .IN2(n107), .QN(n139) );
  AND2X1 U39 ( .IN1(n26), .IN2(n1), .Q(n10) );
  NAND2X1 U40 ( .IN1(n101), .IN2(n102), .QN(n133) );
  INVX0 U41 ( .INP(rst), .ZN(n29) );
  OR2X1 U42 ( .IN1(acc_enable), .IN2(acc_clear), .Q(n26) );
  AO22X1 U43 ( .IN1(out_r[0]), .IN2(n18), .IN3(add_r_out[0]), .IN4(n16), .Q(
        n120) );
  AO22X1 U44 ( .IN1(n9), .IN2(n18), .IN3(add_r_out[1]), .IN4(n16), .Q(n119) );
  AO22X1 U45 ( .IN1(out_r[2]), .IN2(n18), .IN3(add_r_out[2]), .IN4(n16), .Q(
        n118) );
  AO22X1 U46 ( .IN1(n7), .IN2(n18), .IN3(add_r_out[3]), .IN4(n16), .Q(n117) );
  AO22X1 U47 ( .IN1(out_r[4]), .IN2(n18), .IN3(add_r_out[4]), .IN4(n16), .Q(
        n116) );
  AO22X1 U48 ( .IN1(out_r[5]), .IN2(n18), .IN3(add_r_out[5]), .IN4(n16), .Q(
        n115) );
  AO22X1 U49 ( .IN1(n5), .IN2(n18), .IN3(add_r_out[6]), .IN4(n16), .Q(n114) );
  AO22X1 U50 ( .IN1(n3), .IN2(n18), .IN3(add_r_out[7]), .IN4(n16), .Q(n113) );
  AO22X1 U51 ( .IN1(out_r[8]), .IN2(n18), .IN3(add_r_out[8]), .IN4(n16), .Q(
        n112) );
  AO22X1 U52 ( .IN1(out_r[9]), .IN2(n18), .IN3(add_r_out[9]), .IN4(n16), .Q(
        n111) );
  AO22X1 U53 ( .IN1(out_r[10]), .IN2(n18), .IN3(add_r_out[10]), .IN4(n16), .Q(
        n110) );
  AO22X1 U54 ( .IN1(out_r[11]), .IN2(n18), .IN3(add_r_out[11]), .IN4(n16), .Q(
        n109) );
  AO22X1 U55 ( .IN1(n31), .IN2(n96), .IN3(n104), .IN4(in_reg_enable_fsm), .Q(
        n135) );
  AND2X1 U56 ( .IN1(in_b_i[0]), .IN2(n14), .Q(N69) );
  AND2X1 U57 ( .IN1(in_b_i[1]), .IN2(n14), .Q(N70) );
  AND2X1 U58 ( .IN1(in_b_i[2]), .IN2(n14), .Q(N71) );
  AND2X1 U59 ( .IN1(in_b_i[3]), .IN2(n14), .Q(N72) );
  AND2X1 U60 ( .IN1(in_b_i[4]), .IN2(n14), .Q(N73) );
  AND2X1 U61 ( .IN1(in_b_i[5]), .IN2(n14), .Q(N74) );
  AND2X1 U62 ( .IN1(in_b_i[6]), .IN2(n14), .Q(N75) );
  AND2X1 U63 ( .IN1(in_b_i[7]), .IN2(n14), .Q(N76) );
  AND2X1 U64 ( .IN1(in_b_i[8]), .IN2(n14), .Q(N77) );
  AND2X1 U65 ( .IN1(in_b_i[9]), .IN2(n14), .Q(N78) );
  AND2X1 U66 ( .IN1(in_b_i[10]), .IN2(n14), .Q(N79) );
  AND2X1 U67 ( .IN1(in_b_i[11]), .IN2(n14), .Q(N80) );
  AND2X1 U68 ( .IN1(in_b_r[0]), .IN2(n13), .Q(N57) );
  AND2X1 U69 ( .IN1(in_b_r[1]), .IN2(n13), .Q(N58) );
  AND2X1 U70 ( .IN1(in_b_r[2]), .IN2(n13), .Q(N59) );
  AND2X1 U71 ( .IN1(in_b_r[3]), .IN2(n13), .Q(N60) );
  AND2X1 U72 ( .IN1(in_b_r[4]), .IN2(n13), .Q(N61) );
  AND2X1 U73 ( .IN1(in_b_r[5]), .IN2(n13), .Q(N62) );
  AND2X1 U74 ( .IN1(in_b_r[6]), .IN2(n13), .Q(N63) );
  AND2X1 U75 ( .IN1(in_b_r[7]), .IN2(n13), .Q(N64) );
  AND2X1 U76 ( .IN1(in_b_r[8]), .IN2(n13), .Q(N65) );
  AND2X1 U77 ( .IN1(in_b_r[9]), .IN2(n13), .Q(N66) );
  AND2X1 U78 ( .IN1(in_b_r[10]), .IN2(n13), .Q(N67) );
  AND2X1 U79 ( .IN1(in_b_r[11]), .IN2(n13), .Q(N68) );
  AND2X1 U80 ( .IN1(in_a_i[0]), .IN2(n12), .Q(N45) );
  AND2X1 U81 ( .IN1(in_a_i[1]), .IN2(n12), .Q(N46) );
  AND2X1 U82 ( .IN1(in_a_i[2]), .IN2(n12), .Q(N47) );
  AND2X1 U83 ( .IN1(in_a_i[3]), .IN2(n12), .Q(N48) );
  AND2X1 U84 ( .IN1(in_a_i[4]), .IN2(n12), .Q(N49) );
  AND2X1 U85 ( .IN1(in_a_i[5]), .IN2(n12), .Q(N50) );
  AND2X1 U86 ( .IN1(in_a_i[6]), .IN2(n12), .Q(N51) );
  AND2X1 U87 ( .IN1(in_a_i[7]), .IN2(n12), .Q(N52) );
  AND2X1 U88 ( .IN1(in_a_i[8]), .IN2(n12), .Q(N53) );
  AND2X1 U89 ( .IN1(in_a_i[9]), .IN2(n12), .Q(N54) );
  AND2X1 U90 ( .IN1(in_a_i[10]), .IN2(n12), .Q(N55) );
  AND2X1 U91 ( .IN1(in_a_i[11]), .IN2(n12), .Q(N56) );
  AND2X1 U92 ( .IN1(in_a_r[0]), .IN2(n11), .Q(N33) );
  AND2X1 U93 ( .IN1(in_a_r[1]), .IN2(n11), .Q(N34) );
  AND2X1 U94 ( .IN1(in_a_r[2]), .IN2(n11), .Q(N35) );
  AND2X1 U95 ( .IN1(in_a_r[3]), .IN2(n11), .Q(N36) );
  AND2X1 U96 ( .IN1(in_a_r[4]), .IN2(n11), .Q(N37) );
  AND2X1 U97 ( .IN1(in_a_r[5]), .IN2(n11), .Q(N38) );
  AND2X1 U98 ( .IN1(in_a_r[6]), .IN2(n11), .Q(N39) );
  AND2X1 U99 ( .IN1(in_a_r[7]), .IN2(n11), .Q(N40) );
  AND2X1 U100 ( .IN1(in_a_r[8]), .IN2(n11), .Q(N41) );
  AND2X1 U101 ( .IN1(in_a_r[9]), .IN2(n11), .Q(N42) );
  AND2X1 U102 ( .IN1(in_a_r[10]), .IN2(n11), .Q(N43) );
  AND2X1 U103 ( .IN1(in_a_r[11]), .IN2(n11), .Q(N44) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_15_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560;

  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n459), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n461), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n463), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n465), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  XOR3X1 U311 ( .IN1(n27), .IN2(n457), .IN3(n412), .Q(product[21]) );
  DELLN2X2 U312 ( .INP(n18), .Z(n408) );
  INVX0 U313 ( .INP(b[3]), .ZN(n409) );
  INVX0 U314 ( .INP(n409), .ZN(n410) );
  INVX0 U315 ( .INP(n5), .ZN(n411) );
  INVX0 U316 ( .INP(n411), .ZN(n412) );
  INVX0 U317 ( .INP(b[2]), .ZN(n413) );
  INVX0 U318 ( .INP(n413), .ZN(n414) );
  INVX0 U319 ( .INP(b[1]), .ZN(n415) );
  INVX0 U320 ( .INP(n415), .ZN(n416) );
  XOR2X2 U321 ( .IN1(b[10]), .IN2(n456), .Q(n486) );
  XOR2X2 U322 ( .IN1(b[10]), .IN2(n454), .Q(n483) );
  XOR2X2 U323 ( .IN1(b[10]), .IN2(n452), .Q(n480) );
  XOR2X2 U324 ( .IN1(b[10]), .IN2(n450), .Q(n477) );
  XOR2X2 U325 ( .IN1(b[10]), .IN2(n448), .Q(n469) );
  XOR2X2 U326 ( .IN1(b[10]), .IN2(n443), .Q(n496) );
  XOR2X2 U327 ( .IN1(b[8]), .IN2(n456), .Q(n549) );
  XOR2X2 U328 ( .IN1(b[8]), .IN2(n454), .Q(n538) );
  XOR2X2 U329 ( .IN1(b[8]), .IN2(n452), .Q(n527) );
  XOR2X2 U330 ( .IN1(b[8]), .IN2(n450), .Q(n516) );
  XOR2X2 U331 ( .IN1(b[8]), .IN2(n448), .Q(n506) );
  XOR2X2 U332 ( .IN1(b[8]), .IN2(n443), .Q(n494) );
  XOR2X2 U333 ( .IN1(b[6]), .IN2(n456), .Q(n547) );
  XOR2X2 U334 ( .IN1(b[6]), .IN2(n454), .Q(n536) );
  XOR2X2 U335 ( .IN1(b[6]), .IN2(n452), .Q(n525) );
  XOR2X2 U336 ( .IN1(b[6]), .IN2(n450), .Q(n514) );
  XOR2X2 U337 ( .IN1(b[6]), .IN2(n448), .Q(n504) );
  XOR2X2 U338 ( .IN1(b[6]), .IN2(n443), .Q(n492) );
  XOR2X2 U339 ( .IN1(b[5]), .IN2(n456), .Q(n546) );
  XOR2X2 U340 ( .IN1(b[5]), .IN2(n454), .Q(n535) );
  XOR2X2 U341 ( .IN1(b[5]), .IN2(n452), .Q(n524) );
  XOR2X2 U342 ( .IN1(b[5]), .IN2(n450), .Q(n513) );
  XOR2X2 U343 ( .IN1(b[5]), .IN2(n448), .Q(n503) );
  XOR2X2 U344 ( .IN1(b[5]), .IN2(n443), .Q(n491) );
  XOR2X1 U345 ( .IN1(n417), .IN2(n4), .Q(product[22]) );
  XOR2X1 U346 ( .IN1(n25), .IN2(n153), .Q(n417) );
  XNOR2X1 U347 ( .IN1(n418), .IN2(n408), .Q(product[8]) );
  XNOR2X1 U348 ( .IN1(n112), .IN2(n117), .Q(n418) );
  AND3X1 U349 ( .IN1(n431), .IN2(n432), .IN3(n433), .Q(product[23]) );
  INVX0 U350 ( .INP(n55), .ZN(n463) );
  XOR3X1 U351 ( .IN1(n33), .IN2(n30), .IN3(n7), .Q(product[19]) );
  XNOR2X1 U352 ( .IN1(n420), .IN2(n6), .Q(product[20]) );
  XNOR2X1 U353 ( .IN1(n29), .IN2(n28), .Q(n420) );
  INVX0 U354 ( .INP(n25), .ZN(n457) );
  XOR3X1 U355 ( .IN1(n118), .IN2(n123), .IN3(n19), .Q(product[7]) );
  XOR2X1 U356 ( .IN1(n416), .IN2(n443), .Q(n487) );
  XOR2X1 U357 ( .IN1(n410), .IN2(n443), .Q(n489) );
  XOR2X1 U358 ( .IN1(n416), .IN2(n448), .Q(n498) );
  XOR2X1 U359 ( .IN1(n416), .IN2(n450), .Q(n508) );
  XOR2X1 U360 ( .IN1(n410), .IN2(n448), .Q(n501) );
  INVX0 U361 ( .INP(n73), .ZN(n465) );
  XOR2X1 U362 ( .IN1(n416), .IN2(n452), .Q(n519) );
  XOR2X1 U363 ( .IN1(n416), .IN2(n454), .Q(n530) );
  XOR2X1 U364 ( .IN1(n416), .IN2(n456), .Q(n541) );
  XOR2X1 U365 ( .IN1(n410), .IN2(n450), .Q(n511) );
  XOR2X1 U366 ( .IN1(n410), .IN2(n452), .Q(n522) );
  XOR2X1 U367 ( .IN1(n410), .IN2(n454), .Q(n533) );
  INVX0 U368 ( .INP(n41), .ZN(n461) );
  XOR2X1 U369 ( .IN1(n410), .IN2(n456), .Q(n544) );
  INVX0 U370 ( .INP(n31), .ZN(n459) );
  NBUFFX2 U371 ( .INP(a[1]), .Z(n443) );
  INVX0 U372 ( .INP(n497), .ZN(n466) );
  AND2X1 U373 ( .IN1(n443), .IN2(n447), .Q(n472) );
  XNOR2X1 U374 ( .IN1(n421), .IN2(n20), .Q(product[6]) );
  XNOR2X1 U375 ( .IN1(n127), .IN2(n124), .Q(n421) );
  INVX0 U376 ( .INP(n507), .ZN(n464) );
  INVX0 U377 ( .INP(n518), .ZN(n462) );
  INVX0 U378 ( .INP(n529), .ZN(n460) );
  INVX0 U379 ( .INP(n540), .ZN(n458) );
  NBUFFX2 U380 ( .INP(a[3]), .Z(n449) );
  FADDX1 U381 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  NBUFFX2 U382 ( .INP(a[5]), .Z(n451) );
  AND2X1 U383 ( .IN1(n497), .IN2(n552), .Q(n470) );
  AND2X1 U384 ( .IN1(n518), .IN2(n556), .Q(n479) );
  AND2X1 U385 ( .IN1(n507), .IN2(n554), .Q(n476) );
  AND2X1 U386 ( .IN1(n529), .IN2(n558), .Q(n482) );
  AND2X1 U387 ( .IN1(n540), .IN2(n560), .Q(n485) );
  NBUFFX2 U388 ( .INP(a[7]), .Z(n453) );
  NBUFFX2 U389 ( .INP(a[9]), .Z(n455) );
  NAND2X0 U390 ( .IN1(n33), .IN2(n30), .QN(n422) );
  NAND2X0 U391 ( .IN1(n33), .IN2(n7), .QN(n423) );
  NAND2X0 U392 ( .IN1(n30), .IN2(n7), .QN(n424) );
  NAND3X0 U393 ( .IN1(n422), .IN2(n423), .IN3(n424), .QN(n6) );
  NAND2X0 U394 ( .IN1(n29), .IN2(n28), .QN(n425) );
  NAND2X0 U395 ( .IN1(n29), .IN2(n6), .QN(n426) );
  NAND2X0 U396 ( .IN1(n28), .IN2(n6), .QN(n427) );
  NAND3X0 U397 ( .IN1(n425), .IN2(n426), .IN3(n427), .QN(n5) );
  NAND2X1 U398 ( .IN1(n27), .IN2(n457), .QN(n428) );
  NAND2X0 U399 ( .IN1(n27), .IN2(n5), .QN(n429) );
  NAND2X0 U400 ( .IN1(n457), .IN2(n5), .QN(n430) );
  NAND3X0 U401 ( .IN1(n428), .IN2(n429), .IN3(n430), .QN(n4) );
  NAND2X0 U402 ( .IN1(n25), .IN2(n153), .QN(n431) );
  NAND2X0 U403 ( .IN1(n25), .IN2(n4), .QN(n432) );
  NAND2X0 U404 ( .IN1(n153), .IN2(n4), .QN(n433) );
  NAND2X0 U405 ( .IN1(n118), .IN2(n123), .QN(n434) );
  NAND2X0 U406 ( .IN1(n118), .IN2(n19), .QN(n435) );
  NAND2X0 U407 ( .IN1(n123), .IN2(n19), .QN(n436) );
  NAND3X0 U408 ( .IN1(n434), .IN2(n435), .IN3(n436), .QN(n18) );
  NAND2X0 U409 ( .IN1(n112), .IN2(n117), .QN(n437) );
  NAND2X0 U410 ( .IN1(n112), .IN2(n18), .QN(n438) );
  NAND2X0 U411 ( .IN1(n117), .IN2(n18), .QN(n439) );
  NAND3X0 U412 ( .IN1(n437), .IN2(n438), .IN3(n439), .QN(n17) );
  NAND2X0 U413 ( .IN1(n124), .IN2(n20), .QN(n440) );
  NAND2X0 U414 ( .IN1(n127), .IN2(n20), .QN(n441) );
  NAND2X0 U415 ( .IN1(n127), .IN2(n124), .QN(n442) );
  NAND3X0 U416 ( .IN1(n440), .IN2(n442), .IN3(n441), .QN(n19) );
  DELLN1X2 U417 ( .INP(a[11]), .Z(n456) );
  INVX0 U418 ( .INP(n445), .ZN(n444) );
  INVX0 U419 ( .INP(b[0]), .ZN(n445) );
  INVX0 U420 ( .INP(n447), .ZN(n446) );
  INVX0 U421 ( .INP(a[0]), .ZN(n447) );
  DELLN1X2 U422 ( .INP(a[3]), .Z(n448) );
  DELLN1X2 U423 ( .INP(a[5]), .Z(n450) );
  DELLN1X2 U424 ( .INP(a[7]), .Z(n452) );
  DELLN1X2 U425 ( .INP(a[9]), .Z(n454) );
  NOR2X0 U426 ( .IN1(n447), .IN2(n445), .QN(product[0]) );
  XNOR2X1 U427 ( .IN1(n467), .IN2(n468), .Q(n84) );
  NAND2X0 U428 ( .IN1(n468), .IN2(n467), .QN(n83) );
  AOI22X1 U429 ( .IN1(n469), .IN2(n466), .IN3(n470), .IN4(n471), .QN(n467) );
  OA21X1 U430 ( .IN1(n472), .IN2(n446), .IN3(n473), .Q(n468) );
  AO22X1 U431 ( .IN1(n474), .IN2(n466), .IN3(n470), .IN4(n469), .Q(n73) );
  AO22X1 U432 ( .IN1(n475), .IN2(n464), .IN3(n476), .IN4(n477), .Q(n55) );
  AO22X1 U433 ( .IN1(n478), .IN2(n462), .IN3(n479), .IN4(n480), .Q(n41) );
  AO22X1 U434 ( .IN1(n481), .IN2(n460), .IN3(n482), .IN4(n483), .Q(n31) );
  AO22X1 U435 ( .IN1(n484), .IN2(n458), .IN3(n485), .IN4(n486), .Q(n25) );
  AO22X1 U436 ( .IN1(n446), .IN2(n487), .IN3(n472), .IN4(n445), .Q(n224) );
  AO22X1 U437 ( .IN1(n446), .IN2(n488), .IN3(n472), .IN4(n487), .Q(n223) );
  AO22X1 U438 ( .IN1(n446), .IN2(n489), .IN3(n472), .IN4(n488), .Q(n222) );
  XOR2X1 U439 ( .IN1(n414), .IN2(n443), .Q(n488) );
  AO22X1 U440 ( .IN1(n446), .IN2(n490), .IN3(n472), .IN4(n489), .Q(n221) );
  AO22X1 U441 ( .IN1(n446), .IN2(n491), .IN3(n472), .IN4(n490), .Q(n220) );
  XOR2X1 U442 ( .IN1(b[4]), .IN2(n443), .Q(n490) );
  AO22X1 U443 ( .IN1(n446), .IN2(n492), .IN3(n472), .IN4(n491), .Q(n219) );
  AO22X1 U444 ( .IN1(n446), .IN2(n493), .IN3(n472), .IN4(n492), .Q(n218) );
  AO22X1 U445 ( .IN1(n446), .IN2(n494), .IN3(n472), .IN4(n493), .Q(n217) );
  XOR2X1 U446 ( .IN1(b[7]), .IN2(n443), .Q(n493) );
  AO22X1 U447 ( .IN1(n446), .IN2(n495), .IN3(n472), .IN4(n494), .Q(n216) );
  AO22X1 U448 ( .IN1(n446), .IN2(n496), .IN3(n472), .IN4(n495), .Q(n215) );
  XOR2X1 U449 ( .IN1(b[9]), .IN2(n443), .Q(n495) );
  AO22X1 U450 ( .IN1(n446), .IN2(n473), .IN3(n472), .IN4(n496), .Q(n214) );
  XOR2X1 U451 ( .IN1(b[11]), .IN2(n443), .Q(n473) );
  NOR2X0 U452 ( .IN1(n497), .IN2(n445), .QN(n212) );
  AO22X1 U453 ( .IN1(n498), .IN2(n466), .IN3(n470), .IN4(n499), .Q(n211) );
  XOR2X1 U454 ( .IN1(n444), .IN2(n448), .Q(n499) );
  AO22X1 U455 ( .IN1(n500), .IN2(n466), .IN3(n470), .IN4(n498), .Q(n210) );
  AO22X1 U456 ( .IN1(n501), .IN2(n466), .IN3(n470), .IN4(n500), .Q(n209) );
  XOR2X1 U457 ( .IN1(n414), .IN2(n448), .Q(n500) );
  AO22X1 U458 ( .IN1(n502), .IN2(n466), .IN3(n470), .IN4(n501), .Q(n208) );
  AO22X1 U459 ( .IN1(n503), .IN2(n466), .IN3(n470), .IN4(n502), .Q(n207) );
  XOR2X1 U460 ( .IN1(b[4]), .IN2(n448), .Q(n502) );
  AO22X1 U461 ( .IN1(n504), .IN2(n466), .IN3(n470), .IN4(n503), .Q(n206) );
  AO22X1 U462 ( .IN1(n505), .IN2(n466), .IN3(n470), .IN4(n504), .Q(n205) );
  AO22X1 U463 ( .IN1(n506), .IN2(n466), .IN3(n470), .IN4(n505), .Q(n204) );
  XOR2X1 U464 ( .IN1(b[7]), .IN2(n448), .Q(n505) );
  AO22X1 U465 ( .IN1(n471), .IN2(n466), .IN3(n470), .IN4(n506), .Q(n203) );
  XOR2X1 U466 ( .IN1(b[9]), .IN2(n448), .Q(n471) );
  OAI21X1 U467 ( .IN1(n466), .IN2(n470), .IN3(n474), .QN(n201) );
  XOR2X1 U468 ( .IN1(b[11]), .IN2(n448), .Q(n474) );
  NOR2X0 U469 ( .IN1(n507), .IN2(n445), .QN(n200) );
  AO22X1 U470 ( .IN1(n508), .IN2(n464), .IN3(n476), .IN4(n509), .Q(n199) );
  XOR2X1 U471 ( .IN1(n444), .IN2(n450), .Q(n509) );
  AO22X1 U472 ( .IN1(n510), .IN2(n464), .IN3(n476), .IN4(n508), .Q(n198) );
  AO22X1 U473 ( .IN1(n511), .IN2(n464), .IN3(n476), .IN4(n510), .Q(n197) );
  XOR2X1 U474 ( .IN1(n414), .IN2(n450), .Q(n510) );
  AO22X1 U475 ( .IN1(n512), .IN2(n464), .IN3(n476), .IN4(n511), .Q(n196) );
  AO22X1 U476 ( .IN1(n513), .IN2(n464), .IN3(n476), .IN4(n512), .Q(n195) );
  XOR2X1 U477 ( .IN1(b[4]), .IN2(n450), .Q(n512) );
  AO22X1 U478 ( .IN1(n514), .IN2(n464), .IN3(n476), .IN4(n513), .Q(n194) );
  AO22X1 U479 ( .IN1(n515), .IN2(n464), .IN3(n476), .IN4(n514), .Q(n193) );
  AO22X1 U480 ( .IN1(n516), .IN2(n464), .IN3(n476), .IN4(n515), .Q(n192) );
  XOR2X1 U481 ( .IN1(b[7]), .IN2(n450), .Q(n515) );
  AO22X1 U482 ( .IN1(n517), .IN2(n464), .IN3(n476), .IN4(n516), .Q(n191) );
  AO22X1 U483 ( .IN1(n477), .IN2(n464), .IN3(n476), .IN4(n517), .Q(n190) );
  XOR2X1 U484 ( .IN1(b[9]), .IN2(n450), .Q(n517) );
  OAI21X1 U485 ( .IN1(n464), .IN2(n476), .IN3(n475), .QN(n189) );
  XOR2X1 U486 ( .IN1(b[11]), .IN2(n450), .Q(n475) );
  NOR2X0 U487 ( .IN1(n518), .IN2(n445), .QN(n188) );
  AO22X1 U488 ( .IN1(n519), .IN2(n462), .IN3(n479), .IN4(n520), .Q(n187) );
  XOR2X1 U489 ( .IN1(n444), .IN2(n452), .Q(n520) );
  AO22X1 U490 ( .IN1(n521), .IN2(n462), .IN3(n479), .IN4(n519), .Q(n186) );
  AO22X1 U491 ( .IN1(n522), .IN2(n462), .IN3(n479), .IN4(n521), .Q(n185) );
  XOR2X1 U492 ( .IN1(n414), .IN2(n452), .Q(n521) );
  AO22X1 U493 ( .IN1(n523), .IN2(n462), .IN3(n479), .IN4(n522), .Q(n184) );
  AO22X1 U494 ( .IN1(n524), .IN2(n462), .IN3(n479), .IN4(n523), .Q(n183) );
  XOR2X1 U495 ( .IN1(b[4]), .IN2(n452), .Q(n523) );
  AO22X1 U496 ( .IN1(n525), .IN2(n462), .IN3(n479), .IN4(n524), .Q(n182) );
  AO22X1 U497 ( .IN1(n526), .IN2(n462), .IN3(n479), .IN4(n525), .Q(n181) );
  AO22X1 U498 ( .IN1(n527), .IN2(n462), .IN3(n479), .IN4(n526), .Q(n180) );
  XOR2X1 U499 ( .IN1(b[7]), .IN2(n452), .Q(n526) );
  AO22X1 U500 ( .IN1(n528), .IN2(n462), .IN3(n479), .IN4(n527), .Q(n179) );
  AO22X1 U501 ( .IN1(n480), .IN2(n462), .IN3(n479), .IN4(n528), .Q(n178) );
  XOR2X1 U502 ( .IN1(b[9]), .IN2(n452), .Q(n528) );
  OAI21X1 U503 ( .IN1(n462), .IN2(n479), .IN3(n478), .QN(n177) );
  XOR2X1 U504 ( .IN1(b[11]), .IN2(n452), .Q(n478) );
  NOR2X0 U505 ( .IN1(n529), .IN2(n445), .QN(n176) );
  AO22X1 U506 ( .IN1(n530), .IN2(n460), .IN3(n482), .IN4(n531), .Q(n175) );
  XOR2X1 U507 ( .IN1(n444), .IN2(n454), .Q(n531) );
  AO22X1 U508 ( .IN1(n532), .IN2(n460), .IN3(n482), .IN4(n530), .Q(n174) );
  AO22X1 U509 ( .IN1(n533), .IN2(n460), .IN3(n482), .IN4(n532), .Q(n173) );
  XOR2X1 U510 ( .IN1(n414), .IN2(n454), .Q(n532) );
  AO22X1 U511 ( .IN1(n534), .IN2(n460), .IN3(n482), .IN4(n533), .Q(n172) );
  AO22X1 U512 ( .IN1(n535), .IN2(n460), .IN3(n482), .IN4(n534), .Q(n171) );
  XOR2X1 U513 ( .IN1(b[4]), .IN2(n454), .Q(n534) );
  AO22X1 U514 ( .IN1(n536), .IN2(n460), .IN3(n482), .IN4(n535), .Q(n170) );
  AO22X1 U515 ( .IN1(n537), .IN2(n460), .IN3(n482), .IN4(n536), .Q(n169) );
  AO22X1 U516 ( .IN1(n538), .IN2(n460), .IN3(n482), .IN4(n537), .Q(n168) );
  XOR2X1 U517 ( .IN1(b[7]), .IN2(n454), .Q(n537) );
  AO22X1 U518 ( .IN1(n539), .IN2(n460), .IN3(n482), .IN4(n538), .Q(n167) );
  AO22X1 U519 ( .IN1(n483), .IN2(n460), .IN3(n482), .IN4(n539), .Q(n166) );
  XOR2X1 U520 ( .IN1(b[9]), .IN2(n454), .Q(n539) );
  OAI21X1 U521 ( .IN1(n460), .IN2(n482), .IN3(n481), .QN(n165) );
  XOR2X1 U522 ( .IN1(b[11]), .IN2(n454), .Q(n481) );
  NOR2X0 U523 ( .IN1(n540), .IN2(n445), .QN(n164) );
  AO22X1 U524 ( .IN1(n541), .IN2(n458), .IN3(n485), .IN4(n542), .Q(n163) );
  XOR2X1 U525 ( .IN1(n444), .IN2(n456), .Q(n542) );
  AO22X1 U526 ( .IN1(n543), .IN2(n458), .IN3(n485), .IN4(n541), .Q(n162) );
  AO22X1 U527 ( .IN1(n544), .IN2(n458), .IN3(n485), .IN4(n543), .Q(n161) );
  XOR2X1 U528 ( .IN1(n414), .IN2(n456), .Q(n543) );
  AO22X1 U529 ( .IN1(n545), .IN2(n458), .IN3(n485), .IN4(n544), .Q(n160) );
  AO22X1 U530 ( .IN1(n546), .IN2(n458), .IN3(n485), .IN4(n545), .Q(n159) );
  XOR2X1 U531 ( .IN1(b[4]), .IN2(n456), .Q(n545) );
  AO22X1 U532 ( .IN1(n547), .IN2(n458), .IN3(n485), .IN4(n546), .Q(n158) );
  AO22X1 U533 ( .IN1(n548), .IN2(n458), .IN3(n485), .IN4(n547), .Q(n157) );
  AO22X1 U534 ( .IN1(n549), .IN2(n458), .IN3(n485), .IN4(n548), .Q(n156) );
  XOR2X1 U535 ( .IN1(b[7]), .IN2(n456), .Q(n548) );
  AO22X1 U536 ( .IN1(n550), .IN2(n458), .IN3(n485), .IN4(n549), .Q(n155) );
  AO22X1 U537 ( .IN1(n486), .IN2(n458), .IN3(n485), .IN4(n550), .Q(n154) );
  XOR2X1 U538 ( .IN1(b[9]), .IN2(n456), .Q(n550) );
  OAI21X1 U539 ( .IN1(n458), .IN2(n485), .IN3(n484), .QN(n153) );
  XOR2X1 U540 ( .IN1(b[11]), .IN2(n456), .Q(n484) );
  AO21X1 U541 ( .IN1(n443), .IN2(n445), .IN3(n472), .Q(n152) );
  AO22X1 U542 ( .IN1(n551), .IN2(n449), .IN3(n470), .IN4(n449), .Q(n151) );
  XOR2X1 U543 ( .IN1(n448), .IN2(a[2]), .Q(n552) );
  NOR2X0 U544 ( .IN1(n444), .IN2(n497), .QN(n551) );
  XNOR2X1 U545 ( .IN1(a[2]), .IN2(n443), .Q(n497) );
  AO22X1 U546 ( .IN1(n553), .IN2(n451), .IN3(n476), .IN4(n451), .Q(n150) );
  XOR2X1 U547 ( .IN1(n450), .IN2(a[4]), .Q(n554) );
  NOR2X0 U548 ( .IN1(n444), .IN2(n507), .QN(n553) );
  XNOR2X1 U549 ( .IN1(a[4]), .IN2(n448), .Q(n507) );
  AO22X1 U550 ( .IN1(n555), .IN2(n453), .IN3(n479), .IN4(n453), .Q(n149) );
  XOR2X1 U551 ( .IN1(n452), .IN2(a[6]), .Q(n556) );
  NOR2X0 U552 ( .IN1(n444), .IN2(n518), .QN(n555) );
  XNOR2X1 U553 ( .IN1(a[6]), .IN2(n450), .Q(n518) );
  AO22X1 U554 ( .IN1(n557), .IN2(n455), .IN3(n482), .IN4(n455), .Q(n148) );
  XOR2X1 U555 ( .IN1(n454), .IN2(a[8]), .Q(n558) );
  NOR2X0 U556 ( .IN1(n444), .IN2(n529), .QN(n557) );
  XNOR2X1 U557 ( .IN1(a[8]), .IN2(n452), .Q(n529) );
  AO22X1 U558 ( .IN1(n559), .IN2(n456), .IN3(n485), .IN4(n456), .Q(n147) );
  XOR2X1 U559 ( .IN1(n456), .IN2(a[10]), .Q(n560) );
  NOR2X0 U560 ( .IN1(n444), .IN2(n540), .QN(n559) );
  XNOR2X1 U561 ( .IN1(a[10]), .IN2(n454), .Q(n540) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_15 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;
  wire   n1, n2;
  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_15_DW_mult_tc_0 mult_30 ( .a(in_a), .b({
        in_b[11:5], n2, in_b[3:0]}), .product(pre_out) );
  INVX0 U3 ( .INP(in_b[4]), .ZN(n1) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_14_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n461), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n23), .B(n151), .CI(n134), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n463), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n465), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n467), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n469), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  XOR3X1 U311 ( .IN1(n49), .IN2(n44), .IN3(n410), .Q(product[16]) );
  FADDX1 U312 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  INVX0 U313 ( .INP(b[6]), .ZN(n408) );
  INVX0 U314 ( .INP(n408), .ZN(n409) );
  DELLN2X2 U315 ( .INP(n10), .Z(n410) );
  INVX0 U316 ( .INP(b[5]), .ZN(n411) );
  INVX0 U317 ( .INP(n411), .ZN(n412) );
  DELLN2X2 U318 ( .INP(n18), .Z(n413) );
  INVX0 U319 ( .INP(b[1]), .ZN(n414) );
  INVX0 U320 ( .INP(n414), .ZN(n415) );
  DELLN2X2 U321 ( .INP(n9), .Z(n416) );
  INVX0 U322 ( .INP(b[4]), .ZN(n417) );
  INVX0 U323 ( .INP(n417), .ZN(n418) );
  INVX0 U324 ( .INP(b[2]), .ZN(n419) );
  INVX0 U325 ( .INP(n419), .ZN(n420) );
  XOR2X2 U326 ( .IN1(b[11]), .IN2(n459), .Q(n488) );
  XOR2X2 U327 ( .IN1(b[11]), .IN2(n457), .Q(n485) );
  XOR2X2 U328 ( .IN1(b[11]), .IN2(n455), .Q(n482) );
  XOR2X2 U329 ( .IN1(b[11]), .IN2(n453), .Q(n479) );
  XOR2X2 U330 ( .IN1(b[11]), .IN2(n451), .Q(n478) );
  XOR2X2 U331 ( .IN1(b[11]), .IN2(n446), .Q(n477) );
  XOR2X2 U332 ( .IN1(b[10]), .IN2(n459), .Q(n490) );
  XOR2X2 U333 ( .IN1(b[10]), .IN2(n457), .Q(n487) );
  XOR2X2 U334 ( .IN1(b[10]), .IN2(n455), .Q(n484) );
  XOR2X2 U335 ( .IN1(b[10]), .IN2(n453), .Q(n481) );
  XOR2X2 U336 ( .IN1(b[10]), .IN2(n451), .Q(n473) );
  XOR2X2 U337 ( .IN1(b[10]), .IN2(n446), .Q(n500) );
  XOR3X2 U338 ( .IN1(n65), .IN2(n58), .IN3(n12), .Q(product[14]) );
  XOR2X2 U339 ( .IN1(n420), .IN2(n459), .Q(n547) );
  XOR2X2 U340 ( .IN1(n420), .IN2(n457), .Q(n536) );
  XOR2X2 U341 ( .IN1(n420), .IN2(n455), .Q(n525) );
  XOR2X2 U342 ( .IN1(n420), .IN2(n453), .Q(n514) );
  XOR2X2 U343 ( .IN1(n420), .IN2(n451), .Q(n504) );
  XOR2X2 U344 ( .IN1(n420), .IN2(n446), .Q(n492) );
  XOR2X2 U345 ( .IN1(b[9]), .IN2(n459), .Q(n554) );
  XOR2X2 U346 ( .IN1(b[9]), .IN2(n457), .Q(n543) );
  XOR2X2 U347 ( .IN1(b[9]), .IN2(n455), .Q(n532) );
  XOR2X2 U348 ( .IN1(b[9]), .IN2(n453), .Q(n521) );
  XOR2X2 U349 ( .IN1(b[9]), .IN2(n451), .Q(n475) );
  XOR2X2 U350 ( .IN1(b[9]), .IN2(n446), .Q(n499) );
  XOR3X2 U351 ( .IN1(n118), .IN2(n123), .IN3(n19), .Q(product[7]) );
  NAND2X0 U352 ( .IN1(n118), .IN2(n123), .QN(n421) );
  NAND2X0 U353 ( .IN1(n118), .IN2(n19), .QN(n422) );
  NAND2X0 U354 ( .IN1(n123), .IN2(n19), .QN(n423) );
  NAND3X0 U355 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n18) );
  XOR2X1 U356 ( .IN1(n112), .IN2(n117), .Q(n424) );
  XOR2X1 U357 ( .IN1(n424), .IN2(n413), .Q(product[8]) );
  NAND2X0 U358 ( .IN1(n112), .IN2(n117), .QN(n425) );
  NAND2X0 U359 ( .IN1(n112), .IN2(n18), .QN(n426) );
  NAND2X0 U360 ( .IN1(n117), .IN2(n18), .QN(n427) );
  NAND3X0 U361 ( .IN1(n425), .IN2(n426), .IN3(n427), .QN(n17) );
  XOR2X2 U362 ( .IN1(b[8]), .IN2(n459), .Q(n553) );
  XOR2X2 U363 ( .IN1(b[8]), .IN2(n457), .Q(n542) );
  XOR2X2 U364 ( .IN1(b[8]), .IN2(n455), .Q(n531) );
  XOR2X2 U365 ( .IN1(b[8]), .IN2(n453), .Q(n520) );
  XOR2X2 U366 ( .IN1(b[8]), .IN2(n451), .Q(n510) );
  XOR2X2 U367 ( .IN1(b[8]), .IN2(n446), .Q(n498) );
  XOR2X2 U368 ( .IN1(b[7]), .IN2(n459), .Q(n552) );
  XOR2X2 U369 ( .IN1(b[7]), .IN2(n457), .Q(n541) );
  XOR2X2 U370 ( .IN1(b[7]), .IN2(n455), .Q(n530) );
  XOR2X2 U371 ( .IN1(b[7]), .IN2(n453), .Q(n519) );
  XOR2X2 U372 ( .IN1(b[7]), .IN2(n451), .Q(n509) );
  XOR2X2 U373 ( .IN1(b[7]), .IN2(n446), .Q(n497) );
  XOR2X2 U374 ( .IN1(n409), .IN2(n459), .Q(n551) );
  XOR2X2 U375 ( .IN1(n409), .IN2(n457), .Q(n540) );
  XOR2X2 U376 ( .IN1(n409), .IN2(n455), .Q(n529) );
  XOR2X2 U377 ( .IN1(n409), .IN2(n453), .Q(n518) );
  XOR2X2 U378 ( .IN1(n409), .IN2(n451), .Q(n508) );
  XOR2X2 U379 ( .IN1(n409), .IN2(n446), .Q(n496) );
  XOR2X2 U380 ( .IN1(b[3]), .IN2(n459), .Q(n548) );
  XOR2X2 U381 ( .IN1(b[3]), .IN2(n457), .Q(n537) );
  XOR2X2 U382 ( .IN1(b[3]), .IN2(n455), .Q(n526) );
  XOR2X2 U383 ( .IN1(b[3]), .IN2(n453), .Q(n515) );
  XOR2X2 U384 ( .IN1(b[3]), .IN2(n451), .Q(n505) );
  XOR2X2 U385 ( .IN1(b[3]), .IN2(n446), .Q(n493) );
  XOR2X2 U386 ( .IN1(n415), .IN2(n459), .Q(n545) );
  XOR2X2 U387 ( .IN1(n415), .IN2(n457), .Q(n534) );
  XOR2X2 U388 ( .IN1(n415), .IN2(n455), .Q(n523) );
  XOR2X2 U389 ( .IN1(n415), .IN2(n453), .Q(n512) );
  XOR2X2 U390 ( .IN1(n415), .IN2(n451), .Q(n502) );
  XOR2X2 U391 ( .IN1(n415), .IN2(n446), .Q(n491) );
  XOR2X2 U392 ( .IN1(n412), .IN2(n459), .Q(n550) );
  XOR2X2 U393 ( .IN1(n412), .IN2(n457), .Q(n539) );
  XOR2X2 U394 ( .IN1(n412), .IN2(n455), .Q(n528) );
  XOR2X2 U395 ( .IN1(n412), .IN2(n453), .Q(n517) );
  XOR2X2 U396 ( .IN1(n412), .IN2(n451), .Q(n507) );
  XOR2X2 U397 ( .IN1(n418), .IN2(n459), .Q(n549) );
  XOR2X2 U398 ( .IN1(n418), .IN2(n457), .Q(n538) );
  XOR2X2 U399 ( .IN1(n418), .IN2(n455), .Q(n527) );
  XOR2X2 U400 ( .IN1(n418), .IN2(n453), .Q(n516) );
  XOR2X2 U401 ( .IN1(n418), .IN2(n451), .Q(n506) );
  XOR2X2 U402 ( .IN1(n418), .IN2(n446), .Q(n494) );
  NAND2X1 U403 ( .IN1(n49), .IN2(n44), .QN(n428) );
  NAND2X0 U404 ( .IN1(n49), .IN2(n10), .QN(n429) );
  NAND2X0 U405 ( .IN1(n44), .IN2(n10), .QN(n430) );
  NAND3X0 U406 ( .IN1(n428), .IN2(n429), .IN3(n430), .QN(n9) );
  XOR2X1 U407 ( .IN1(n43), .IN2(n38), .Q(n431) );
  XOR2X1 U408 ( .IN1(n431), .IN2(n416), .Q(product[17]) );
  NAND2X1 U409 ( .IN1(n43), .IN2(n38), .QN(n432) );
  NAND2X0 U410 ( .IN1(n43), .IN2(n9), .QN(n433) );
  NAND2X0 U411 ( .IN1(n38), .IN2(n9), .QN(n434) );
  NAND3X0 U412 ( .IN1(n432), .IN2(n433), .IN3(n434), .QN(n8) );
  FADDX1 U413 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U414 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U415 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  XNOR2X1 U416 ( .IN1(n435), .IN2(n11), .Q(product[15]) );
  XNOR2X1 U417 ( .IN1(n57), .IN2(n50), .Q(n435) );
  XNOR2X1 U418 ( .IN1(n436), .IN2(n13), .Q(product[13]) );
  XNOR2X1 U419 ( .IN1(n66), .IN2(n75), .Q(n436) );
  INVX0 U420 ( .INP(n25), .ZN(n461) );
  INVX0 U421 ( .INP(n3), .ZN(product[23]) );
  INVX0 U422 ( .INP(n55), .ZN(n467) );
  FADDX1 U423 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  INVX0 U424 ( .INP(n73), .ZN(n469) );
  FADDX1 U425 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U426 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  INVX0 U427 ( .INP(n31), .ZN(n463) );
  INVX0 U428 ( .INP(n41), .ZN(n465) );
  DELLN1X2 U429 ( .INP(a[1]), .Z(n446) );
  AND2X1 U430 ( .IN1(n446), .IN2(n450), .Q(n476) );
  INVX0 U431 ( .INP(n501), .ZN(n470) );
  INVX0 U432 ( .INP(n522), .ZN(n466) );
  INVX0 U433 ( .INP(n511), .ZN(n468) );
  INVX0 U434 ( .INP(n533), .ZN(n464) );
  INVX0 U435 ( .INP(n544), .ZN(n462) );
  NBUFFX2 U436 ( .INP(a[3]), .Z(n452) );
  FADDX1 U437 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  NBUFFX2 U438 ( .INP(a[5]), .Z(n454) );
  NBUFFX2 U439 ( .INP(a[7]), .Z(n456) );
  NBUFFX2 U440 ( .INP(a[9]), .Z(n458) );
  XOR2X2 U441 ( .IN1(n412), .IN2(n446), .Q(n495) );
  NAND2X0 U442 ( .IN1(n65), .IN2(n58), .QN(n437) );
  NAND2X0 U443 ( .IN1(n65), .IN2(n12), .QN(n438) );
  NAND2X0 U444 ( .IN1(n58), .IN2(n12), .QN(n439) );
  NAND3X0 U445 ( .IN1(n439), .IN2(n438), .IN3(n437), .QN(n11) );
  NAND2X0 U446 ( .IN1(n57), .IN2(n50), .QN(n440) );
  NAND2X0 U447 ( .IN1(n57), .IN2(n11), .QN(n441) );
  NAND2X0 U448 ( .IN1(n50), .IN2(n11), .QN(n442) );
  NAND3X0 U449 ( .IN1(n442), .IN2(n441), .IN3(n440), .QN(n10) );
  NAND2X0 U450 ( .IN1(n75), .IN2(n13), .QN(n443) );
  NAND2X0 U451 ( .IN1(n66), .IN2(n13), .QN(n444) );
  NAND2X0 U452 ( .IN1(n66), .IN2(n75), .QN(n445) );
  NAND3X0 U453 ( .IN1(n443), .IN2(n445), .IN3(n444), .QN(n12) );
  DELLN1X2 U454 ( .INP(a[11]), .Z(n459) );
  AND2X2 U455 ( .IN1(n501), .IN2(n556), .Q(n474) );
  AND2X2 U456 ( .IN1(n511), .IN2(n558), .Q(n480) );
  AND2X2 U457 ( .IN1(n522), .IN2(n560), .Q(n483) );
  AND2X2 U458 ( .IN1(n533), .IN2(n562), .Q(n486) );
  AND2X2 U459 ( .IN1(n544), .IN2(n564), .Q(n489) );
  INVX0 U460 ( .INP(n448), .ZN(n447) );
  INVX0 U461 ( .INP(b[0]), .ZN(n448) );
  INVX0 U462 ( .INP(n450), .ZN(n449) );
  INVX0 U463 ( .INP(a[0]), .ZN(n450) );
  DELLN1X2 U464 ( .INP(a[3]), .Z(n451) );
  DELLN1X2 U465 ( .INP(a[5]), .Z(n453) );
  DELLN1X2 U466 ( .INP(a[7]), .Z(n455) );
  DELLN1X2 U467 ( .INP(a[9]), .Z(n457) );
  NOR2X0 U468 ( .IN1(n450), .IN2(n448), .QN(product[0]) );
  XNOR2X1 U469 ( .IN1(n471), .IN2(n472), .Q(n84) );
  NAND2X0 U470 ( .IN1(n472), .IN2(n471), .QN(n83) );
  AOI22X1 U471 ( .IN1(n473), .IN2(n470), .IN3(n474), .IN4(n475), .QN(n471) );
  OA21X1 U472 ( .IN1(n476), .IN2(n449), .IN3(n477), .Q(n472) );
  AO22X1 U473 ( .IN1(n478), .IN2(n470), .IN3(n474), .IN4(n473), .Q(n73) );
  AO22X1 U474 ( .IN1(n479), .IN2(n468), .IN3(n480), .IN4(n481), .Q(n55) );
  AO22X1 U475 ( .IN1(n482), .IN2(n466), .IN3(n483), .IN4(n484), .Q(n41) );
  AO22X1 U476 ( .IN1(n485), .IN2(n464), .IN3(n486), .IN4(n487), .Q(n31) );
  AO22X1 U477 ( .IN1(n488), .IN2(n462), .IN3(n489), .IN4(n490), .Q(n25) );
  AO22X1 U478 ( .IN1(n449), .IN2(n491), .IN3(n476), .IN4(n448), .Q(n224) );
  AO22X1 U479 ( .IN1(n449), .IN2(n492), .IN3(n476), .IN4(n491), .Q(n223) );
  AO22X1 U480 ( .IN1(n449), .IN2(n493), .IN3(n476), .IN4(n492), .Q(n222) );
  AO22X1 U481 ( .IN1(n449), .IN2(n494), .IN3(n476), .IN4(n493), .Q(n221) );
  AO22X1 U482 ( .IN1(n449), .IN2(n495), .IN3(n476), .IN4(n494), .Q(n220) );
  AO22X1 U483 ( .IN1(n449), .IN2(n496), .IN3(n476), .IN4(n495), .Q(n219) );
  AO22X1 U484 ( .IN1(n449), .IN2(n497), .IN3(n476), .IN4(n496), .Q(n218) );
  AO22X1 U485 ( .IN1(n449), .IN2(n498), .IN3(n476), .IN4(n497), .Q(n217) );
  AO22X1 U486 ( .IN1(n449), .IN2(n499), .IN3(n476), .IN4(n498), .Q(n216) );
  AO22X1 U487 ( .IN1(n449), .IN2(n500), .IN3(n476), .IN4(n499), .Q(n215) );
  AO22X1 U488 ( .IN1(n449), .IN2(n477), .IN3(n476), .IN4(n500), .Q(n214) );
  NOR2X0 U489 ( .IN1(n501), .IN2(n448), .QN(n212) );
  AO22X1 U490 ( .IN1(n502), .IN2(n470), .IN3(n474), .IN4(n503), .Q(n211) );
  XOR2X1 U491 ( .IN1(n447), .IN2(n451), .Q(n503) );
  AO22X1 U492 ( .IN1(n504), .IN2(n470), .IN3(n474), .IN4(n502), .Q(n210) );
  AO22X1 U493 ( .IN1(n505), .IN2(n470), .IN3(n474), .IN4(n504), .Q(n209) );
  AO22X1 U494 ( .IN1(n506), .IN2(n470), .IN3(n474), .IN4(n505), .Q(n208) );
  AO22X1 U495 ( .IN1(n507), .IN2(n470), .IN3(n474), .IN4(n506), .Q(n207) );
  AO22X1 U496 ( .IN1(n508), .IN2(n470), .IN3(n474), .IN4(n507), .Q(n206) );
  AO22X1 U497 ( .IN1(n509), .IN2(n470), .IN3(n474), .IN4(n508), .Q(n205) );
  AO22X1 U498 ( .IN1(n510), .IN2(n470), .IN3(n474), .IN4(n509), .Q(n204) );
  AO22X1 U499 ( .IN1(n475), .IN2(n470), .IN3(n474), .IN4(n510), .Q(n203) );
  OAI21X1 U500 ( .IN1(n470), .IN2(n474), .IN3(n478), .QN(n201) );
  NOR2X0 U501 ( .IN1(n511), .IN2(n448), .QN(n200) );
  AO22X1 U502 ( .IN1(n512), .IN2(n468), .IN3(n480), .IN4(n513), .Q(n199) );
  XOR2X1 U503 ( .IN1(n447), .IN2(n453), .Q(n513) );
  AO22X1 U504 ( .IN1(n514), .IN2(n468), .IN3(n480), .IN4(n512), .Q(n198) );
  AO22X1 U505 ( .IN1(n515), .IN2(n468), .IN3(n480), .IN4(n514), .Q(n197) );
  AO22X1 U506 ( .IN1(n516), .IN2(n468), .IN3(n480), .IN4(n515), .Q(n196) );
  AO22X1 U507 ( .IN1(n517), .IN2(n468), .IN3(n480), .IN4(n516), .Q(n195) );
  AO22X1 U508 ( .IN1(n518), .IN2(n468), .IN3(n480), .IN4(n517), .Q(n194) );
  AO22X1 U509 ( .IN1(n519), .IN2(n468), .IN3(n480), .IN4(n518), .Q(n193) );
  AO22X1 U510 ( .IN1(n520), .IN2(n468), .IN3(n480), .IN4(n519), .Q(n192) );
  AO22X1 U511 ( .IN1(n521), .IN2(n468), .IN3(n480), .IN4(n520), .Q(n191) );
  AO22X1 U512 ( .IN1(n481), .IN2(n468), .IN3(n480), .IN4(n521), .Q(n190) );
  OAI21X1 U513 ( .IN1(n468), .IN2(n480), .IN3(n479), .QN(n189) );
  NOR2X0 U514 ( .IN1(n522), .IN2(n448), .QN(n188) );
  AO22X1 U515 ( .IN1(n523), .IN2(n466), .IN3(n483), .IN4(n524), .Q(n187) );
  XOR2X1 U516 ( .IN1(n447), .IN2(n455), .Q(n524) );
  AO22X1 U517 ( .IN1(n525), .IN2(n466), .IN3(n483), .IN4(n523), .Q(n186) );
  AO22X1 U518 ( .IN1(n526), .IN2(n466), .IN3(n483), .IN4(n525), .Q(n185) );
  AO22X1 U519 ( .IN1(n527), .IN2(n466), .IN3(n483), .IN4(n526), .Q(n184) );
  AO22X1 U520 ( .IN1(n528), .IN2(n466), .IN3(n483), .IN4(n527), .Q(n183) );
  AO22X1 U521 ( .IN1(n529), .IN2(n466), .IN3(n483), .IN4(n528), .Q(n182) );
  AO22X1 U522 ( .IN1(n530), .IN2(n466), .IN3(n483), .IN4(n529), .Q(n181) );
  AO22X1 U523 ( .IN1(n531), .IN2(n466), .IN3(n483), .IN4(n530), .Q(n180) );
  AO22X1 U524 ( .IN1(n532), .IN2(n466), .IN3(n483), .IN4(n531), .Q(n179) );
  AO22X1 U525 ( .IN1(n484), .IN2(n466), .IN3(n483), .IN4(n532), .Q(n178) );
  OAI21X1 U526 ( .IN1(n466), .IN2(n483), .IN3(n482), .QN(n177) );
  NOR2X0 U527 ( .IN1(n533), .IN2(n448), .QN(n176) );
  AO22X1 U528 ( .IN1(n534), .IN2(n464), .IN3(n486), .IN4(n535), .Q(n175) );
  XOR2X1 U529 ( .IN1(n447), .IN2(n457), .Q(n535) );
  AO22X1 U530 ( .IN1(n536), .IN2(n464), .IN3(n486), .IN4(n534), .Q(n174) );
  AO22X1 U531 ( .IN1(n537), .IN2(n464), .IN3(n486), .IN4(n536), .Q(n173) );
  AO22X1 U532 ( .IN1(n538), .IN2(n464), .IN3(n486), .IN4(n537), .Q(n172) );
  AO22X1 U533 ( .IN1(n539), .IN2(n464), .IN3(n486), .IN4(n538), .Q(n171) );
  AO22X1 U534 ( .IN1(n540), .IN2(n464), .IN3(n486), .IN4(n539), .Q(n170) );
  AO22X1 U535 ( .IN1(n541), .IN2(n464), .IN3(n486), .IN4(n540), .Q(n169) );
  AO22X1 U536 ( .IN1(n542), .IN2(n464), .IN3(n486), .IN4(n541), .Q(n168) );
  AO22X1 U537 ( .IN1(n543), .IN2(n464), .IN3(n486), .IN4(n542), .Q(n167) );
  AO22X1 U538 ( .IN1(n487), .IN2(n464), .IN3(n486), .IN4(n543), .Q(n166) );
  OAI21X1 U539 ( .IN1(n464), .IN2(n486), .IN3(n485), .QN(n165) );
  NOR2X0 U540 ( .IN1(n544), .IN2(n448), .QN(n164) );
  AO22X1 U541 ( .IN1(n545), .IN2(n462), .IN3(n489), .IN4(n546), .Q(n163) );
  XOR2X1 U542 ( .IN1(n447), .IN2(n459), .Q(n546) );
  AO22X1 U543 ( .IN1(n547), .IN2(n462), .IN3(n489), .IN4(n545), .Q(n162) );
  AO22X1 U544 ( .IN1(n548), .IN2(n462), .IN3(n489), .IN4(n547), .Q(n161) );
  AO22X1 U545 ( .IN1(n549), .IN2(n462), .IN3(n489), .IN4(n548), .Q(n160) );
  AO22X1 U546 ( .IN1(n550), .IN2(n462), .IN3(n489), .IN4(n549), .Q(n159) );
  AO22X1 U547 ( .IN1(n551), .IN2(n462), .IN3(n489), .IN4(n550), .Q(n158) );
  AO22X1 U548 ( .IN1(n552), .IN2(n462), .IN3(n489), .IN4(n551), .Q(n157) );
  AO22X1 U549 ( .IN1(n553), .IN2(n462), .IN3(n489), .IN4(n552), .Q(n156) );
  AO22X1 U550 ( .IN1(n554), .IN2(n462), .IN3(n489), .IN4(n553), .Q(n155) );
  AO22X1 U551 ( .IN1(n490), .IN2(n462), .IN3(n489), .IN4(n554), .Q(n154) );
  OAI21X1 U552 ( .IN1(n462), .IN2(n489), .IN3(n488), .QN(n153) );
  AO21X1 U553 ( .IN1(n446), .IN2(n448), .IN3(n476), .Q(n152) );
  AO22X1 U554 ( .IN1(n555), .IN2(n452), .IN3(n474), .IN4(n452), .Q(n151) );
  XOR2X1 U555 ( .IN1(n451), .IN2(a[2]), .Q(n556) );
  NOR2X0 U556 ( .IN1(n447), .IN2(n501), .QN(n555) );
  XNOR2X1 U557 ( .IN1(a[2]), .IN2(n446), .Q(n501) );
  AO22X1 U558 ( .IN1(n557), .IN2(n454), .IN3(n480), .IN4(n454), .Q(n150) );
  XOR2X1 U559 ( .IN1(n453), .IN2(a[4]), .Q(n558) );
  NOR2X0 U560 ( .IN1(n447), .IN2(n511), .QN(n557) );
  XNOR2X1 U561 ( .IN1(a[4]), .IN2(n451), .Q(n511) );
  AO22X1 U562 ( .IN1(n559), .IN2(n456), .IN3(n483), .IN4(n456), .Q(n149) );
  XOR2X1 U563 ( .IN1(n455), .IN2(a[6]), .Q(n560) );
  NOR2X0 U564 ( .IN1(n447), .IN2(n522), .QN(n559) );
  XNOR2X1 U565 ( .IN1(a[6]), .IN2(n453), .Q(n522) );
  AO22X1 U566 ( .IN1(n561), .IN2(n458), .IN3(n486), .IN4(n458), .Q(n148) );
  XOR2X1 U567 ( .IN1(n457), .IN2(a[8]), .Q(n562) );
  NOR2X0 U568 ( .IN1(n447), .IN2(n533), .QN(n561) );
  XNOR2X1 U569 ( .IN1(a[8]), .IN2(n455), .Q(n533) );
  AO22X1 U570 ( .IN1(n563), .IN2(n459), .IN3(n489), .IN4(n459), .Q(n147) );
  XOR2X1 U571 ( .IN1(n459), .IN2(a[10]), .Q(n564) );
  NOR2X0 U572 ( .IN1(n447), .IN2(n544), .QN(n563) );
  XNOR2X1 U573 ( .IN1(a[10]), .IN2(n457), .Q(n544) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_14 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_14_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_13_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555;

  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n454), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n456), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n458), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n460), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  AND3X1 U311 ( .IN1(n413), .IN2(n414), .IN3(n415), .Q(product[23]) );
  XOR2X2 U312 ( .IN1(b[11]), .IN2(n451), .Q(n479) );
  XOR2X2 U313 ( .IN1(b[11]), .IN2(n449), .Q(n476) );
  XOR2X2 U314 ( .IN1(b[11]), .IN2(n447), .Q(n473) );
  XOR2X2 U315 ( .IN1(b[11]), .IN2(n445), .Q(n470) );
  XOR2X2 U316 ( .IN1(b[11]), .IN2(n443), .Q(n469) );
  XOR2X2 U317 ( .IN1(b[11]), .IN2(a[1]), .Q(n468) );
  XOR2X2 U318 ( .IN1(b[10]), .IN2(n451), .Q(n481) );
  XOR2X2 U319 ( .IN1(b[10]), .IN2(n449), .Q(n478) );
  XOR2X2 U320 ( .IN1(b[10]), .IN2(n447), .Q(n475) );
  XOR2X2 U321 ( .IN1(b[10]), .IN2(n445), .Q(n472) );
  XOR2X2 U322 ( .IN1(b[10]), .IN2(n443), .Q(n464) );
  XOR2X2 U323 ( .IN1(b[10]), .IN2(a[1]), .Q(n491) );
  XOR2X2 U324 ( .IN1(b[2]), .IN2(n451), .Q(n538) );
  XOR2X2 U325 ( .IN1(b[2]), .IN2(n449), .Q(n527) );
  XOR2X2 U326 ( .IN1(b[2]), .IN2(n447), .Q(n516) );
  XOR2X2 U327 ( .IN1(b[2]), .IN2(n445), .Q(n505) );
  XOR2X2 U328 ( .IN1(b[2]), .IN2(n443), .Q(n495) );
  XOR2X2 U329 ( .IN1(b[2]), .IN2(a[1]), .Q(n483) );
  XOR2X2 U330 ( .IN1(b[9]), .IN2(n451), .Q(n545) );
  XOR2X2 U331 ( .IN1(b[9]), .IN2(n449), .Q(n534) );
  XOR2X2 U332 ( .IN1(b[9]), .IN2(n447), .Q(n523) );
  XOR2X2 U333 ( .IN1(b[9]), .IN2(n445), .Q(n512) );
  XOR2X2 U334 ( .IN1(b[9]), .IN2(n443), .Q(n466) );
  XOR2X2 U335 ( .IN1(b[9]), .IN2(a[1]), .Q(n490) );
  XOR2X2 U336 ( .IN1(b[8]), .IN2(n451), .Q(n544) );
  XOR2X2 U337 ( .IN1(b[8]), .IN2(n449), .Q(n533) );
  XOR2X2 U338 ( .IN1(b[8]), .IN2(n447), .Q(n522) );
  XOR2X2 U339 ( .IN1(b[8]), .IN2(n445), .Q(n511) );
  XOR2X2 U340 ( .IN1(b[8]), .IN2(n443), .Q(n501) );
  XOR2X2 U341 ( .IN1(b[8]), .IN2(a[1]), .Q(n489) );
  XOR2X2 U342 ( .IN1(b[7]), .IN2(n451), .Q(n543) );
  XOR2X2 U343 ( .IN1(b[7]), .IN2(n449), .Q(n532) );
  XOR2X2 U344 ( .IN1(b[7]), .IN2(n447), .Q(n521) );
  XOR2X2 U345 ( .IN1(b[7]), .IN2(n445), .Q(n510) );
  XOR2X2 U346 ( .IN1(b[7]), .IN2(n443), .Q(n500) );
  XOR2X2 U347 ( .IN1(b[7]), .IN2(a[1]), .Q(n488) );
  XOR2X2 U348 ( .IN1(b[6]), .IN2(n451), .Q(n542) );
  XOR2X2 U349 ( .IN1(b[6]), .IN2(n449), .Q(n531) );
  XOR2X2 U350 ( .IN1(b[6]), .IN2(n447), .Q(n520) );
  XOR2X2 U351 ( .IN1(b[6]), .IN2(n445), .Q(n509) );
  XOR2X2 U352 ( .IN1(b[6]), .IN2(n443), .Q(n499) );
  XOR2X2 U353 ( .IN1(b[6]), .IN2(a[1]), .Q(n487) );
  XOR2X2 U354 ( .IN1(b[3]), .IN2(n451), .Q(n539) );
  XOR2X2 U355 ( .IN1(b[3]), .IN2(n449), .Q(n528) );
  XOR2X2 U356 ( .IN1(b[3]), .IN2(n447), .Q(n517) );
  XOR2X2 U357 ( .IN1(b[3]), .IN2(n445), .Q(n506) );
  XOR2X2 U358 ( .IN1(b[3]), .IN2(n443), .Q(n496) );
  XOR2X2 U359 ( .IN1(b[3]), .IN2(a[1]), .Q(n484) );
  XOR3X2 U360 ( .IN1(n27), .IN2(n452), .IN3(n5), .Q(product[21]) );
  NAND2X0 U361 ( .IN1(n27), .IN2(n452), .QN(n409) );
  NAND2X0 U362 ( .IN1(n27), .IN2(n5), .QN(n410) );
  NAND2X0 U363 ( .IN1(n452), .IN2(n5), .QN(n411) );
  NAND3X0 U364 ( .IN1(n409), .IN2(n410), .IN3(n411), .QN(n4) );
  XOR2X2 U365 ( .IN1(n25), .IN2(n153), .Q(n412) );
  XOR2X1 U366 ( .IN1(n412), .IN2(n4), .Q(product[22]) );
  NAND2X0 U367 ( .IN1(n25), .IN2(n153), .QN(n413) );
  NAND2X0 U368 ( .IN1(n25), .IN2(n4), .QN(n414) );
  NAND2X0 U369 ( .IN1(n153), .IN2(n4), .QN(n415) );
  XOR3X2 U370 ( .IN1(n76), .IN2(n85), .IN3(n14), .Q(product[12]) );
  NAND2X1 U371 ( .IN1(n76), .IN2(n85), .QN(n416) );
  NAND2X0 U372 ( .IN1(n76), .IN2(n14), .QN(n417) );
  NAND2X0 U373 ( .IN1(n85), .IN2(n14), .QN(n418) );
  NAND3X0 U374 ( .IN1(n416), .IN2(n417), .IN3(n418), .QN(n13) );
  XOR2X1 U375 ( .IN1(n66), .IN2(n75), .Q(n419) );
  XOR2X1 U376 ( .IN1(n419), .IN2(n13), .Q(product[13]) );
  NAND2X0 U377 ( .IN1(n66), .IN2(n75), .QN(n420) );
  NAND2X0 U378 ( .IN1(n66), .IN2(n13), .QN(n421) );
  NAND2X0 U379 ( .IN1(n75), .IN2(n13), .QN(n422) );
  NAND3X0 U380 ( .IN1(n420), .IN2(n421), .IN3(n422), .QN(n12) );
  INVX0 U381 ( .INP(n15), .ZN(n423) );
  INVX0 U382 ( .INP(n423), .ZN(n424) );
  XOR2X2 U383 ( .IN1(b[1]), .IN2(n451), .Q(n536) );
  XOR2X2 U384 ( .IN1(b[1]), .IN2(n449), .Q(n525) );
  XOR2X2 U385 ( .IN1(b[1]), .IN2(n447), .Q(n514) );
  XOR2X2 U386 ( .IN1(b[1]), .IN2(n445), .Q(n503) );
  XOR2X2 U387 ( .IN1(b[1]), .IN2(n443), .Q(n493) );
  XOR2X2 U388 ( .IN1(b[1]), .IN2(a[1]), .Q(n482) );
  XOR2X2 U389 ( .IN1(b[5]), .IN2(n451), .Q(n541) );
  XOR2X2 U390 ( .IN1(b[5]), .IN2(n449), .Q(n530) );
  XOR2X2 U391 ( .IN1(b[5]), .IN2(n447), .Q(n519) );
  XOR2X2 U392 ( .IN1(b[5]), .IN2(n445), .Q(n508) );
  XOR2X2 U393 ( .IN1(b[5]), .IN2(n443), .Q(n498) );
  AO22X2 U394 ( .IN1(n441), .IN2(n487), .IN3(n467), .IN4(n486), .Q(n219) );
  AO22X1 U395 ( .IN1(n441), .IN2(n486), .IN3(n467), .IN4(n485), .Q(n220) );
  XOR2X2 U396 ( .IN1(b[5]), .IN2(a[1]), .Q(n486) );
  XOR2X2 U397 ( .IN1(b[4]), .IN2(n451), .Q(n540) );
  XOR2X2 U398 ( .IN1(b[4]), .IN2(n449), .Q(n529) );
  XOR2X2 U399 ( .IN1(b[4]), .IN2(n447), .Q(n518) );
  XOR2X2 U400 ( .IN1(b[4]), .IN2(n445), .Q(n507) );
  XOR2X2 U401 ( .IN1(b[4]), .IN2(n443), .Q(n497) );
  XOR2X2 U402 ( .IN1(b[4]), .IN2(a[1]), .Q(n485) );
  XOR3X1 U403 ( .IN1(n49), .IN2(n44), .IN3(n10), .Q(product[16]) );
  XNOR2X1 U404 ( .IN1(n9), .IN2(n425), .Q(product[17]) );
  XNOR2X1 U405 ( .IN1(n43), .IN2(n38), .Q(n425) );
  XOR3X1 U406 ( .IN1(n96), .IN2(n103), .IN3(n16), .Q(product[10]) );
  XNOR2X1 U407 ( .IN1(n426), .IN2(n424), .Q(product[11]) );
  XNOR2X1 U408 ( .IN1(n86), .IN2(n95), .Q(n426) );
  INVX0 U409 ( .INP(n25), .ZN(n452) );
  FADDX1 U410 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  INVX0 U411 ( .INP(n55), .ZN(n458) );
  INVX0 U412 ( .INP(n73), .ZN(n460) );
  FADDX1 U413 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U414 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  INVX0 U415 ( .INP(n31), .ZN(n454) );
  INVX0 U416 ( .INP(n41), .ZN(n456) );
  INVX0 U417 ( .INP(n492), .ZN(n461) );
  INVX0 U418 ( .INP(n502), .ZN(n459) );
  INVX0 U419 ( .INP(n513), .ZN(n457) );
  INVX0 U420 ( .INP(n524), .ZN(n455) );
  AND2X1 U421 ( .IN1(a[1]), .IN2(n442), .Q(n467) );
  INVX0 U422 ( .INP(n535), .ZN(n453) );
  NBUFFX2 U423 ( .INP(a[5]), .Z(n446) );
  FADDX1 U424 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  NBUFFX2 U425 ( .INP(a[3]), .Z(n444) );
  AND2X1 U426 ( .IN1(n492), .IN2(n547), .Q(n465) );
  AND2X1 U427 ( .IN1(n513), .IN2(n551), .Q(n474) );
  AND2X1 U428 ( .IN1(n502), .IN2(n549), .Q(n471) );
  AND2X1 U429 ( .IN1(n524), .IN2(n553), .Q(n477) );
  AND2X1 U430 ( .IN1(n535), .IN2(n555), .Q(n480) );
  NBUFFX2 U431 ( .INP(a[7]), .Z(n448) );
  NBUFFX2 U432 ( .INP(a[9]), .Z(n450) );
  NAND2X0 U433 ( .IN1(n49), .IN2(n44), .QN(n427) );
  NAND2X0 U434 ( .IN1(n49), .IN2(n10), .QN(n428) );
  NAND2X0 U435 ( .IN1(n44), .IN2(n10), .QN(n429) );
  NAND3X0 U436 ( .IN1(n427), .IN2(n428), .IN3(n429), .QN(n9) );
  NAND2X0 U437 ( .IN1(n43), .IN2(n38), .QN(n430) );
  NAND2X0 U438 ( .IN1(n43), .IN2(n9), .QN(n431) );
  NAND2X0 U439 ( .IN1(n38), .IN2(n9), .QN(n432) );
  NAND3X0 U440 ( .IN1(n432), .IN2(n431), .IN3(n430), .QN(n8) );
  NAND2X0 U441 ( .IN1(n96), .IN2(n103), .QN(n433) );
  NAND2X0 U442 ( .IN1(n96), .IN2(n16), .QN(n434) );
  NAND2X0 U443 ( .IN1(n103), .IN2(n16), .QN(n435) );
  NAND3X0 U444 ( .IN1(n433), .IN2(n434), .IN3(n435), .QN(n15) );
  NAND2X0 U445 ( .IN1(n86), .IN2(n95), .QN(n436) );
  NAND2X0 U446 ( .IN1(n86), .IN2(n15), .QN(n437) );
  NAND2X0 U447 ( .IN1(n95), .IN2(n15), .QN(n438) );
  NAND3X0 U448 ( .IN1(n438), .IN2(n437), .IN3(n436), .QN(n14) );
  DELLN1X2 U449 ( .INP(a[11]), .Z(n451) );
  INVX0 U450 ( .INP(n440), .ZN(n439) );
  INVX0 U451 ( .INP(b[0]), .ZN(n440) );
  INVX0 U452 ( .INP(n442), .ZN(n441) );
  INVX0 U453 ( .INP(a[0]), .ZN(n442) );
  DELLN1X2 U454 ( .INP(a[3]), .Z(n443) );
  DELLN1X2 U455 ( .INP(a[5]), .Z(n445) );
  DELLN1X2 U456 ( .INP(a[7]), .Z(n447) );
  DELLN1X2 U457 ( .INP(a[9]), .Z(n449) );
  NOR2X0 U458 ( .IN1(n442), .IN2(n440), .QN(product[0]) );
  XNOR2X1 U459 ( .IN1(n462), .IN2(n463), .Q(n84) );
  NAND2X0 U460 ( .IN1(n463), .IN2(n462), .QN(n83) );
  AOI22X1 U461 ( .IN1(n464), .IN2(n461), .IN3(n465), .IN4(n466), .QN(n462) );
  OA21X1 U462 ( .IN1(n467), .IN2(n441), .IN3(n468), .Q(n463) );
  AO22X1 U463 ( .IN1(n469), .IN2(n461), .IN3(n465), .IN4(n464), .Q(n73) );
  AO22X1 U464 ( .IN1(n470), .IN2(n459), .IN3(n471), .IN4(n472), .Q(n55) );
  AO22X1 U465 ( .IN1(n473), .IN2(n457), .IN3(n474), .IN4(n475), .Q(n41) );
  AO22X1 U466 ( .IN1(n476), .IN2(n455), .IN3(n477), .IN4(n478), .Q(n31) );
  AO22X1 U467 ( .IN1(n479), .IN2(n453), .IN3(n480), .IN4(n481), .Q(n25) );
  AO22X1 U468 ( .IN1(n441), .IN2(n482), .IN3(n467), .IN4(n440), .Q(n224) );
  AO22X1 U469 ( .IN1(n441), .IN2(n483), .IN3(n467), .IN4(n482), .Q(n223) );
  AO22X1 U470 ( .IN1(n441), .IN2(n484), .IN3(n467), .IN4(n483), .Q(n222) );
  AO22X1 U471 ( .IN1(n441), .IN2(n485), .IN3(n467), .IN4(n484), .Q(n221) );
  AO22X1 U472 ( .IN1(n441), .IN2(n488), .IN3(n467), .IN4(n487), .Q(n218) );
  AO22X1 U473 ( .IN1(n441), .IN2(n489), .IN3(n467), .IN4(n488), .Q(n217) );
  AO22X1 U474 ( .IN1(n441), .IN2(n490), .IN3(n467), .IN4(n489), .Q(n216) );
  AO22X1 U475 ( .IN1(n441), .IN2(n491), .IN3(n467), .IN4(n490), .Q(n215) );
  AO22X1 U476 ( .IN1(n441), .IN2(n468), .IN3(n467), .IN4(n491), .Q(n214) );
  NOR2X0 U477 ( .IN1(n492), .IN2(n440), .QN(n212) );
  AO22X1 U478 ( .IN1(n493), .IN2(n461), .IN3(n465), .IN4(n494), .Q(n211) );
  XOR2X1 U479 ( .IN1(n439), .IN2(n443), .Q(n494) );
  AO22X1 U480 ( .IN1(n495), .IN2(n461), .IN3(n465), .IN4(n493), .Q(n210) );
  AO22X1 U481 ( .IN1(n496), .IN2(n461), .IN3(n465), .IN4(n495), .Q(n209) );
  AO22X1 U482 ( .IN1(n497), .IN2(n461), .IN3(n465), .IN4(n496), .Q(n208) );
  AO22X1 U483 ( .IN1(n498), .IN2(n461), .IN3(n465), .IN4(n497), .Q(n207) );
  AO22X1 U484 ( .IN1(n499), .IN2(n461), .IN3(n465), .IN4(n498), .Q(n206) );
  AO22X1 U485 ( .IN1(n500), .IN2(n461), .IN3(n465), .IN4(n499), .Q(n205) );
  AO22X1 U486 ( .IN1(n501), .IN2(n461), .IN3(n465), .IN4(n500), .Q(n204) );
  AO22X1 U487 ( .IN1(n466), .IN2(n461), .IN3(n465), .IN4(n501), .Q(n203) );
  OAI21X1 U488 ( .IN1(n461), .IN2(n465), .IN3(n469), .QN(n201) );
  NOR2X0 U489 ( .IN1(n502), .IN2(n440), .QN(n200) );
  AO22X1 U490 ( .IN1(n503), .IN2(n459), .IN3(n471), .IN4(n504), .Q(n199) );
  XOR2X1 U491 ( .IN1(n439), .IN2(n445), .Q(n504) );
  AO22X1 U492 ( .IN1(n505), .IN2(n459), .IN3(n471), .IN4(n503), .Q(n198) );
  AO22X1 U493 ( .IN1(n506), .IN2(n459), .IN3(n471), .IN4(n505), .Q(n197) );
  AO22X1 U494 ( .IN1(n507), .IN2(n459), .IN3(n471), .IN4(n506), .Q(n196) );
  AO22X1 U495 ( .IN1(n508), .IN2(n459), .IN3(n471), .IN4(n507), .Q(n195) );
  AO22X1 U496 ( .IN1(n509), .IN2(n459), .IN3(n471), .IN4(n508), .Q(n194) );
  AO22X1 U497 ( .IN1(n510), .IN2(n459), .IN3(n471), .IN4(n509), .Q(n193) );
  AO22X1 U498 ( .IN1(n511), .IN2(n459), .IN3(n471), .IN4(n510), .Q(n192) );
  AO22X1 U499 ( .IN1(n512), .IN2(n459), .IN3(n471), .IN4(n511), .Q(n191) );
  AO22X1 U500 ( .IN1(n472), .IN2(n459), .IN3(n471), .IN4(n512), .Q(n190) );
  OAI21X1 U501 ( .IN1(n459), .IN2(n471), .IN3(n470), .QN(n189) );
  NOR2X0 U502 ( .IN1(n513), .IN2(n440), .QN(n188) );
  AO22X1 U503 ( .IN1(n514), .IN2(n457), .IN3(n474), .IN4(n515), .Q(n187) );
  XOR2X1 U504 ( .IN1(n439), .IN2(n447), .Q(n515) );
  AO22X1 U505 ( .IN1(n516), .IN2(n457), .IN3(n474), .IN4(n514), .Q(n186) );
  AO22X1 U506 ( .IN1(n517), .IN2(n457), .IN3(n474), .IN4(n516), .Q(n185) );
  AO22X1 U507 ( .IN1(n518), .IN2(n457), .IN3(n474), .IN4(n517), .Q(n184) );
  AO22X1 U508 ( .IN1(n519), .IN2(n457), .IN3(n474), .IN4(n518), .Q(n183) );
  AO22X1 U509 ( .IN1(n520), .IN2(n457), .IN3(n474), .IN4(n519), .Q(n182) );
  AO22X1 U510 ( .IN1(n521), .IN2(n457), .IN3(n474), .IN4(n520), .Q(n181) );
  AO22X1 U511 ( .IN1(n522), .IN2(n457), .IN3(n474), .IN4(n521), .Q(n180) );
  AO22X1 U512 ( .IN1(n523), .IN2(n457), .IN3(n474), .IN4(n522), .Q(n179) );
  AO22X1 U513 ( .IN1(n475), .IN2(n457), .IN3(n474), .IN4(n523), .Q(n178) );
  OAI21X1 U514 ( .IN1(n457), .IN2(n474), .IN3(n473), .QN(n177) );
  NOR2X0 U515 ( .IN1(n524), .IN2(n440), .QN(n176) );
  AO22X1 U516 ( .IN1(n525), .IN2(n455), .IN3(n477), .IN4(n526), .Q(n175) );
  XOR2X1 U517 ( .IN1(n439), .IN2(n449), .Q(n526) );
  AO22X1 U518 ( .IN1(n527), .IN2(n455), .IN3(n477), .IN4(n525), .Q(n174) );
  AO22X1 U519 ( .IN1(n528), .IN2(n455), .IN3(n477), .IN4(n527), .Q(n173) );
  AO22X1 U520 ( .IN1(n529), .IN2(n455), .IN3(n477), .IN4(n528), .Q(n172) );
  AO22X1 U521 ( .IN1(n530), .IN2(n455), .IN3(n477), .IN4(n529), .Q(n171) );
  AO22X1 U522 ( .IN1(n531), .IN2(n455), .IN3(n477), .IN4(n530), .Q(n170) );
  AO22X1 U523 ( .IN1(n532), .IN2(n455), .IN3(n477), .IN4(n531), .Q(n169) );
  AO22X1 U524 ( .IN1(n533), .IN2(n455), .IN3(n477), .IN4(n532), .Q(n168) );
  AO22X1 U525 ( .IN1(n534), .IN2(n455), .IN3(n477), .IN4(n533), .Q(n167) );
  AO22X1 U526 ( .IN1(n478), .IN2(n455), .IN3(n477), .IN4(n534), .Q(n166) );
  OAI21X1 U527 ( .IN1(n455), .IN2(n477), .IN3(n476), .QN(n165) );
  NOR2X0 U528 ( .IN1(n535), .IN2(n440), .QN(n164) );
  AO22X1 U529 ( .IN1(n536), .IN2(n453), .IN3(n480), .IN4(n537), .Q(n163) );
  XOR2X1 U530 ( .IN1(n439), .IN2(n451), .Q(n537) );
  AO22X1 U531 ( .IN1(n538), .IN2(n453), .IN3(n480), .IN4(n536), .Q(n162) );
  AO22X1 U532 ( .IN1(n539), .IN2(n453), .IN3(n480), .IN4(n538), .Q(n161) );
  AO22X1 U533 ( .IN1(n540), .IN2(n453), .IN3(n480), .IN4(n539), .Q(n160) );
  AO22X1 U534 ( .IN1(n541), .IN2(n453), .IN3(n480), .IN4(n540), .Q(n159) );
  AO22X1 U535 ( .IN1(n542), .IN2(n453), .IN3(n480), .IN4(n541), .Q(n158) );
  AO22X1 U536 ( .IN1(n543), .IN2(n453), .IN3(n480), .IN4(n542), .Q(n157) );
  AO22X1 U537 ( .IN1(n544), .IN2(n453), .IN3(n480), .IN4(n543), .Q(n156) );
  AO22X1 U538 ( .IN1(n545), .IN2(n453), .IN3(n480), .IN4(n544), .Q(n155) );
  AO22X1 U539 ( .IN1(n481), .IN2(n453), .IN3(n480), .IN4(n545), .Q(n154) );
  OAI21X1 U540 ( .IN1(n453), .IN2(n480), .IN3(n479), .QN(n153) );
  AO21X1 U541 ( .IN1(a[1]), .IN2(n440), .IN3(n467), .Q(n152) );
  AO22X1 U542 ( .IN1(n546), .IN2(n444), .IN3(n465), .IN4(n444), .Q(n151) );
  XOR2X1 U543 ( .IN1(n443), .IN2(a[2]), .Q(n547) );
  NOR2X0 U544 ( .IN1(n439), .IN2(n492), .QN(n546) );
  XNOR2X1 U545 ( .IN1(a[2]), .IN2(a[1]), .Q(n492) );
  AO22X1 U546 ( .IN1(n548), .IN2(n446), .IN3(n471), .IN4(n446), .Q(n150) );
  XOR2X1 U547 ( .IN1(n445), .IN2(a[4]), .Q(n549) );
  NOR2X0 U548 ( .IN1(n439), .IN2(n502), .QN(n548) );
  XNOR2X1 U549 ( .IN1(a[4]), .IN2(n443), .Q(n502) );
  AO22X1 U550 ( .IN1(n550), .IN2(n448), .IN3(n474), .IN4(n448), .Q(n149) );
  XOR2X1 U551 ( .IN1(n447), .IN2(a[6]), .Q(n551) );
  NOR2X0 U552 ( .IN1(n439), .IN2(n513), .QN(n550) );
  XNOR2X1 U553 ( .IN1(a[6]), .IN2(n445), .Q(n513) );
  AO22X1 U554 ( .IN1(n552), .IN2(n450), .IN3(n477), .IN4(n450), .Q(n148) );
  XOR2X1 U555 ( .IN1(n449), .IN2(a[8]), .Q(n553) );
  NOR2X0 U556 ( .IN1(n439), .IN2(n524), .QN(n552) );
  XNOR2X1 U557 ( .IN1(a[8]), .IN2(n447), .Q(n524) );
  AO22X1 U558 ( .IN1(n554), .IN2(n451), .IN3(n480), .IN4(n451), .Q(n147) );
  XOR2X1 U559 ( .IN1(n451), .IN2(a[10]), .Q(n555) );
  NOR2X0 U560 ( .IN1(n439), .IN2(n535), .QN(n554) );
  XNOR2X1 U561 ( .IN1(a[10]), .IN2(n449), .Q(n535) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_13 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_13_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_12_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n456), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n458), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n460), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n462), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  DELLN1X2 U311 ( .INP(b[2]), .Z(n408) );
  DELLN1X2 U312 ( .INP(b[7]), .Z(n409) );
  FADDX1 U313 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U314 ( .A(n27), .B(n454), .CI(n5), .CO(n4), .S(product[21]) );
  DELLN1X2 U315 ( .INP(b[1]), .Z(n410) );
  INVX0 U316 ( .INP(b[8]), .ZN(n411) );
  INVX0 U317 ( .INP(n411), .ZN(n412) );
  DELLN2X2 U318 ( .INP(n12), .Z(n413) );
  INVX0 U319 ( .INP(b[6]), .ZN(n414) );
  INVX0 U320 ( .INP(n414), .ZN(n415) );
  INVX0 U321 ( .INP(b[5]), .ZN(n416) );
  INVX0 U322 ( .INP(n416), .ZN(n417) );
  XOR2X2 U323 ( .IN1(b[10]), .IN2(n452), .Q(n483) );
  XOR2X2 U324 ( .IN1(b[10]), .IN2(n450), .Q(n480) );
  XOR2X2 U325 ( .IN1(b[10]), .IN2(n448), .Q(n477) );
  XOR2X2 U326 ( .IN1(b[10]), .IN2(n446), .Q(n474) );
  XOR2X2 U327 ( .IN1(b[10]), .IN2(n444), .Q(n466) );
  XOR2X2 U328 ( .IN1(n412), .IN2(n452), .Q(n546) );
  XOR2X2 U329 ( .IN1(n412), .IN2(n450), .Q(n535) );
  XOR2X2 U330 ( .IN1(n412), .IN2(n448), .Q(n524) );
  XOR2X2 U331 ( .IN1(n412), .IN2(n446), .Q(n513) );
  XOR2X2 U332 ( .IN1(n412), .IN2(n444), .Q(n503) );
  XOR2X2 U333 ( .IN1(n412), .IN2(a[1]), .Q(n491) );
  XOR2X2 U334 ( .IN1(n415), .IN2(n452), .Q(n544) );
  XOR2X2 U335 ( .IN1(n415), .IN2(n450), .Q(n533) );
  XOR2X2 U336 ( .IN1(n415), .IN2(n448), .Q(n522) );
  XOR2X2 U337 ( .IN1(n415), .IN2(n446), .Q(n511) );
  XOR2X2 U338 ( .IN1(n415), .IN2(n444), .Q(n501) );
  XOR2X2 U339 ( .IN1(n417), .IN2(n452), .Q(n543) );
  XOR2X2 U340 ( .IN1(n417), .IN2(n450), .Q(n532) );
  XOR2X2 U341 ( .IN1(n417), .IN2(n448), .Q(n521) );
  XOR2X2 U342 ( .IN1(n417), .IN2(n446), .Q(n510) );
  XOR2X2 U343 ( .IN1(n417), .IN2(n444), .Q(n500) );
  XOR3X1 U344 ( .IN1(n66), .IN2(n75), .IN3(n13), .Q(product[13]) );
  NAND2X0 U345 ( .IN1(n66), .IN2(n75), .QN(n418) );
  NAND2X0 U346 ( .IN1(n65), .IN2(n58), .QN(n422) );
  XOR2X1 U347 ( .IN1(n132), .IN2(n133), .Q(n435) );
  NAND2X0 U348 ( .IN1(n151), .IN2(n23), .QN(n434) );
  NAND2X0 U349 ( .IN1(n66), .IN2(n13), .QN(n419) );
  NAND2X0 U350 ( .IN1(n75), .IN2(n13), .QN(n420) );
  NAND3X0 U351 ( .IN1(n418), .IN2(n419), .IN3(n420), .QN(n12) );
  XOR2X1 U352 ( .IN1(n65), .IN2(n58), .Q(n421) );
  XOR2X1 U353 ( .IN1(n421), .IN2(n413), .Q(product[14]) );
  NAND2X0 U354 ( .IN1(n65), .IN2(n12), .QN(n423) );
  NAND2X0 U355 ( .IN1(n58), .IN2(n12), .QN(n424) );
  NAND3X0 U356 ( .IN1(n422), .IN2(n423), .IN3(n424), .QN(n11) );
  XOR3X1 U357 ( .IN1(n124), .IN2(n127), .IN3(n20), .Q(product[6]) );
  NAND2X0 U358 ( .IN1(n124), .IN2(n127), .QN(n425) );
  NAND2X0 U359 ( .IN1(n124), .IN2(n20), .QN(n426) );
  NAND2X0 U360 ( .IN1(n127), .IN2(n20), .QN(n427) );
  NAND3X0 U361 ( .IN1(n425), .IN2(n426), .IN3(n427), .QN(n19) );
  XOR2X1 U362 ( .IN1(n118), .IN2(n123), .Q(n428) );
  XOR2X1 U363 ( .IN1(n428), .IN2(n19), .Q(product[7]) );
  NAND2X0 U364 ( .IN1(n118), .IN2(n123), .QN(n429) );
  NAND2X0 U365 ( .IN1(n118), .IN2(n19), .QN(n430) );
  NAND2X0 U366 ( .IN1(n123), .IN2(n19), .QN(n431) );
  NAND3X0 U367 ( .IN1(n429), .IN2(n430), .IN3(n431), .QN(n18) );
  XOR3X1 U368 ( .IN1(n134), .IN2(n151), .IN3(n23), .Q(product[3]) );
  NAND2X0 U369 ( .IN1(n134), .IN2(n151), .QN(n432) );
  NAND2X0 U370 ( .IN1(n134), .IN2(n23), .QN(n433) );
  NAND3X0 U371 ( .IN1(n432), .IN2(n433), .IN3(n434), .QN(n22) );
  XOR2X1 U372 ( .IN1(n435), .IN2(n22), .Q(product[4]) );
  NAND2X0 U373 ( .IN1(n132), .IN2(n133), .QN(n436) );
  NAND2X0 U374 ( .IN1(n132), .IN2(n22), .QN(n437) );
  NAND2X0 U375 ( .IN1(n133), .IN2(n22), .QN(n438) );
  NAND3X0 U376 ( .IN1(n436), .IN2(n437), .IN3(n438), .QN(n21) );
  FADDX1 U377 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U378 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  INVX0 U379 ( .INP(n25), .ZN(n454) );
  INVX0 U380 ( .INP(n3), .ZN(product[23]) );
  INVX0 U381 ( .INP(n55), .ZN(n460) );
  XOR2X1 U382 ( .IN1(n410), .IN2(n444), .Q(n495) );
  INVX0 U383 ( .INP(n73), .ZN(n462) );
  XOR2X1 U384 ( .IN1(n410), .IN2(n448), .Q(n516) );
  XOR2X1 U385 ( .IN1(n410), .IN2(n450), .Q(n527) );
  XOR2X1 U386 ( .IN1(n410), .IN2(n446), .Q(n505) );
  XOR2X1 U387 ( .IN1(b[3]), .IN2(n448), .Q(n519) );
  XOR2X1 U388 ( .IN1(n410), .IN2(n452), .Q(n538) );
  XOR2X1 U389 ( .IN1(b[3]), .IN2(n450), .Q(n530) );
  XOR2X1 U390 ( .IN1(b[3]), .IN2(n452), .Q(n541) );
  INVX0 U391 ( .INP(n31), .ZN(n456) );
  INVX0 U392 ( .INP(n41), .ZN(n458) );
  INVX0 U393 ( .INP(n504), .ZN(n461) );
  INVX0 U394 ( .INP(n494), .ZN(n463) );
  AND2X1 U395 ( .IN1(a[1]), .IN2(n443), .Q(n469) );
  INVX0 U396 ( .INP(n515), .ZN(n459) );
  INVX0 U397 ( .INP(n526), .ZN(n457) );
  INVX0 U398 ( .INP(n537), .ZN(n455) );
  NBUFFX2 U399 ( .INP(a[3]), .Z(n445) );
  FADDX1 U400 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  NBUFFX2 U401 ( .INP(a[5]), .Z(n447) );
  NBUFFX2 U402 ( .INP(a[9]), .Z(n451) );
  XOR2X2 U403 ( .IN1(b[3]), .IN2(n446), .Q(n508) );
  XOR2X2 U404 ( .IN1(b[3]), .IN2(n444), .Q(n498) );
  XOR2X2 U405 ( .IN1(b[3]), .IN2(a[1]), .Q(n486) );
  XOR2X2 U406 ( .IN1(n410), .IN2(a[1]), .Q(n484) );
  XOR2X2 U407 ( .IN1(b[10]), .IN2(a[1]), .Q(n493) );
  XOR2X2 U408 ( .IN1(n409), .IN2(a[1]), .Q(n490) );
  XOR2X2 U409 ( .IN1(n417), .IN2(a[1]), .Q(n488) );
  XOR2X2 U410 ( .IN1(n415), .IN2(a[1]), .Q(n489) );
  FADDX1 U411 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X2 U412 ( .IN1(b[4]), .IN2(a[1]), .Q(n487) );
  XOR2X2 U413 ( .IN1(n408), .IN2(a[1]), .Q(n485) );
  DELLN1X2 U414 ( .INP(a[11]), .Z(n452) );
  AND2X2 U415 ( .IN1(n494), .IN2(n549), .Q(n467) );
  AND2X2 U416 ( .IN1(n504), .IN2(n551), .Q(n473) );
  AND2X2 U417 ( .IN1(n515), .IN2(n553), .Q(n476) );
  AND2X2 U418 ( .IN1(n526), .IN2(n555), .Q(n479) );
  AND2X2 U419 ( .IN1(n537), .IN2(n557), .Q(n482) );
  INVX0 U420 ( .INP(n441), .ZN(n439) );
  INVX0 U421 ( .INP(b[0]), .ZN(n440) );
  INVX0 U422 ( .INP(b[0]), .ZN(n441) );
  INVX0 U423 ( .INP(n443), .ZN(n442) );
  INVX0 U424 ( .INP(a[0]), .ZN(n443) );
  DELLN1X2 U425 ( .INP(a[3]), .Z(n444) );
  DELLN1X2 U426 ( .INP(a[5]), .Z(n446) );
  DELLN1X2 U427 ( .INP(a[7]), .Z(n448) );
  DELLN1X2 U428 ( .INP(a[7]), .Z(n449) );
  DELLN1X2 U429 ( .INP(a[9]), .Z(n450) );
  NOR2X0 U430 ( .IN1(n443), .IN2(n440), .QN(product[0]) );
  XNOR2X1 U431 ( .IN1(n464), .IN2(n465), .Q(n84) );
  NAND2X0 U432 ( .IN1(n465), .IN2(n464), .QN(n83) );
  AOI22X1 U433 ( .IN1(n466), .IN2(n463), .IN3(n467), .IN4(n468), .QN(n464) );
  OA21X1 U434 ( .IN1(n469), .IN2(n442), .IN3(n470), .Q(n465) );
  AO22X1 U435 ( .IN1(n471), .IN2(n463), .IN3(n467), .IN4(n466), .Q(n73) );
  AO22X1 U436 ( .IN1(n472), .IN2(n461), .IN3(n473), .IN4(n474), .Q(n55) );
  AO22X1 U437 ( .IN1(n475), .IN2(n459), .IN3(n476), .IN4(n477), .Q(n41) );
  AO22X1 U438 ( .IN1(n478), .IN2(n457), .IN3(n479), .IN4(n480), .Q(n31) );
  AO22X1 U439 ( .IN1(n481), .IN2(n455), .IN3(n482), .IN4(n483), .Q(n25) );
  AO22X1 U440 ( .IN1(n442), .IN2(n484), .IN3(n469), .IN4(n441), .Q(n224) );
  AO22X1 U441 ( .IN1(n442), .IN2(n485), .IN3(n469), .IN4(n484), .Q(n223) );
  AO22X1 U442 ( .IN1(n442), .IN2(n486), .IN3(n469), .IN4(n485), .Q(n222) );
  AO22X1 U443 ( .IN1(n442), .IN2(n487), .IN3(n469), .IN4(n486), .Q(n221) );
  AO22X1 U444 ( .IN1(n442), .IN2(n488), .IN3(n469), .IN4(n487), .Q(n220) );
  AO22X1 U445 ( .IN1(n442), .IN2(n489), .IN3(n469), .IN4(n488), .Q(n219) );
  AO22X1 U446 ( .IN1(n442), .IN2(n490), .IN3(n469), .IN4(n489), .Q(n218) );
  AO22X1 U447 ( .IN1(n442), .IN2(n491), .IN3(n469), .IN4(n490), .Q(n217) );
  AO22X1 U448 ( .IN1(n442), .IN2(n492), .IN3(n469), .IN4(n491), .Q(n216) );
  AO22X1 U449 ( .IN1(n442), .IN2(n493), .IN3(n469), .IN4(n492), .Q(n215) );
  XOR2X1 U450 ( .IN1(b[9]), .IN2(a[1]), .Q(n492) );
  AO22X1 U451 ( .IN1(n442), .IN2(n470), .IN3(n469), .IN4(n493), .Q(n214) );
  XOR2X1 U452 ( .IN1(b[11]), .IN2(a[1]), .Q(n470) );
  NOR2X0 U453 ( .IN1(n494), .IN2(n440), .QN(n212) );
  AO22X1 U454 ( .IN1(n495), .IN2(n463), .IN3(n467), .IN4(n496), .Q(n211) );
  XOR2X1 U455 ( .IN1(n439), .IN2(n444), .Q(n496) );
  AO22X1 U456 ( .IN1(n497), .IN2(n463), .IN3(n467), .IN4(n495), .Q(n210) );
  AO22X1 U457 ( .IN1(n498), .IN2(n463), .IN3(n467), .IN4(n497), .Q(n209) );
  XOR2X1 U458 ( .IN1(n408), .IN2(n444), .Q(n497) );
  AO22X1 U459 ( .IN1(n499), .IN2(n463), .IN3(n467), .IN4(n498), .Q(n208) );
  AO22X1 U460 ( .IN1(n500), .IN2(n463), .IN3(n467), .IN4(n499), .Q(n207) );
  XOR2X1 U461 ( .IN1(b[4]), .IN2(n444), .Q(n499) );
  AO22X1 U462 ( .IN1(n501), .IN2(n463), .IN3(n467), .IN4(n500), .Q(n206) );
  AO22X1 U463 ( .IN1(n502), .IN2(n463), .IN3(n467), .IN4(n501), .Q(n205) );
  AO22X1 U464 ( .IN1(n503), .IN2(n463), .IN3(n467), .IN4(n502), .Q(n204) );
  XOR2X1 U465 ( .IN1(n409), .IN2(n444), .Q(n502) );
  AO22X1 U466 ( .IN1(n468), .IN2(n463), .IN3(n467), .IN4(n503), .Q(n203) );
  XOR2X1 U467 ( .IN1(b[9]), .IN2(n444), .Q(n468) );
  OAI21X1 U468 ( .IN1(n463), .IN2(n467), .IN3(n471), .QN(n201) );
  XOR2X1 U469 ( .IN1(b[11]), .IN2(n444), .Q(n471) );
  NOR2X0 U470 ( .IN1(n504), .IN2(n440), .QN(n200) );
  AO22X1 U471 ( .IN1(n505), .IN2(n461), .IN3(n473), .IN4(n506), .Q(n199) );
  XOR2X1 U472 ( .IN1(n439), .IN2(n446), .Q(n506) );
  AO22X1 U473 ( .IN1(n507), .IN2(n461), .IN3(n473), .IN4(n505), .Q(n198) );
  AO22X1 U474 ( .IN1(n508), .IN2(n461), .IN3(n473), .IN4(n507), .Q(n197) );
  XOR2X1 U475 ( .IN1(n408), .IN2(n446), .Q(n507) );
  AO22X1 U476 ( .IN1(n509), .IN2(n461), .IN3(n473), .IN4(n508), .Q(n196) );
  AO22X1 U477 ( .IN1(n510), .IN2(n461), .IN3(n473), .IN4(n509), .Q(n195) );
  XOR2X1 U478 ( .IN1(b[4]), .IN2(n446), .Q(n509) );
  AO22X1 U479 ( .IN1(n511), .IN2(n461), .IN3(n473), .IN4(n510), .Q(n194) );
  AO22X1 U480 ( .IN1(n512), .IN2(n461), .IN3(n473), .IN4(n511), .Q(n193) );
  AO22X1 U481 ( .IN1(n513), .IN2(n461), .IN3(n473), .IN4(n512), .Q(n192) );
  XOR2X1 U482 ( .IN1(n409), .IN2(n446), .Q(n512) );
  AO22X1 U483 ( .IN1(n514), .IN2(n461), .IN3(n473), .IN4(n513), .Q(n191) );
  AO22X1 U484 ( .IN1(n474), .IN2(n461), .IN3(n473), .IN4(n514), .Q(n190) );
  XOR2X1 U485 ( .IN1(b[9]), .IN2(n446), .Q(n514) );
  OAI21X1 U486 ( .IN1(n461), .IN2(n473), .IN3(n472), .QN(n189) );
  XOR2X1 U487 ( .IN1(b[11]), .IN2(n446), .Q(n472) );
  NOR2X0 U488 ( .IN1(n515), .IN2(n440), .QN(n188) );
  AO22X1 U489 ( .IN1(n516), .IN2(n459), .IN3(n476), .IN4(n517), .Q(n187) );
  XOR2X1 U490 ( .IN1(n439), .IN2(n448), .Q(n517) );
  AO22X1 U491 ( .IN1(n518), .IN2(n459), .IN3(n476), .IN4(n516), .Q(n186) );
  AO22X1 U492 ( .IN1(n519), .IN2(n459), .IN3(n476), .IN4(n518), .Q(n185) );
  XOR2X1 U493 ( .IN1(n408), .IN2(n448), .Q(n518) );
  AO22X1 U494 ( .IN1(n520), .IN2(n459), .IN3(n476), .IN4(n519), .Q(n184) );
  AO22X1 U495 ( .IN1(n521), .IN2(n459), .IN3(n476), .IN4(n520), .Q(n183) );
  XOR2X1 U496 ( .IN1(b[4]), .IN2(n448), .Q(n520) );
  AO22X1 U497 ( .IN1(n522), .IN2(n459), .IN3(n476), .IN4(n521), .Q(n182) );
  AO22X1 U498 ( .IN1(n523), .IN2(n459), .IN3(n476), .IN4(n522), .Q(n181) );
  AO22X1 U499 ( .IN1(n524), .IN2(n459), .IN3(n476), .IN4(n523), .Q(n180) );
  XOR2X1 U500 ( .IN1(n409), .IN2(n448), .Q(n523) );
  AO22X1 U501 ( .IN1(n525), .IN2(n459), .IN3(n476), .IN4(n524), .Q(n179) );
  AO22X1 U502 ( .IN1(n477), .IN2(n459), .IN3(n476), .IN4(n525), .Q(n178) );
  XOR2X1 U503 ( .IN1(b[9]), .IN2(n448), .Q(n525) );
  OAI21X1 U504 ( .IN1(n459), .IN2(n476), .IN3(n475), .QN(n177) );
  XOR2X1 U505 ( .IN1(b[11]), .IN2(n448), .Q(n475) );
  NOR2X0 U506 ( .IN1(n526), .IN2(n440), .QN(n176) );
  AO22X1 U507 ( .IN1(n527), .IN2(n457), .IN3(n479), .IN4(n528), .Q(n175) );
  XOR2X1 U508 ( .IN1(n439), .IN2(n450), .Q(n528) );
  AO22X1 U509 ( .IN1(n529), .IN2(n457), .IN3(n479), .IN4(n527), .Q(n174) );
  AO22X1 U510 ( .IN1(n530), .IN2(n457), .IN3(n479), .IN4(n529), .Q(n173) );
  XOR2X1 U511 ( .IN1(n408), .IN2(n450), .Q(n529) );
  AO22X1 U512 ( .IN1(n531), .IN2(n457), .IN3(n479), .IN4(n530), .Q(n172) );
  AO22X1 U513 ( .IN1(n532), .IN2(n457), .IN3(n479), .IN4(n531), .Q(n171) );
  XOR2X1 U514 ( .IN1(b[4]), .IN2(n450), .Q(n531) );
  AO22X1 U515 ( .IN1(n533), .IN2(n457), .IN3(n479), .IN4(n532), .Q(n170) );
  AO22X1 U516 ( .IN1(n534), .IN2(n457), .IN3(n479), .IN4(n533), .Q(n169) );
  AO22X1 U517 ( .IN1(n535), .IN2(n457), .IN3(n479), .IN4(n534), .Q(n168) );
  XOR2X1 U518 ( .IN1(n409), .IN2(n450), .Q(n534) );
  AO22X1 U519 ( .IN1(n536), .IN2(n457), .IN3(n479), .IN4(n535), .Q(n167) );
  AO22X1 U520 ( .IN1(n480), .IN2(n457), .IN3(n479), .IN4(n536), .Q(n166) );
  XOR2X1 U521 ( .IN1(b[9]), .IN2(n450), .Q(n536) );
  OAI21X1 U522 ( .IN1(n457), .IN2(n479), .IN3(n478), .QN(n165) );
  XOR2X1 U523 ( .IN1(b[11]), .IN2(n450), .Q(n478) );
  NOR2X0 U524 ( .IN1(n537), .IN2(n440), .QN(n164) );
  AO22X1 U525 ( .IN1(n538), .IN2(n455), .IN3(n482), .IN4(n539), .Q(n163) );
  XOR2X1 U526 ( .IN1(n439), .IN2(n452), .Q(n539) );
  AO22X1 U527 ( .IN1(n540), .IN2(n455), .IN3(n482), .IN4(n538), .Q(n162) );
  AO22X1 U528 ( .IN1(n541), .IN2(n455), .IN3(n482), .IN4(n540), .Q(n161) );
  XOR2X1 U529 ( .IN1(n408), .IN2(n452), .Q(n540) );
  AO22X1 U530 ( .IN1(n542), .IN2(n455), .IN3(n482), .IN4(n541), .Q(n160) );
  AO22X1 U531 ( .IN1(n543), .IN2(n455), .IN3(n482), .IN4(n542), .Q(n159) );
  XOR2X1 U532 ( .IN1(b[4]), .IN2(n452), .Q(n542) );
  AO22X1 U533 ( .IN1(n544), .IN2(n455), .IN3(n482), .IN4(n543), .Q(n158) );
  AO22X1 U534 ( .IN1(n545), .IN2(n455), .IN3(n482), .IN4(n544), .Q(n157) );
  AO22X1 U535 ( .IN1(n546), .IN2(n455), .IN3(n482), .IN4(n545), .Q(n156) );
  XOR2X1 U536 ( .IN1(n409), .IN2(n452), .Q(n545) );
  AO22X1 U537 ( .IN1(n547), .IN2(n455), .IN3(n482), .IN4(n546), .Q(n155) );
  AO22X1 U538 ( .IN1(n483), .IN2(n455), .IN3(n482), .IN4(n547), .Q(n154) );
  XOR2X1 U539 ( .IN1(b[9]), .IN2(n452), .Q(n547) );
  OAI21X1 U540 ( .IN1(n455), .IN2(n482), .IN3(n481), .QN(n153) );
  XOR2X1 U541 ( .IN1(b[11]), .IN2(n452), .Q(n481) );
  AO21X1 U542 ( .IN1(a[1]), .IN2(n441), .IN3(n469), .Q(n152) );
  AO22X1 U543 ( .IN1(n548), .IN2(n445), .IN3(n467), .IN4(n445), .Q(n151) );
  XOR2X1 U544 ( .IN1(n444), .IN2(a[2]), .Q(n549) );
  NOR2X0 U545 ( .IN1(n439), .IN2(n494), .QN(n548) );
  XNOR2X1 U546 ( .IN1(a[2]), .IN2(a[1]), .Q(n494) );
  AO22X1 U547 ( .IN1(n550), .IN2(n447), .IN3(n473), .IN4(n447), .Q(n150) );
  XOR2X1 U548 ( .IN1(n446), .IN2(a[4]), .Q(n551) );
  NOR2X0 U549 ( .IN1(n439), .IN2(n504), .QN(n550) );
  XNOR2X1 U550 ( .IN1(a[4]), .IN2(n444), .Q(n504) );
  AO22X1 U551 ( .IN1(n552), .IN2(n449), .IN3(n476), .IN4(n449), .Q(n149) );
  XOR2X1 U552 ( .IN1(n448), .IN2(a[6]), .Q(n553) );
  NOR2X0 U553 ( .IN1(n439), .IN2(n515), .QN(n552) );
  XNOR2X1 U554 ( .IN1(a[6]), .IN2(n446), .Q(n515) );
  AO22X1 U555 ( .IN1(n554), .IN2(n451), .IN3(n479), .IN4(n451), .Q(n148) );
  XOR2X1 U556 ( .IN1(n450), .IN2(a[8]), .Q(n555) );
  NOR2X0 U557 ( .IN1(n439), .IN2(n526), .QN(n554) );
  XNOR2X1 U558 ( .IN1(a[8]), .IN2(n448), .Q(n526) );
  AO22X1 U559 ( .IN1(n556), .IN2(n452), .IN3(n482), .IN4(n452), .Q(n147) );
  XOR2X1 U560 ( .IN1(n452), .IN2(a[10]), .Q(n557) );
  NOR2X0 U561 ( .IN1(n439), .IN2(n537), .QN(n556) );
  XNOR2X1 U562 ( .IN1(a[10]), .IN2(n450), .Q(n537) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_12 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_12_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_3_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [24:0] carry;

  FADDX1 U2_22 ( .A(A[22]), .B(n7), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n8), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n9), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n10), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n11), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n12), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n13), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n18), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n21), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n22), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XNOR3X1 U1 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(DIFF[23]) );
  INVX0 U2 ( .INP(B[21]), .ZN(n8) );
  INVX0 U3 ( .INP(B[20]), .ZN(n9) );
  INVX0 U4 ( .INP(B[22]), .ZN(n7) );
  INVX0 U5 ( .INP(B[19]), .ZN(n10) );
  INVX0 U6 ( .INP(B[18]), .ZN(n11) );
  INVX0 U7 ( .INP(B[17]), .ZN(n12) );
  INVX0 U8 ( .INP(B[16]), .ZN(n13) );
  INVX0 U9 ( .INP(B[15]), .ZN(n14) );
  INVX0 U10 ( .INP(B[14]), .ZN(n15) );
  INVX0 U11 ( .INP(B[13]), .ZN(n16) );
  INVX0 U12 ( .INP(B[12]), .ZN(n17) );
  INVX0 U13 ( .INP(B[11]), .ZN(n18) );
  INVX0 U14 ( .INP(B[10]), .ZN(n19) );
  INVX0 U15 ( .INP(B[9]), .ZN(n20) );
  INVX0 U16 ( .INP(B[8]), .ZN(n21) );
  INVX0 U17 ( .INP(B[7]), .ZN(n22) );
  INVX0 U18 ( .INP(A[3]), .ZN(n4) );
  INVX0 U19 ( .INP(A[1]), .ZN(n6) );
  INVX0 U20 ( .INP(A[5]), .ZN(n2) );
  INVX0 U21 ( .INP(A[2]), .ZN(n5) );
  INVX0 U22 ( .INP(B[0]), .ZN(n23) );
  INVX0 U23 ( .INP(A[4]), .ZN(n3) );
  INVX0 U24 ( .INP(A[6]), .ZN(n1) );
  OAI22X1 U25 ( .IN1(n24), .IN2(n1), .IN3(B[6]), .IN4(n25), .QN(carry[7]) );
  AND2X1 U26 ( .IN1(n1), .IN2(n24), .Q(n25) );
  OA22X1 U27 ( .IN1(n26), .IN2(n2), .IN3(B[5]), .IN4(n27), .Q(n24) );
  AND2X1 U28 ( .IN1(n2), .IN2(n26), .Q(n27) );
  OA22X1 U29 ( .IN1(n28), .IN2(n3), .IN3(B[4]), .IN4(n29), .Q(n26) );
  AND2X1 U30 ( .IN1(n3), .IN2(n28), .Q(n29) );
  OA22X1 U31 ( .IN1(n30), .IN2(n4), .IN3(B[3]), .IN4(n31), .Q(n28) );
  AND2X1 U32 ( .IN1(n4), .IN2(n30), .Q(n31) );
  OA22X1 U33 ( .IN1(n32), .IN2(n5), .IN3(B[2]), .IN4(n33), .Q(n30) );
  AND2X1 U34 ( .IN1(n5), .IN2(n32), .Q(n33) );
  OA22X1 U35 ( .IN1(n34), .IN2(n6), .IN3(B[1]), .IN4(n35), .Q(n32) );
  AND2X1 U36 ( .IN1(n6), .IN2(n34), .Q(n35) );
  NOR2X0 U37 ( .IN1(n23), .IN2(A[0]), .QN(n34) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_3 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_3_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(\output ) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_3_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AO22X1 U1 ( .IN1(A[6]), .IN2(n1), .IN3(B[6]), .IN4(n2), .Q(carry[7]) );
  OR2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AO22X1 U3 ( .IN1(A[5]), .IN2(n3), .IN3(B[5]), .IN4(n4), .Q(n1) );
  OR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AO22X1 U5 ( .IN1(A[4]), .IN2(n5), .IN3(B[4]), .IN4(n6), .Q(n3) );
  OR2X1 U6 ( .IN1(n5), .IN2(A[4]), .Q(n6) );
  AO22X1 U7 ( .IN1(A[3]), .IN2(n7), .IN3(B[3]), .IN4(n8), .Q(n5) );
  OR2X1 U8 ( .IN1(n7), .IN2(A[3]), .Q(n8) );
  AO22X1 U9 ( .IN1(A[2]), .IN2(n9), .IN3(B[2]), .IN4(n10), .Q(n7) );
  OR2X1 U10 ( .IN1(n9), .IN2(A[2]), .Q(n10) );
  AO22X1 U11 ( .IN1(B[1]), .IN2(A[1]), .IN3(n11), .IN4(B[0]), .Q(n9) );
  OA21X1 U12 ( .IN1(A[1]), .IN2(B[1]), .IN3(A[0]), .Q(n11) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_3 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_3_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(\output ) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3 ( a_r, a_i, b_r, b_i, out_r, 
        out_i, clk );
  input [11:0] a_r;
  input [11:0] a_i;
  input [11:0] b_r;
  input [11:0] b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37;
  wire   [23:0] mult1_out;
  wire   [23:0] mult2_out;
  wire   [23:0] mult3_out;
  wire   [23:0] mult4_out;
  wire   [23:7] pre_out_r;
  wire   [23:7] pre_out_i;
  wire   [11:0] rnd_out_r;
  wire   [11:0] rnd_out_i;
  wire   [11:0] pos_out_r;
  wire   [11:0] pos_out_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFFX1 \out_r_reg_reg[11]  ( .D(pos_out_r[11]), .CLK(clk), .Q(out_r[11]) );
  DFFX1 \out_r_reg_reg[10]  ( .D(pos_out_r[10]), .CLK(clk), .Q(out_r[10]) );
  DFFX1 \out_r_reg_reg[9]  ( .D(pos_out_r[9]), .CLK(clk), .Q(out_r[9]) );
  DFFX1 \out_r_reg_reg[8]  ( .D(pos_out_r[8]), .CLK(clk), .Q(out_r[8]) );
  DFFX1 \out_r_reg_reg[7]  ( .D(pos_out_r[7]), .CLK(clk), .Q(out_r[7]) );
  DFFX1 \out_r_reg_reg[6]  ( .D(pos_out_r[6]), .CLK(clk), .Q(out_r[6]) );
  DFFX1 \out_r_reg_reg[5]  ( .D(pos_out_r[5]), .CLK(clk), .Q(out_r[5]) );
  DFFX1 \out_r_reg_reg[4]  ( .D(pos_out_r[4]), .CLK(clk), .Q(out_r[4]) );
  DFFX1 \out_r_reg_reg[3]  ( .D(pos_out_r[3]), .CLK(clk), .Q(out_r[3]) );
  DFFX1 \out_r_reg_reg[2]  ( .D(pos_out_r[2]), .CLK(clk), .Q(out_r[2]) );
  DFFX1 \out_r_reg_reg[1]  ( .D(pos_out_r[1]), .CLK(clk), .Q(out_r[1]) );
  DFFX1 \out_r_reg_reg[0]  ( .D(pos_out_r[0]), .CLK(clk), .Q(out_r[0]) );
  DFFX1 \out_i_reg_reg[11]  ( .D(pos_out_i[11]), .CLK(clk), .Q(out_i[11]) );
  DFFX1 \out_i_reg_reg[10]  ( .D(pos_out_i[10]), .CLK(clk), .Q(out_i[10]) );
  DFFX1 \out_i_reg_reg[9]  ( .D(pos_out_i[9]), .CLK(clk), .Q(out_i[9]) );
  DFFX1 \out_i_reg_reg[8]  ( .D(pos_out_i[8]), .CLK(clk), .Q(out_i[8]) );
  DFFX1 \out_i_reg_reg[7]  ( .D(pos_out_i[7]), .CLK(clk), .Q(out_i[7]) );
  DFFX1 \out_i_reg_reg[6]  ( .D(pos_out_i[6]), .CLK(clk), .Q(out_i[6]) );
  DFFX1 \out_i_reg_reg[5]  ( .D(pos_out_i[5]), .CLK(clk), .Q(out_i[5]) );
  DFFX1 \out_i_reg_reg[4]  ( .D(pos_out_i[4]), .CLK(clk), .Q(out_i[4]) );
  DFFX1 \out_i_reg_reg[3]  ( .D(pos_out_i[3]), .CLK(clk), .Q(out_i[3]) );
  DFFX1 \out_i_reg_reg[2]  ( .D(pos_out_i[2]), .CLK(clk), .Q(out_i[2]) );
  DFFX1 \out_i_reg_reg[1]  ( .D(pos_out_i[1]), .CLK(clk), .Q(out_i[1]) );
  DFFX1 \out_i_reg_reg[0]  ( .D(pos_out_i[0]), .CLK(clk), .Q(out_i[0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_15 mult1 ( .in_a({a_r[11:2], n7, a_r[0]}), 
        .in_b({b_r[11:10], n5, b_r[8:0]}), .clk(clk), .\output (mult1_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_14 mult2 ( .in_a({a_i[11:2], n6, a_i[0]}), 
        .in_b(b_i), .clk(clk), .\output (mult2_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_13 mult3 ( .in_a({a_r[11:2], n7, a_r[0]}), 
        .in_b(b_i), .clk(clk), .\output (mult3_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_12 mult4 ( .in_a({a_i[11:2], n6, a_i[0]}), 
        .in_b({b_r[11:10], n5, b_r[8:0]}), .clk(clk), .\output (mult4_out) );
  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_3 sub ( .a(mult1_out), .b(mult2_out), .\output ({pre_out_r, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_3 add ( .a(mult3_out), .b(mult4_out), .\output ({pre_out_i, SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_DW01_inc_0 add_154_round ( .A(
        pre_out_i[19:7]), .SUM({rnd_out_i, SYNOPSYS_UNCONNECTED__14}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3_DW01_inc_1 add_140_round ( .A(
        pre_out_r[19:7]), .SUM({rnd_out_r, SYNOPSYS_UNCONNECTED__15}) );
  INVX0 U3 ( .INP(pre_out_r[23]), .ZN(n30) );
  INVX0 U4 ( .INP(pre_out_i[23]), .ZN(n15) );
  INVX0 U5 ( .INP(n31), .ZN(n33) );
  INVX0 U6 ( .INP(n16), .ZN(n18) );
  AND2X1 U7 ( .IN1(n17), .IN2(n19), .Q(n1) );
  AND2X1 U8 ( .IN1(n32), .IN2(n34), .Q(n2) );
  AND2X1 U9 ( .IN1(n18), .IN2(n19), .Q(n3) );
  AND2X1 U10 ( .IN1(n33), .IN2(n34), .Q(n4) );
  NOR2X0 U11 ( .IN1(pre_out_r[21]), .IN2(pre_out_r[22]), .QN(n23) );
  NOR2X0 U12 ( .IN1(pre_out_i[21]), .IN2(pre_out_i[22]), .QN(n8) );
  NAND2X0 U13 ( .IN1(n24), .IN2(n23), .QN(n26) );
  NOR2X0 U14 ( .IN1(pre_out_r[19]), .IN2(pre_out_r[20]), .QN(n24) );
  NAND2X0 U15 ( .IN1(n9), .IN2(n8), .QN(n11) );
  NOR2X0 U16 ( .IN1(pre_out_i[19]), .IN2(pre_out_i[20]), .QN(n9) );
  INVX0 U17 ( .INP(n21), .ZN(n14) );
  INVX0 U18 ( .INP(n19), .ZN(n20) );
  INVX0 U19 ( .INP(n34), .ZN(n35) );
  INVX0 U20 ( .INP(n36), .ZN(n29) );
  DELLN1X2 U21 ( .INP(b_r[9]), .Z(n5) );
  XNOR2X1 U22 ( .IN1(mult3_out[23]), .IN2(mult4_out[23]), .Q(n13) );
  NAND2X0 U23 ( .IN1(n28), .IN2(n27), .QN(n36) );
  DELLN1X2 U24 ( .INP(a_i[1]), .Z(n6) );
  DELLN1X2 U25 ( .INP(a_r[1]), .Z(n7) );
  NAND4X0 U26 ( .IN1(pre_out_i[22]), .IN2(pre_out_i[21]), .IN3(pre_out_i[20]), 
        .IN4(pre_out_i[19]), .QN(n10) );
  MUX21X1 U27 ( .IN1(n11), .IN2(n10), .S(pre_out_i[23]), .Q(n16) );
  XOR2X1 U28 ( .IN1(pre_out_i[23]), .IN2(mult3_out[23]), .Q(n12) );
  NAND2X1 U29 ( .IN1(n13), .IN2(n12), .QN(n21) );
  NAND2X1 U30 ( .IN1(mult3_out[23]), .IN2(n14), .QN(n19) );
  AO21X1 U31 ( .IN1(n16), .IN2(n15), .IN3(n14), .Q(n17) );
  AO21X1 U32 ( .IN1(rnd_out_i[0]), .IN2(n3), .IN3(n1), .Q(pos_out_i[0]) );
  AO21X1 U33 ( .IN1(rnd_out_i[1]), .IN2(n3), .IN3(n1), .Q(pos_out_i[1]) );
  AO21X1 U34 ( .IN1(rnd_out_i[2]), .IN2(n3), .IN3(n1), .Q(pos_out_i[2]) );
  AO21X1 U35 ( .IN1(rnd_out_i[3]), .IN2(n3), .IN3(n1), .Q(pos_out_i[3]) );
  AO21X1 U36 ( .IN1(rnd_out_i[4]), .IN2(n3), .IN3(n1), .Q(pos_out_i[4]) );
  AO21X1 U37 ( .IN1(rnd_out_i[5]), .IN2(n3), .IN3(n1), .Q(pos_out_i[5]) );
  AO21X1 U38 ( .IN1(rnd_out_i[6]), .IN2(n3), .IN3(n1), .Q(pos_out_i[6]) );
  AO21X1 U39 ( .IN1(rnd_out_i[7]), .IN2(n3), .IN3(n1), .Q(pos_out_i[7]) );
  AO21X1 U40 ( .IN1(rnd_out_i[8]), .IN2(n3), .IN3(n1), .Q(pos_out_i[8]) );
  AO21X1 U41 ( .IN1(rnd_out_i[9]), .IN2(n3), .IN3(n1), .Q(pos_out_i[9]) );
  AO21X1 U42 ( .IN1(rnd_out_i[10]), .IN2(n3), .IN3(n1), .Q(pos_out_i[10]) );
  MUX21X1 U43 ( .IN1(pre_out_i[23]), .IN2(rnd_out_i[11]), .S(n18), .Q(n22) );
  AO21X1 U44 ( .IN1(n22), .IN2(n21), .IN3(n20), .Q(pos_out_i[11]) );
  NAND4X0 U45 ( .IN1(pre_out_r[22]), .IN2(pre_out_r[21]), .IN3(pre_out_r[20]), 
        .IN4(pre_out_r[19]), .QN(n25) );
  MUX21X1 U46 ( .IN1(n26), .IN2(n25), .S(pre_out_r[23]), .Q(n31) );
  XOR2X1 U47 ( .IN1(mult2_out[23]), .IN2(mult1_out[23]), .Q(n28) );
  XOR2X1 U48 ( .IN1(pre_out_r[23]), .IN2(mult1_out[23]), .Q(n27) );
  NAND2X1 U49 ( .IN1(mult1_out[23]), .IN2(n29), .QN(n34) );
  AO21X1 U50 ( .IN1(n31), .IN2(n30), .IN3(n29), .Q(n32) );
  AO21X1 U51 ( .IN1(rnd_out_r[0]), .IN2(n4), .IN3(n2), .Q(pos_out_r[0]) );
  AO21X1 U52 ( .IN1(rnd_out_r[1]), .IN2(n4), .IN3(n2), .Q(pos_out_r[1]) );
  AO21X1 U53 ( .IN1(rnd_out_r[2]), .IN2(n4), .IN3(n2), .Q(pos_out_r[2]) );
  AO21X1 U54 ( .IN1(rnd_out_r[3]), .IN2(n4), .IN3(n2), .Q(pos_out_r[3]) );
  AO21X1 U55 ( .IN1(rnd_out_r[4]), .IN2(n4), .IN3(n2), .Q(pos_out_r[4]) );
  AO21X1 U56 ( .IN1(rnd_out_r[5]), .IN2(n4), .IN3(n2), .Q(pos_out_r[5]) );
  AO21X1 U57 ( .IN1(rnd_out_r[6]), .IN2(n4), .IN3(n2), .Q(pos_out_r[6]) );
  AO21X1 U58 ( .IN1(rnd_out_r[7]), .IN2(n4), .IN3(n2), .Q(pos_out_r[7]) );
  AO21X1 U59 ( .IN1(rnd_out_r[8]), .IN2(n4), .IN3(n2), .Q(pos_out_r[8]) );
  AO21X1 U60 ( .IN1(rnd_out_r[9]), .IN2(n4), .IN3(n2), .Q(pos_out_r[9]) );
  AO21X1 U61 ( .IN1(rnd_out_r[10]), .IN2(n4), .IN3(n2), .Q(pos_out_r[10]) );
  MUX21X1 U62 ( .IN1(pre_out_r[23]), .IN2(rnd_out_r[11]), .S(n33), .Q(n37) );
  AO21X1 U63 ( .IN1(n37), .IN2(n36), .IN3(n35), .Q(pos_out_r[11]) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_11_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n450), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n452), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n454), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n456), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  DELLN1X2 U311 ( .INP(b[4]), .Z(n408) );
  FADDX1 U312 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  XOR2X1 U313 ( .IN1(b[2]), .IN2(n431), .Q(n479) );
  FADDX1 U314 ( .A(n27), .B(n448), .CI(n5), .CO(n4), .S(product[21]) );
  DELLN1X2 U315 ( .INP(b[3]), .Z(n409) );
  INVX0 U316 ( .INP(n435), .ZN(n410) );
  INVX0 U317 ( .INP(n435), .ZN(n411) );
  XOR2X2 U318 ( .IN1(n432), .IN2(n446), .Q(n533) );
  XOR2X2 U319 ( .IN1(n432), .IN2(n444), .Q(n522) );
  XOR2X2 U320 ( .IN1(n411), .IN2(n442), .Q(n511) );
  XOR2X2 U321 ( .IN1(n411), .IN2(n440), .Q(n500) );
  XOR2X2 U322 ( .IN1(n432), .IN2(n438), .Q(n490) );
  XOR2X2 U323 ( .IN1(b[2]), .IN2(n446), .Q(n534) );
  XOR2X2 U324 ( .IN1(b[2]), .IN2(n444), .Q(n523) );
  XOR2X2 U325 ( .IN1(b[2]), .IN2(n442), .Q(n512) );
  XOR2X2 U326 ( .IN1(b[2]), .IN2(n440), .Q(n501) );
  XOR2X2 U327 ( .IN1(b[2]), .IN2(n438), .Q(n491) );
  XOR2X2 U328 ( .IN1(b[10]), .IN2(n446), .Q(n477) );
  XOR2X2 U329 ( .IN1(b[10]), .IN2(n444), .Q(n474) );
  XOR2X2 U330 ( .IN1(b[10]), .IN2(n442), .Q(n471) );
  XOR2X2 U331 ( .IN1(b[10]), .IN2(n440), .Q(n468) );
  XOR2X2 U332 ( .IN1(b[10]), .IN2(n438), .Q(n460) );
  XOR3X2 U333 ( .IN1(n57), .IN2(n50), .IN3(n11), .Q(product[15]) );
  NAND2X0 U334 ( .IN1(n57), .IN2(n50), .QN(n412) );
  NAND2X0 U335 ( .IN1(n57), .IN2(n11), .QN(n413) );
  NAND2X0 U336 ( .IN1(n50), .IN2(n11), .QN(n414) );
  NAND3X0 U337 ( .IN1(n412), .IN2(n413), .IN3(n414), .QN(n10) );
  XOR2X1 U338 ( .IN1(n49), .IN2(n44), .Q(n415) );
  XOR2X1 U339 ( .IN1(n415), .IN2(n10), .Q(product[16]) );
  NAND2X0 U340 ( .IN1(n49), .IN2(n44), .QN(n416) );
  NAND2X0 U341 ( .IN1(n49), .IN2(n10), .QN(n417) );
  NAND2X0 U342 ( .IN1(n44), .IN2(n10), .QN(n418) );
  NAND3X0 U343 ( .IN1(n416), .IN2(n417), .IN3(n418), .QN(n9) );
  XOR2X2 U344 ( .IN1(b[9]), .IN2(n446), .Q(n541) );
  XOR2X2 U345 ( .IN1(b[9]), .IN2(n444), .Q(n530) );
  XOR2X2 U346 ( .IN1(b[9]), .IN2(n442), .Q(n519) );
  XOR2X2 U347 ( .IN1(b[9]), .IN2(n440), .Q(n508) );
  XOR2X2 U348 ( .IN1(b[9]), .IN2(n438), .Q(n462) );
  XOR2X2 U349 ( .IN1(b[9]), .IN2(n431), .Q(n486) );
  AO22X1 U350 ( .IN1(n436), .IN2(n484), .IN3(n463), .IN4(n483), .Q(n218) );
  XOR2X2 U351 ( .IN1(b[8]), .IN2(n446), .Q(n540) );
  XOR2X2 U352 ( .IN1(b[8]), .IN2(n444), .Q(n529) );
  XOR2X2 U353 ( .IN1(b[8]), .IN2(n442), .Q(n518) );
  XOR2X2 U354 ( .IN1(b[8]), .IN2(n440), .Q(n507) );
  XOR2X2 U355 ( .IN1(b[8]), .IN2(n438), .Q(n497) );
  XOR2X2 U356 ( .IN1(b[8]), .IN2(n431), .Q(n485) );
  XOR2X2 U357 ( .IN1(b[6]), .IN2(n446), .Q(n538) );
  XOR2X2 U358 ( .IN1(b[6]), .IN2(n444), .Q(n527) );
  XOR2X2 U359 ( .IN1(b[6]), .IN2(n442), .Q(n516) );
  XOR2X2 U360 ( .IN1(b[6]), .IN2(n440), .Q(n505) );
  XOR2X2 U361 ( .IN1(b[6]), .IN2(n438), .Q(n495) );
  XOR2X2 U362 ( .IN1(b[6]), .IN2(n431), .Q(n483) );
  XOR2X2 U363 ( .IN1(b[10]), .IN2(n431), .Q(n487) );
  XOR2X2 U364 ( .IN1(b[1]), .IN2(n446), .Q(n532) );
  XOR2X2 U365 ( .IN1(b[1]), .IN2(n444), .Q(n521) );
  XOR2X2 U366 ( .IN1(b[1]), .IN2(n442), .Q(n510) );
  XOR2X2 U367 ( .IN1(b[1]), .IN2(n440), .Q(n499) );
  XOR2X2 U368 ( .IN1(b[1]), .IN2(n438), .Q(n489) );
  XOR2X2 U369 ( .IN1(b[1]), .IN2(n431), .Q(n478) );
  DELLN2X2 U370 ( .INP(b[5]), .Z(n430) );
  FADDX1 U371 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U372 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  XOR3X1 U373 ( .IN1(n76), .IN2(n85), .IN3(n14), .Q(product[12]) );
  XNOR2X1 U374 ( .IN1(n419), .IN2(n13), .Q(product[13]) );
  XNOR2X1 U375 ( .IN1(n66), .IN2(n75), .Q(n419) );
  XNOR2X1 U376 ( .IN1(n420), .IN2(n15), .Q(product[11]) );
  XNOR2X1 U377 ( .IN1(n95), .IN2(n86), .Q(n420) );
  INVX0 U378 ( .INP(n25), .ZN(n448) );
  FADDX1 U379 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U380 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  INVX0 U381 ( .INP(n3), .ZN(product[23]) );
  INVX0 U382 ( .INP(n55), .ZN(n454) );
  FADDX1 U383 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U384 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X1 U385 ( .IN1(n408), .IN2(n431), .Q(n481) );
  XOR2X1 U386 ( .IN1(n409), .IN2(n431), .Q(n480) );
  XOR2X1 U387 ( .IN1(n409), .IN2(n438), .Q(n492) );
  XOR2X1 U388 ( .IN1(n409), .IN2(n440), .Q(n502) );
  INVX0 U389 ( .INP(n73), .ZN(n456) );
  XOR2X1 U390 ( .IN1(n409), .IN2(n442), .Q(n513) );
  XOR2X1 U391 ( .IN1(n409), .IN2(n444), .Q(n524) );
  XOR2X1 U392 ( .IN1(n409), .IN2(n446), .Q(n535) );
  INVX0 U393 ( .INP(n31), .ZN(n450) );
  INVX0 U394 ( .INP(n41), .ZN(n452) );
  NBUFFX2 U395 ( .INP(a[1]), .Z(n431) );
  INVX0 U396 ( .INP(n488), .ZN(n457) );
  AND2X1 U397 ( .IN1(n431), .IN2(n437), .Q(n463) );
  INVX0 U398 ( .INP(n498), .ZN(n455) );
  INVX0 U399 ( .INP(n509), .ZN(n453) );
  INVX0 U400 ( .INP(n520), .ZN(n451) );
  INVX0 U401 ( .INP(n531), .ZN(n449) );
  NBUFFX2 U402 ( .INP(a[3]), .Z(n439) );
  NBUFFX2 U403 ( .INP(a[5]), .Z(n441) );
  AND2X1 U404 ( .IN1(n488), .IN2(n543), .Q(n461) );
  AND2X1 U405 ( .IN1(n509), .IN2(n547), .Q(n470) );
  AND2X1 U406 ( .IN1(n498), .IN2(n545), .Q(n467) );
  AND2X1 U407 ( .IN1(n520), .IN2(n549), .Q(n473) );
  AND2X1 U408 ( .IN1(n531), .IN2(n551), .Q(n476) );
  NBUFFX2 U409 ( .INP(a[7]), .Z(n443) );
  NBUFFX2 U410 ( .INP(a[9]), .Z(n445) );
  NAND2X0 U411 ( .IN1(n76), .IN2(n85), .QN(n421) );
  NAND2X0 U412 ( .IN1(n76), .IN2(n14), .QN(n422) );
  NAND2X0 U413 ( .IN1(n85), .IN2(n14), .QN(n423) );
  NAND3X0 U414 ( .IN1(n423), .IN2(n422), .IN3(n421), .QN(n13) );
  NAND2X0 U415 ( .IN1(n66), .IN2(n75), .QN(n424) );
  NAND2X0 U416 ( .IN1(n66), .IN2(n13), .QN(n425) );
  NAND2X0 U417 ( .IN1(n75), .IN2(n13), .QN(n426) );
  NAND3X0 U418 ( .IN1(n424), .IN2(n425), .IN3(n426), .QN(n12) );
  NAND2X0 U419 ( .IN1(n86), .IN2(n15), .QN(n427) );
  NAND2X0 U420 ( .IN1(n95), .IN2(n15), .QN(n428) );
  NAND2X0 U421 ( .IN1(n95), .IN2(n86), .QN(n429) );
  NAND3X0 U422 ( .IN1(n427), .IN2(n428), .IN3(n429), .QN(n14) );
  DELLN1X2 U423 ( .INP(a[11]), .Z(n446) );
  INVX0 U424 ( .INP(n435), .ZN(n432) );
  INVX0 U425 ( .INP(b[0]), .ZN(n433) );
  INVX0 U426 ( .INP(b[0]), .ZN(n434) );
  INVX0 U427 ( .INP(b[0]), .ZN(n435) );
  INVX0 U428 ( .INP(n437), .ZN(n436) );
  INVX0 U429 ( .INP(a[0]), .ZN(n437) );
  DELLN1X2 U430 ( .INP(a[3]), .Z(n438) );
  DELLN1X2 U431 ( .INP(a[5]), .Z(n440) );
  DELLN1X2 U432 ( .INP(a[7]), .Z(n442) );
  DELLN1X2 U433 ( .INP(a[9]), .Z(n444) );
  NOR2X0 U434 ( .IN1(n437), .IN2(n434), .QN(product[0]) );
  XNOR2X1 U435 ( .IN1(n458), .IN2(n459), .Q(n84) );
  NAND2X0 U436 ( .IN1(n459), .IN2(n458), .QN(n83) );
  AOI22X1 U437 ( .IN1(n460), .IN2(n457), .IN3(n461), .IN4(n462), .QN(n458) );
  OA21X1 U438 ( .IN1(n463), .IN2(n436), .IN3(n464), .Q(n459) );
  AO22X1 U439 ( .IN1(n465), .IN2(n457), .IN3(n461), .IN4(n460), .Q(n73) );
  AO22X1 U440 ( .IN1(n466), .IN2(n455), .IN3(n467), .IN4(n468), .Q(n55) );
  AO22X1 U441 ( .IN1(n469), .IN2(n453), .IN3(n470), .IN4(n471), .Q(n41) );
  AO22X1 U442 ( .IN1(n472), .IN2(n451), .IN3(n473), .IN4(n474), .Q(n31) );
  AO22X1 U443 ( .IN1(n475), .IN2(n449), .IN3(n476), .IN4(n477), .Q(n25) );
  AO22X1 U444 ( .IN1(n436), .IN2(n478), .IN3(n463), .IN4(n435), .Q(n224) );
  AO22X1 U445 ( .IN1(n436), .IN2(n479), .IN3(n463), .IN4(n478), .Q(n223) );
  AO22X1 U446 ( .IN1(n436), .IN2(n480), .IN3(n463), .IN4(n479), .Q(n222) );
  AO22X1 U447 ( .IN1(n436), .IN2(n481), .IN3(n463), .IN4(n480), .Q(n221) );
  AO22X1 U448 ( .IN1(n436), .IN2(n482), .IN3(n463), .IN4(n481), .Q(n220) );
  AO22X1 U449 ( .IN1(n436), .IN2(n483), .IN3(n463), .IN4(n482), .Q(n219) );
  XOR2X1 U450 ( .IN1(n430), .IN2(n431), .Q(n482) );
  AO22X1 U451 ( .IN1(n436), .IN2(n485), .IN3(n463), .IN4(n484), .Q(n217) );
  XOR2X1 U452 ( .IN1(b[7]), .IN2(n431), .Q(n484) );
  AO22X1 U453 ( .IN1(n436), .IN2(n486), .IN3(n463), .IN4(n485), .Q(n216) );
  AO22X1 U454 ( .IN1(n436), .IN2(n487), .IN3(n463), .IN4(n486), .Q(n215) );
  AO22X1 U455 ( .IN1(n436), .IN2(n464), .IN3(n463), .IN4(n487), .Q(n214) );
  XOR2X1 U456 ( .IN1(b[11]), .IN2(n431), .Q(n464) );
  NOR2X0 U457 ( .IN1(n488), .IN2(n434), .QN(n212) );
  AO22X1 U458 ( .IN1(n489), .IN2(n457), .IN3(n461), .IN4(n490), .Q(n211) );
  AO22X1 U459 ( .IN1(n491), .IN2(n457), .IN3(n461), .IN4(n489), .Q(n210) );
  AO22X1 U460 ( .IN1(n492), .IN2(n457), .IN3(n461), .IN4(n491), .Q(n209) );
  AO22X1 U461 ( .IN1(n493), .IN2(n457), .IN3(n461), .IN4(n492), .Q(n208) );
  AO22X1 U462 ( .IN1(n494), .IN2(n457), .IN3(n461), .IN4(n493), .Q(n207) );
  XOR2X1 U463 ( .IN1(n408), .IN2(n438), .Q(n493) );
  AO22X1 U464 ( .IN1(n495), .IN2(n457), .IN3(n461), .IN4(n494), .Q(n206) );
  XOR2X1 U465 ( .IN1(n430), .IN2(n438), .Q(n494) );
  AO22X1 U466 ( .IN1(n496), .IN2(n457), .IN3(n461), .IN4(n495), .Q(n205) );
  AO22X1 U467 ( .IN1(n497), .IN2(n457), .IN3(n461), .IN4(n496), .Q(n204) );
  XOR2X1 U468 ( .IN1(b[7]), .IN2(n438), .Q(n496) );
  AO22X1 U469 ( .IN1(n462), .IN2(n457), .IN3(n461), .IN4(n497), .Q(n203) );
  OAI21X1 U470 ( .IN1(n457), .IN2(n461), .IN3(n465), .QN(n201) );
  XOR2X1 U471 ( .IN1(b[11]), .IN2(n438), .Q(n465) );
  NOR2X0 U472 ( .IN1(n498), .IN2(n434), .QN(n200) );
  AO22X1 U473 ( .IN1(n499), .IN2(n455), .IN3(n467), .IN4(n500), .Q(n199) );
  AO22X1 U474 ( .IN1(n501), .IN2(n455), .IN3(n467), .IN4(n499), .Q(n198) );
  AO22X1 U475 ( .IN1(n502), .IN2(n455), .IN3(n467), .IN4(n501), .Q(n197) );
  AO22X1 U476 ( .IN1(n503), .IN2(n455), .IN3(n467), .IN4(n502), .Q(n196) );
  AO22X1 U477 ( .IN1(n504), .IN2(n455), .IN3(n467), .IN4(n503), .Q(n195) );
  XOR2X1 U478 ( .IN1(n408), .IN2(n440), .Q(n503) );
  AO22X1 U479 ( .IN1(n505), .IN2(n455), .IN3(n467), .IN4(n504), .Q(n194) );
  XOR2X1 U480 ( .IN1(n430), .IN2(n440), .Q(n504) );
  AO22X1 U481 ( .IN1(n506), .IN2(n455), .IN3(n467), .IN4(n505), .Q(n193) );
  AO22X1 U482 ( .IN1(n507), .IN2(n455), .IN3(n467), .IN4(n506), .Q(n192) );
  XOR2X1 U483 ( .IN1(b[7]), .IN2(n440), .Q(n506) );
  AO22X1 U484 ( .IN1(n508), .IN2(n455), .IN3(n467), .IN4(n507), .Q(n191) );
  AO22X1 U485 ( .IN1(n468), .IN2(n455), .IN3(n467), .IN4(n508), .Q(n190) );
  OAI21X1 U486 ( .IN1(n455), .IN2(n467), .IN3(n466), .QN(n189) );
  XOR2X1 U487 ( .IN1(b[11]), .IN2(n440), .Q(n466) );
  NOR2X0 U488 ( .IN1(n509), .IN2(n433), .QN(n188) );
  AO22X1 U489 ( .IN1(n510), .IN2(n453), .IN3(n470), .IN4(n511), .Q(n187) );
  AO22X1 U490 ( .IN1(n512), .IN2(n453), .IN3(n470), .IN4(n510), .Q(n186) );
  AO22X1 U491 ( .IN1(n513), .IN2(n453), .IN3(n470), .IN4(n512), .Q(n185) );
  AO22X1 U492 ( .IN1(n514), .IN2(n453), .IN3(n470), .IN4(n513), .Q(n184) );
  AO22X1 U493 ( .IN1(n515), .IN2(n453), .IN3(n470), .IN4(n514), .Q(n183) );
  XOR2X1 U494 ( .IN1(n408), .IN2(n442), .Q(n514) );
  AO22X1 U495 ( .IN1(n516), .IN2(n453), .IN3(n470), .IN4(n515), .Q(n182) );
  XOR2X1 U496 ( .IN1(n430), .IN2(n442), .Q(n515) );
  AO22X1 U497 ( .IN1(n517), .IN2(n453), .IN3(n470), .IN4(n516), .Q(n181) );
  AO22X1 U498 ( .IN1(n518), .IN2(n453), .IN3(n470), .IN4(n517), .Q(n180) );
  XOR2X1 U499 ( .IN1(b[7]), .IN2(n442), .Q(n517) );
  AO22X1 U500 ( .IN1(n519), .IN2(n453), .IN3(n470), .IN4(n518), .Q(n179) );
  AO22X1 U501 ( .IN1(n471), .IN2(n453), .IN3(n470), .IN4(n519), .Q(n178) );
  OAI21X1 U502 ( .IN1(n453), .IN2(n470), .IN3(n469), .QN(n177) );
  XOR2X1 U503 ( .IN1(b[11]), .IN2(n442), .Q(n469) );
  NOR2X0 U504 ( .IN1(n520), .IN2(n433), .QN(n176) );
  AO22X1 U505 ( .IN1(n521), .IN2(n451), .IN3(n473), .IN4(n522), .Q(n175) );
  AO22X1 U506 ( .IN1(n523), .IN2(n451), .IN3(n473), .IN4(n521), .Q(n174) );
  AO22X1 U507 ( .IN1(n524), .IN2(n451), .IN3(n473), .IN4(n523), .Q(n173) );
  AO22X1 U508 ( .IN1(n525), .IN2(n451), .IN3(n473), .IN4(n524), .Q(n172) );
  AO22X1 U509 ( .IN1(n526), .IN2(n451), .IN3(n473), .IN4(n525), .Q(n171) );
  XOR2X1 U510 ( .IN1(n408), .IN2(n444), .Q(n525) );
  AO22X1 U511 ( .IN1(n527), .IN2(n451), .IN3(n473), .IN4(n526), .Q(n170) );
  XOR2X1 U512 ( .IN1(n430), .IN2(n444), .Q(n526) );
  AO22X1 U513 ( .IN1(n528), .IN2(n451), .IN3(n473), .IN4(n527), .Q(n169) );
  AO22X1 U514 ( .IN1(n529), .IN2(n451), .IN3(n473), .IN4(n528), .Q(n168) );
  XOR2X1 U515 ( .IN1(b[7]), .IN2(n444), .Q(n528) );
  AO22X1 U516 ( .IN1(n530), .IN2(n451), .IN3(n473), .IN4(n529), .Q(n167) );
  AO22X1 U517 ( .IN1(n474), .IN2(n451), .IN3(n473), .IN4(n530), .Q(n166) );
  OAI21X1 U518 ( .IN1(n451), .IN2(n473), .IN3(n472), .QN(n165) );
  XOR2X1 U519 ( .IN1(b[11]), .IN2(n444), .Q(n472) );
  NOR2X0 U520 ( .IN1(n531), .IN2(n433), .QN(n164) );
  AO22X1 U521 ( .IN1(n532), .IN2(n449), .IN3(n476), .IN4(n533), .Q(n163) );
  AO22X1 U522 ( .IN1(n534), .IN2(n449), .IN3(n476), .IN4(n532), .Q(n162) );
  AO22X1 U523 ( .IN1(n535), .IN2(n449), .IN3(n476), .IN4(n534), .Q(n161) );
  AO22X1 U524 ( .IN1(n536), .IN2(n449), .IN3(n476), .IN4(n535), .Q(n160) );
  AO22X1 U525 ( .IN1(n537), .IN2(n449), .IN3(n476), .IN4(n536), .Q(n159) );
  XOR2X1 U526 ( .IN1(n408), .IN2(n446), .Q(n536) );
  AO22X1 U527 ( .IN1(n538), .IN2(n449), .IN3(n476), .IN4(n537), .Q(n158) );
  XOR2X1 U528 ( .IN1(n430), .IN2(n446), .Q(n537) );
  AO22X1 U529 ( .IN1(n539), .IN2(n449), .IN3(n476), .IN4(n538), .Q(n157) );
  AO22X1 U530 ( .IN1(n540), .IN2(n449), .IN3(n476), .IN4(n539), .Q(n156) );
  XOR2X1 U531 ( .IN1(b[7]), .IN2(n446), .Q(n539) );
  AO22X1 U532 ( .IN1(n541), .IN2(n449), .IN3(n476), .IN4(n540), .Q(n155) );
  AO22X1 U533 ( .IN1(n477), .IN2(n449), .IN3(n476), .IN4(n541), .Q(n154) );
  OAI21X1 U534 ( .IN1(n449), .IN2(n476), .IN3(n475), .QN(n153) );
  XOR2X1 U535 ( .IN1(b[11]), .IN2(n446), .Q(n475) );
  AO21X1 U536 ( .IN1(n431), .IN2(n435), .IN3(n463), .Q(n152) );
  AO22X1 U537 ( .IN1(n542), .IN2(n439), .IN3(n461), .IN4(n439), .Q(n151) );
  XOR2X1 U538 ( .IN1(n438), .IN2(a[2]), .Q(n543) );
  NOR2X0 U539 ( .IN1(n410), .IN2(n488), .QN(n542) );
  XNOR2X1 U540 ( .IN1(a[2]), .IN2(n431), .Q(n488) );
  AO22X1 U541 ( .IN1(n544), .IN2(n441), .IN3(n467), .IN4(n441), .Q(n150) );
  XOR2X1 U542 ( .IN1(n440), .IN2(a[4]), .Q(n545) );
  NOR2X0 U543 ( .IN1(n432), .IN2(n498), .QN(n544) );
  XNOR2X1 U544 ( .IN1(a[4]), .IN2(n438), .Q(n498) );
  AO22X1 U545 ( .IN1(n546), .IN2(n443), .IN3(n470), .IN4(n443), .Q(n149) );
  XOR2X1 U546 ( .IN1(n442), .IN2(a[6]), .Q(n547) );
  NOR2X0 U547 ( .IN1(n410), .IN2(n509), .QN(n546) );
  XNOR2X1 U548 ( .IN1(a[6]), .IN2(n440), .Q(n509) );
  AO22X1 U549 ( .IN1(n548), .IN2(n445), .IN3(n473), .IN4(n445), .Q(n148) );
  XOR2X1 U550 ( .IN1(n444), .IN2(a[8]), .Q(n549) );
  NOR2X0 U551 ( .IN1(n410), .IN2(n520), .QN(n548) );
  XNOR2X1 U552 ( .IN1(a[8]), .IN2(n442), .Q(n520) );
  AO22X1 U553 ( .IN1(n550), .IN2(n446), .IN3(n476), .IN4(n446), .Q(n147) );
  XOR2X1 U554 ( .IN1(n446), .IN2(a[10]), .Q(n551) );
  NOR2X0 U555 ( .IN1(n411), .IN2(n531), .QN(n550) );
  XNOR2X1 U556 ( .IN1(a[10]), .IN2(n444), .Q(n531) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_11 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_11_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_10_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567;

  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n466), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n468), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n470), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n472), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(b[5]), .ZN(n408) );
  INVX0 U312 ( .INP(n408), .ZN(n409) );
  XOR2X2 U313 ( .IN1(b[10]), .IN2(n463), .Q(n493) );
  XOR2X2 U314 ( .IN1(b[10]), .IN2(n461), .Q(n490) );
  XOR2X2 U315 ( .IN1(b[10]), .IN2(n459), .Q(n487) );
  XOR2X2 U316 ( .IN1(b[10]), .IN2(n457), .Q(n484) );
  XOR2X2 U317 ( .IN1(b[10]), .IN2(n455), .Q(n476) );
  XOR2X2 U318 ( .IN1(b[10]), .IN2(n450), .Q(n503) );
  XOR2X2 U319 ( .IN1(b[2]), .IN2(n463), .Q(n550) );
  XOR2X2 U320 ( .IN1(b[2]), .IN2(n461), .Q(n539) );
  XOR2X2 U321 ( .IN1(b[2]), .IN2(n459), .Q(n528) );
  XOR2X2 U322 ( .IN1(b[2]), .IN2(n457), .Q(n517) );
  XOR2X2 U323 ( .IN1(b[2]), .IN2(n455), .Q(n507) );
  XOR2X2 U324 ( .IN1(b[2]), .IN2(n450), .Q(n495) );
  XOR3X1 U325 ( .IN1(n105), .IN2(n100), .IN3(n98), .Q(n96) );
  XOR2X1 U326 ( .IN1(n103), .IN2(n16), .Q(n410) );
  XOR2X2 U327 ( .IN1(n410), .IN2(n96), .Q(product[10]) );
  NAND2X0 U328 ( .IN1(n105), .IN2(n100), .QN(n411) );
  NAND2X0 U329 ( .IN1(n105), .IN2(n98), .QN(n412) );
  NAND2X0 U330 ( .IN1(n100), .IN2(n98), .QN(n413) );
  NAND3X0 U331 ( .IN1(n411), .IN2(n412), .IN3(n413), .QN(n95) );
  NAND2X0 U332 ( .IN1(n103), .IN2(n16), .QN(n414) );
  NAND2X0 U333 ( .IN1(n103), .IN2(n96), .QN(n415) );
  NAND2X0 U334 ( .IN1(n16), .IN2(n96), .QN(n416) );
  NAND3X0 U335 ( .IN1(n414), .IN2(n415), .IN3(n416), .QN(n15) );
  XOR3X1 U336 ( .IN1(n215), .IN2(n164), .IN3(n204), .Q(n102) );
  XOR2X1 U337 ( .IN1(n109), .IN2(n107), .Q(n417) );
  XOR2X1 U338 ( .IN1(n417), .IN2(n102), .Q(n98) );
  NAND2X0 U339 ( .IN1(n215), .IN2(n164), .QN(n418) );
  NAND2X0 U340 ( .IN1(n215), .IN2(n204), .QN(n419) );
  NAND2X1 U341 ( .IN1(n164), .IN2(n204), .QN(n420) );
  NAND3X0 U342 ( .IN1(n418), .IN2(n419), .IN3(n420), .QN(n101) );
  NAND2X1 U343 ( .IN1(n109), .IN2(n107), .QN(n421) );
  NAND2X0 U344 ( .IN1(n109), .IN2(n102), .QN(n422) );
  NAND2X0 U345 ( .IN1(n107), .IN2(n102), .QN(n423) );
  NAND3X0 U346 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n97) );
  XOR3X2 U347 ( .IN1(n27), .IN2(n464), .IN3(n5), .Q(product[21]) );
  XOR2X2 U348 ( .IN1(b[9]), .IN2(n463), .Q(n557) );
  XOR2X2 U349 ( .IN1(b[9]), .IN2(n461), .Q(n546) );
  XOR2X2 U350 ( .IN1(b[9]), .IN2(n459), .Q(n535) );
  XOR2X2 U351 ( .IN1(b[9]), .IN2(n457), .Q(n524) );
  XOR2X2 U352 ( .IN1(b[9]), .IN2(n455), .Q(n478) );
  XOR2X2 U353 ( .IN1(b[9]), .IN2(n450), .Q(n502) );
  XOR2X2 U354 ( .IN1(b[8]), .IN2(n463), .Q(n556) );
  XOR2X2 U355 ( .IN1(b[8]), .IN2(n461), .Q(n545) );
  XOR2X2 U356 ( .IN1(b[8]), .IN2(n459), .Q(n534) );
  XOR2X2 U357 ( .IN1(b[8]), .IN2(n457), .Q(n523) );
  XOR2X2 U358 ( .IN1(b[8]), .IN2(n455), .Q(n513) );
  XOR2X2 U359 ( .IN1(b[8]), .IN2(n450), .Q(n501) );
  XOR2X2 U360 ( .IN1(b[7]), .IN2(n463), .Q(n555) );
  XOR2X2 U361 ( .IN1(b[7]), .IN2(n461), .Q(n544) );
  XOR2X2 U362 ( .IN1(b[7]), .IN2(n459), .Q(n533) );
  XOR2X2 U363 ( .IN1(b[7]), .IN2(n457), .Q(n522) );
  XOR2X2 U364 ( .IN1(b[7]), .IN2(n455), .Q(n512) );
  XOR2X2 U365 ( .IN1(b[7]), .IN2(n450), .Q(n500) );
  XOR2X2 U366 ( .IN1(b[4]), .IN2(n463), .Q(n552) );
  XOR2X2 U367 ( .IN1(b[4]), .IN2(n461), .Q(n541) );
  XOR2X2 U368 ( .IN1(b[4]), .IN2(n459), .Q(n530) );
  XOR2X2 U369 ( .IN1(b[4]), .IN2(n457), .Q(n519) );
  XOR2X2 U370 ( .IN1(b[4]), .IN2(n455), .Q(n509) );
  XOR2X2 U371 ( .IN1(b[4]), .IN2(n450), .Q(n497) );
  XOR2X2 U372 ( .IN1(b[6]), .IN2(n463), .Q(n554) );
  XOR2X2 U373 ( .IN1(b[6]), .IN2(n461), .Q(n543) );
  XOR2X2 U374 ( .IN1(b[6]), .IN2(n459), .Q(n532) );
  XOR2X2 U375 ( .IN1(b[6]), .IN2(n457), .Q(n521) );
  XOR2X2 U376 ( .IN1(b[6]), .IN2(n455), .Q(n511) );
  XOR2X2 U377 ( .IN1(b[6]), .IN2(n450), .Q(n499) );
  XOR2X2 U378 ( .IN1(b[1]), .IN2(n463), .Q(n548) );
  XOR2X2 U379 ( .IN1(b[1]), .IN2(n461), .Q(n537) );
  XOR2X2 U380 ( .IN1(b[1]), .IN2(n459), .Q(n526) );
  XOR2X2 U381 ( .IN1(b[1]), .IN2(n457), .Q(n515) );
  XOR2X2 U382 ( .IN1(b[1]), .IN2(n455), .Q(n505) );
  XOR2X2 U383 ( .IN1(b[1]), .IN2(n450), .Q(n494) );
  XOR2X2 U384 ( .IN1(n409), .IN2(n463), .Q(n553) );
  XOR2X2 U385 ( .IN1(n409), .IN2(n461), .Q(n542) );
  XOR2X2 U386 ( .IN1(n409), .IN2(n459), .Q(n531) );
  XOR2X2 U387 ( .IN1(n409), .IN2(n457), .Q(n520) );
  XOR2X2 U388 ( .IN1(n409), .IN2(n455), .Q(n510) );
  XOR2X2 U389 ( .IN1(n409), .IN2(n450), .Q(n498) );
  XOR2X1 U390 ( .IN1(n424), .IN2(n4), .Q(product[22]) );
  XOR2X1 U391 ( .IN1(n25), .IN2(n153), .Q(n424) );
  AND3X1 U392 ( .IN1(n437), .IN2(n438), .IN3(n439), .Q(product[23]) );
  INVX0 U393 ( .INP(n55), .ZN(n470) );
  XOR3X1 U394 ( .IN1(n33), .IN2(n30), .IN3(n7), .Q(product[19]) );
  XNOR2X1 U395 ( .IN1(n426), .IN2(n6), .Q(product[20]) );
  XNOR2X1 U396 ( .IN1(n29), .IN2(n28), .Q(n426) );
  INVX0 U397 ( .INP(n25), .ZN(n464) );
  XOR3X1 U398 ( .IN1(n118), .IN2(n123), .IN3(n19), .Q(product[7]) );
  XOR2X1 U399 ( .IN1(b[3]), .IN2(n450), .Q(n496) );
  XOR2X1 U400 ( .IN1(b[3]), .IN2(n455), .Q(n508) );
  INVX0 U401 ( .INP(n73), .ZN(n472) );
  XOR2X1 U402 ( .IN1(b[3]), .IN2(n457), .Q(n518) );
  XOR2X1 U403 ( .IN1(b[3]), .IN2(n459), .Q(n529) );
  XOR2X1 U404 ( .IN1(b[3]), .IN2(n461), .Q(n540) );
  INVX0 U405 ( .INP(n41), .ZN(n468) );
  XOR2X1 U406 ( .IN1(b[3]), .IN2(n463), .Q(n551) );
  INVX0 U407 ( .INP(n31), .ZN(n466) );
  NBUFFX2 U408 ( .INP(a[1]), .Z(n450) );
  INVX0 U409 ( .INP(n504), .ZN(n473) );
  AND2X1 U410 ( .IN1(n450), .IN2(n454), .Q(n479) );
  INVX0 U411 ( .INP(n514), .ZN(n471) );
  INVX0 U412 ( .INP(n525), .ZN(n469) );
  INVX0 U413 ( .INP(n536), .ZN(n467) );
  XNOR2X1 U414 ( .IN1(n427), .IN2(n20), .Q(product[6]) );
  XNOR2X1 U415 ( .IN1(n127), .IN2(n124), .Q(n427) );
  INVX0 U416 ( .INP(n547), .ZN(n465) );
  NBUFFX2 U417 ( .INP(a[3]), .Z(n456) );
  FADDX1 U418 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  NBUFFX2 U419 ( .INP(a[5]), .Z(n458) );
  AND2X1 U420 ( .IN1(n504), .IN2(n559), .Q(n477) );
  AND2X1 U421 ( .IN1(n525), .IN2(n563), .Q(n486) );
  AND2X1 U422 ( .IN1(n514), .IN2(n561), .Q(n483) );
  AND2X1 U423 ( .IN1(n536), .IN2(n565), .Q(n489) );
  AND2X1 U424 ( .IN1(n547), .IN2(n567), .Q(n492) );
  NBUFFX2 U425 ( .INP(a[7]), .Z(n460) );
  NBUFFX2 U426 ( .INP(a[9]), .Z(n462) );
  NAND2X0 U427 ( .IN1(n33), .IN2(n30), .QN(n428) );
  NAND2X0 U428 ( .IN1(n33), .IN2(n7), .QN(n429) );
  NAND2X0 U429 ( .IN1(n30), .IN2(n7), .QN(n430) );
  NAND3X0 U430 ( .IN1(n428), .IN2(n429), .IN3(n430), .QN(n6) );
  NAND2X0 U431 ( .IN1(n29), .IN2(n28), .QN(n431) );
  NAND2X0 U432 ( .IN1(n29), .IN2(n6), .QN(n432) );
  NAND2X0 U433 ( .IN1(n28), .IN2(n6), .QN(n433) );
  NAND3X0 U434 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(n5) );
  NAND2X1 U435 ( .IN1(n27), .IN2(n464), .QN(n434) );
  NAND2X0 U436 ( .IN1(n27), .IN2(n5), .QN(n435) );
  NAND2X0 U437 ( .IN1(n464), .IN2(n5), .QN(n436) );
  NAND3X0 U438 ( .IN1(n434), .IN2(n435), .IN3(n436), .QN(n4) );
  NAND2X0 U439 ( .IN1(n25), .IN2(n153), .QN(n437) );
  NAND2X0 U440 ( .IN1(n25), .IN2(n4), .QN(n438) );
  NAND2X0 U441 ( .IN1(n153), .IN2(n4), .QN(n439) );
  NAND2X0 U442 ( .IN1(n118), .IN2(n123), .QN(n440) );
  NAND2X0 U443 ( .IN1(n118), .IN2(n19), .QN(n441) );
  NAND2X0 U444 ( .IN1(n123), .IN2(n19), .QN(n442) );
  NAND3X0 U445 ( .IN1(n440), .IN2(n441), .IN3(n442), .QN(n18) );
  XOR2X1 U446 ( .IN1(n112), .IN2(n117), .Q(n443) );
  XOR2X1 U447 ( .IN1(n443), .IN2(n18), .Q(product[8]) );
  NAND2X0 U448 ( .IN1(n112), .IN2(n117), .QN(n444) );
  NAND2X0 U449 ( .IN1(n112), .IN2(n18), .QN(n445) );
  NAND2X0 U450 ( .IN1(n117), .IN2(n18), .QN(n446) );
  NAND3X0 U451 ( .IN1(n444), .IN2(n445), .IN3(n446), .QN(n17) );
  NAND2X0 U452 ( .IN1(n124), .IN2(n20), .QN(n447) );
  NAND2X0 U453 ( .IN1(n127), .IN2(n20), .QN(n448) );
  NAND2X0 U454 ( .IN1(n127), .IN2(n124), .QN(n449) );
  NAND3X0 U455 ( .IN1(n447), .IN2(n449), .IN3(n448), .QN(n19) );
  DELLN1X2 U456 ( .INP(a[11]), .Z(n463) );
  INVX0 U457 ( .INP(n452), .ZN(n451) );
  INVX0 U458 ( .INP(b[0]), .ZN(n452) );
  INVX0 U459 ( .INP(n454), .ZN(n453) );
  INVX0 U460 ( .INP(a[0]), .ZN(n454) );
  DELLN1X2 U461 ( .INP(a[3]), .Z(n455) );
  DELLN1X2 U462 ( .INP(a[5]), .Z(n457) );
  DELLN1X2 U463 ( .INP(a[7]), .Z(n459) );
  DELLN1X2 U464 ( .INP(a[9]), .Z(n461) );
  NOR2X0 U465 ( .IN1(n454), .IN2(n452), .QN(product[0]) );
  XNOR2X1 U466 ( .IN1(n474), .IN2(n475), .Q(n84) );
  NAND2X0 U467 ( .IN1(n475), .IN2(n474), .QN(n83) );
  AOI22X1 U468 ( .IN1(n476), .IN2(n473), .IN3(n477), .IN4(n478), .QN(n474) );
  OA21X1 U469 ( .IN1(n479), .IN2(n453), .IN3(n480), .Q(n475) );
  AO22X1 U470 ( .IN1(n481), .IN2(n473), .IN3(n477), .IN4(n476), .Q(n73) );
  AO22X1 U471 ( .IN1(n482), .IN2(n471), .IN3(n483), .IN4(n484), .Q(n55) );
  AO22X1 U472 ( .IN1(n485), .IN2(n469), .IN3(n486), .IN4(n487), .Q(n41) );
  AO22X1 U473 ( .IN1(n488), .IN2(n467), .IN3(n489), .IN4(n490), .Q(n31) );
  AO22X1 U474 ( .IN1(n491), .IN2(n465), .IN3(n492), .IN4(n493), .Q(n25) );
  AO22X1 U475 ( .IN1(n453), .IN2(n494), .IN3(n479), .IN4(n452), .Q(n224) );
  AO22X1 U476 ( .IN1(n453), .IN2(n495), .IN3(n479), .IN4(n494), .Q(n223) );
  AO22X1 U477 ( .IN1(n453), .IN2(n496), .IN3(n479), .IN4(n495), .Q(n222) );
  AO22X1 U478 ( .IN1(n453), .IN2(n497), .IN3(n479), .IN4(n496), .Q(n221) );
  AO22X1 U479 ( .IN1(n453), .IN2(n498), .IN3(n479), .IN4(n497), .Q(n220) );
  AO22X1 U480 ( .IN1(n453), .IN2(n499), .IN3(n479), .IN4(n498), .Q(n219) );
  AO22X1 U481 ( .IN1(n453), .IN2(n500), .IN3(n479), .IN4(n499), .Q(n218) );
  AO22X1 U482 ( .IN1(n453), .IN2(n501), .IN3(n479), .IN4(n500), .Q(n217) );
  AO22X1 U483 ( .IN1(n453), .IN2(n502), .IN3(n479), .IN4(n501), .Q(n216) );
  AO22X1 U484 ( .IN1(n453), .IN2(n503), .IN3(n479), .IN4(n502), .Q(n215) );
  AO22X1 U485 ( .IN1(n453), .IN2(n480), .IN3(n479), .IN4(n503), .Q(n214) );
  XOR2X1 U486 ( .IN1(b[11]), .IN2(n450), .Q(n480) );
  NOR2X0 U487 ( .IN1(n504), .IN2(n452), .QN(n212) );
  AO22X1 U488 ( .IN1(n505), .IN2(n473), .IN3(n477), .IN4(n506), .Q(n211) );
  XOR2X1 U489 ( .IN1(n451), .IN2(n455), .Q(n506) );
  AO22X1 U490 ( .IN1(n507), .IN2(n473), .IN3(n477), .IN4(n505), .Q(n210) );
  AO22X1 U491 ( .IN1(n508), .IN2(n473), .IN3(n477), .IN4(n507), .Q(n209) );
  AO22X1 U492 ( .IN1(n509), .IN2(n473), .IN3(n477), .IN4(n508), .Q(n208) );
  AO22X1 U493 ( .IN1(n510), .IN2(n473), .IN3(n477), .IN4(n509), .Q(n207) );
  AO22X1 U494 ( .IN1(n511), .IN2(n473), .IN3(n477), .IN4(n510), .Q(n206) );
  AO22X1 U495 ( .IN1(n512), .IN2(n473), .IN3(n477), .IN4(n511), .Q(n205) );
  AO22X1 U496 ( .IN1(n513), .IN2(n473), .IN3(n477), .IN4(n512), .Q(n204) );
  AO22X1 U497 ( .IN1(n478), .IN2(n473), .IN3(n477), .IN4(n513), .Q(n203) );
  OAI21X1 U498 ( .IN1(n473), .IN2(n477), .IN3(n481), .QN(n201) );
  XOR2X1 U499 ( .IN1(b[11]), .IN2(n455), .Q(n481) );
  NOR2X0 U500 ( .IN1(n514), .IN2(n452), .QN(n200) );
  AO22X1 U501 ( .IN1(n515), .IN2(n471), .IN3(n483), .IN4(n516), .Q(n199) );
  XOR2X1 U502 ( .IN1(n451), .IN2(n457), .Q(n516) );
  AO22X1 U503 ( .IN1(n517), .IN2(n471), .IN3(n483), .IN4(n515), .Q(n198) );
  AO22X1 U504 ( .IN1(n518), .IN2(n471), .IN3(n483), .IN4(n517), .Q(n197) );
  AO22X1 U505 ( .IN1(n519), .IN2(n471), .IN3(n483), .IN4(n518), .Q(n196) );
  AO22X1 U506 ( .IN1(n520), .IN2(n471), .IN3(n483), .IN4(n519), .Q(n195) );
  AO22X1 U507 ( .IN1(n521), .IN2(n471), .IN3(n483), .IN4(n520), .Q(n194) );
  AO22X1 U508 ( .IN1(n522), .IN2(n471), .IN3(n483), .IN4(n521), .Q(n193) );
  AO22X1 U509 ( .IN1(n523), .IN2(n471), .IN3(n483), .IN4(n522), .Q(n192) );
  AO22X1 U510 ( .IN1(n524), .IN2(n471), .IN3(n483), .IN4(n523), .Q(n191) );
  AO22X1 U511 ( .IN1(n484), .IN2(n471), .IN3(n483), .IN4(n524), .Q(n190) );
  OAI21X1 U512 ( .IN1(n471), .IN2(n483), .IN3(n482), .QN(n189) );
  XOR2X1 U513 ( .IN1(b[11]), .IN2(n457), .Q(n482) );
  NOR2X0 U514 ( .IN1(n525), .IN2(n452), .QN(n188) );
  AO22X1 U515 ( .IN1(n526), .IN2(n469), .IN3(n486), .IN4(n527), .Q(n187) );
  XOR2X1 U516 ( .IN1(n451), .IN2(n459), .Q(n527) );
  AO22X1 U517 ( .IN1(n528), .IN2(n469), .IN3(n486), .IN4(n526), .Q(n186) );
  AO22X1 U518 ( .IN1(n529), .IN2(n469), .IN3(n486), .IN4(n528), .Q(n185) );
  AO22X1 U519 ( .IN1(n530), .IN2(n469), .IN3(n486), .IN4(n529), .Q(n184) );
  AO22X1 U520 ( .IN1(n531), .IN2(n469), .IN3(n486), .IN4(n530), .Q(n183) );
  AO22X1 U521 ( .IN1(n532), .IN2(n469), .IN3(n486), .IN4(n531), .Q(n182) );
  AO22X1 U522 ( .IN1(n533), .IN2(n469), .IN3(n486), .IN4(n532), .Q(n181) );
  AO22X1 U523 ( .IN1(n534), .IN2(n469), .IN3(n486), .IN4(n533), .Q(n180) );
  AO22X1 U524 ( .IN1(n535), .IN2(n469), .IN3(n486), .IN4(n534), .Q(n179) );
  AO22X1 U525 ( .IN1(n487), .IN2(n469), .IN3(n486), .IN4(n535), .Q(n178) );
  OAI21X1 U526 ( .IN1(n469), .IN2(n486), .IN3(n485), .QN(n177) );
  XOR2X1 U527 ( .IN1(b[11]), .IN2(n459), .Q(n485) );
  NOR2X0 U528 ( .IN1(n536), .IN2(n452), .QN(n176) );
  AO22X1 U529 ( .IN1(n537), .IN2(n467), .IN3(n489), .IN4(n538), .Q(n175) );
  XOR2X1 U530 ( .IN1(n451), .IN2(n461), .Q(n538) );
  AO22X1 U531 ( .IN1(n539), .IN2(n467), .IN3(n489), .IN4(n537), .Q(n174) );
  AO22X1 U532 ( .IN1(n540), .IN2(n467), .IN3(n489), .IN4(n539), .Q(n173) );
  AO22X1 U533 ( .IN1(n541), .IN2(n467), .IN3(n489), .IN4(n540), .Q(n172) );
  AO22X1 U534 ( .IN1(n542), .IN2(n467), .IN3(n489), .IN4(n541), .Q(n171) );
  AO22X1 U535 ( .IN1(n543), .IN2(n467), .IN3(n489), .IN4(n542), .Q(n170) );
  AO22X1 U536 ( .IN1(n544), .IN2(n467), .IN3(n489), .IN4(n543), .Q(n169) );
  AO22X1 U537 ( .IN1(n545), .IN2(n467), .IN3(n489), .IN4(n544), .Q(n168) );
  AO22X1 U538 ( .IN1(n546), .IN2(n467), .IN3(n489), .IN4(n545), .Q(n167) );
  AO22X1 U539 ( .IN1(n490), .IN2(n467), .IN3(n489), .IN4(n546), .Q(n166) );
  OAI21X1 U540 ( .IN1(n467), .IN2(n489), .IN3(n488), .QN(n165) );
  XOR2X1 U541 ( .IN1(b[11]), .IN2(n461), .Q(n488) );
  NOR2X0 U542 ( .IN1(n547), .IN2(n452), .QN(n164) );
  AO22X1 U543 ( .IN1(n548), .IN2(n465), .IN3(n492), .IN4(n549), .Q(n163) );
  XOR2X1 U544 ( .IN1(n451), .IN2(n463), .Q(n549) );
  AO22X1 U545 ( .IN1(n550), .IN2(n465), .IN3(n492), .IN4(n548), .Q(n162) );
  AO22X1 U546 ( .IN1(n551), .IN2(n465), .IN3(n492), .IN4(n550), .Q(n161) );
  AO22X1 U547 ( .IN1(n552), .IN2(n465), .IN3(n492), .IN4(n551), .Q(n160) );
  AO22X1 U548 ( .IN1(n553), .IN2(n465), .IN3(n492), .IN4(n552), .Q(n159) );
  AO22X1 U549 ( .IN1(n554), .IN2(n465), .IN3(n492), .IN4(n553), .Q(n158) );
  AO22X1 U550 ( .IN1(n555), .IN2(n465), .IN3(n492), .IN4(n554), .Q(n157) );
  AO22X1 U551 ( .IN1(n556), .IN2(n465), .IN3(n492), .IN4(n555), .Q(n156) );
  AO22X1 U552 ( .IN1(n557), .IN2(n465), .IN3(n492), .IN4(n556), .Q(n155) );
  AO22X1 U553 ( .IN1(n493), .IN2(n465), .IN3(n492), .IN4(n557), .Q(n154) );
  OAI21X1 U554 ( .IN1(n465), .IN2(n492), .IN3(n491), .QN(n153) );
  XOR2X1 U555 ( .IN1(b[11]), .IN2(n463), .Q(n491) );
  AO21X1 U556 ( .IN1(n450), .IN2(n452), .IN3(n479), .Q(n152) );
  AO22X1 U557 ( .IN1(n558), .IN2(n456), .IN3(n477), .IN4(n456), .Q(n151) );
  XOR2X1 U558 ( .IN1(n455), .IN2(a[2]), .Q(n559) );
  NOR2X0 U559 ( .IN1(n451), .IN2(n504), .QN(n558) );
  XNOR2X1 U560 ( .IN1(a[2]), .IN2(n450), .Q(n504) );
  AO22X1 U561 ( .IN1(n560), .IN2(n458), .IN3(n483), .IN4(n458), .Q(n150) );
  XOR2X1 U562 ( .IN1(n457), .IN2(a[4]), .Q(n561) );
  NOR2X0 U563 ( .IN1(n451), .IN2(n514), .QN(n560) );
  XNOR2X1 U564 ( .IN1(a[4]), .IN2(n455), .Q(n514) );
  AO22X1 U565 ( .IN1(n562), .IN2(n460), .IN3(n486), .IN4(n460), .Q(n149) );
  XOR2X1 U566 ( .IN1(n459), .IN2(a[6]), .Q(n563) );
  NOR2X0 U567 ( .IN1(n451), .IN2(n525), .QN(n562) );
  XNOR2X1 U568 ( .IN1(a[6]), .IN2(n457), .Q(n525) );
  AO22X1 U569 ( .IN1(n564), .IN2(n462), .IN3(n489), .IN4(n462), .Q(n148) );
  XOR2X1 U570 ( .IN1(n461), .IN2(a[8]), .Q(n565) );
  NOR2X0 U571 ( .IN1(n451), .IN2(n536), .QN(n564) );
  XNOR2X1 U572 ( .IN1(a[8]), .IN2(n459), .Q(n536) );
  AO22X1 U573 ( .IN1(n566), .IN2(n463), .IN3(n492), .IN4(n463), .Q(n147) );
  XOR2X1 U574 ( .IN1(n463), .IN2(a[10]), .Q(n567) );
  NOR2X0 U575 ( .IN1(n451), .IN2(n547), .QN(n566) );
  XNOR2X1 U576 ( .IN1(a[10]), .IN2(n461), .Q(n547) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_10 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_10_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_9_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n463), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n465), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n467), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n469), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n209), .B0(n220), .C1(n129), .SO(n130) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(b[4]), .ZN(n408) );
  INVX0 U312 ( .INP(n408), .ZN(n409) );
  FADDX1 U313 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U314 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U315 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U316 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U317 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR3X1 U318 ( .IN1(n96), .IN2(n103), .IN3(n410), .Q(product[10]) );
  XNOR2X1 U319 ( .IN1(n414), .IN2(n423), .Q(product[13]) );
  FADDX1 U320 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  XNOR2X1 U321 ( .IN1(n411), .IN2(n424), .Q(product[19]) );
  FADDX1 U322 ( .A(n27), .B(n461), .CI(n5), .CO(n4), .S(product[21]) );
  DELLN2X2 U323 ( .INP(n16), .Z(n410) );
  DELLN1X2 U324 ( .INP(n15), .Z(n415) );
  DELLN2X2 U325 ( .INP(n7), .Z(n411) );
  INVX0 U326 ( .INP(b[3]), .ZN(n412) );
  INVX0 U327 ( .INP(n412), .ZN(n413) );
  DELLN2X2 U328 ( .INP(n13), .Z(n414) );
  XOR2X2 U329 ( .IN1(b[10]), .IN2(n459), .Q(n490) );
  XOR2X2 U330 ( .IN1(b[10]), .IN2(n457), .Q(n487) );
  XOR2X2 U331 ( .IN1(b[10]), .IN2(n455), .Q(n484) );
  XOR2X2 U332 ( .IN1(b[10]), .IN2(n453), .Q(n481) );
  XOR2X2 U333 ( .IN1(b[10]), .IN2(n451), .Q(n473) );
  XOR2X2 U334 ( .IN1(b[10]), .IN2(a[1]), .Q(n500) );
  DELLN1X2 U335 ( .INP(b[2]), .Z(n444) );
  XOR2X2 U336 ( .IN1(b[9]), .IN2(n459), .Q(n554) );
  XOR2X2 U337 ( .IN1(b[9]), .IN2(n457), .Q(n543) );
  XOR2X2 U338 ( .IN1(b[9]), .IN2(n455), .Q(n532) );
  XOR2X2 U339 ( .IN1(b[9]), .IN2(n453), .Q(n521) );
  XOR2X2 U340 ( .IN1(b[9]), .IN2(n451), .Q(n475) );
  XOR2X2 U341 ( .IN1(b[9]), .IN2(a[1]), .Q(n499) );
  NAND2X0 U342 ( .IN1(n96), .IN2(n103), .QN(n416) );
  NAND2X0 U343 ( .IN1(n96), .IN2(n16), .QN(n417) );
  NAND2X0 U344 ( .IN1(n103), .IN2(n16), .QN(n418) );
  NAND3X0 U345 ( .IN1(n418), .IN2(n417), .IN3(n416), .QN(n15) );
  XOR2X1 U346 ( .IN1(n86), .IN2(n95), .Q(n419) );
  XOR2X1 U347 ( .IN1(n419), .IN2(n415), .Q(product[11]) );
  NAND2X0 U348 ( .IN1(n86), .IN2(n95), .QN(n420) );
  NAND2X0 U349 ( .IN1(n86), .IN2(n15), .QN(n421) );
  NAND2X0 U350 ( .IN1(n95), .IN2(n15), .QN(n422) );
  NAND3X0 U351 ( .IN1(n422), .IN2(n421), .IN3(n420), .QN(n14) );
  XOR2X2 U352 ( .IN1(b[8]), .IN2(n459), .Q(n553) );
  XOR2X2 U353 ( .IN1(b[8]), .IN2(n457), .Q(n542) );
  XOR2X2 U354 ( .IN1(b[8]), .IN2(n455), .Q(n531) );
  XOR2X2 U355 ( .IN1(b[8]), .IN2(n453), .Q(n520) );
  AO22X2 U356 ( .IN1(n449), .IN2(n499), .IN3(n476), .IN4(n498), .Q(n216) );
  XOR2X2 U357 ( .IN1(b[8]), .IN2(n451), .Q(n510) );
  XOR2X2 U358 ( .IN1(b[8]), .IN2(a[1]), .Q(n498) );
  XOR2X2 U359 ( .IN1(b[7]), .IN2(n459), .Q(n552) );
  XOR2X2 U360 ( .IN1(b[7]), .IN2(n457), .Q(n541) );
  XOR2X2 U361 ( .IN1(b[7]), .IN2(n455), .Q(n530) );
  XOR2X2 U362 ( .IN1(b[7]), .IN2(n453), .Q(n519) );
  XOR2X2 U363 ( .IN1(b[7]), .IN2(n451), .Q(n509) );
  XOR2X2 U364 ( .IN1(b[7]), .IN2(a[1]), .Q(n497) );
  XOR2X2 U365 ( .IN1(n409), .IN2(n459), .Q(n549) );
  XOR2X2 U366 ( .IN1(n409), .IN2(n457), .Q(n538) );
  XOR2X2 U367 ( .IN1(n409), .IN2(n455), .Q(n527) );
  XOR2X2 U368 ( .IN1(n409), .IN2(n453), .Q(n516) );
  XOR2X2 U369 ( .IN1(n409), .IN2(n451), .Q(n506) );
  XOR2X2 U370 ( .IN1(n409), .IN2(a[1]), .Q(n494) );
  XOR2X2 U371 ( .IN1(b[6]), .IN2(n459), .Q(n551) );
  XOR2X2 U372 ( .IN1(b[6]), .IN2(n457), .Q(n540) );
  XOR2X2 U373 ( .IN1(b[6]), .IN2(n455), .Q(n529) );
  XOR2X2 U374 ( .IN1(b[6]), .IN2(n453), .Q(n518) );
  XOR2X2 U375 ( .IN1(b[6]), .IN2(n451), .Q(n508) );
  XOR2X2 U376 ( .IN1(b[6]), .IN2(a[1]), .Q(n496) );
  XOR2X2 U377 ( .IN1(b[1]), .IN2(n459), .Q(n545) );
  XOR2X2 U378 ( .IN1(b[1]), .IN2(n457), .Q(n534) );
  XOR2X2 U379 ( .IN1(b[1]), .IN2(n455), .Q(n523) );
  XOR2X2 U380 ( .IN1(b[1]), .IN2(n453), .Q(n512) );
  XOR2X2 U381 ( .IN1(b[1]), .IN2(n451), .Q(n502) );
  XOR2X2 U382 ( .IN1(b[1]), .IN2(a[1]), .Q(n491) );
  XOR2X2 U383 ( .IN1(b[5]), .IN2(n459), .Q(n550) );
  XOR2X2 U384 ( .IN1(b[5]), .IN2(n457), .Q(n539) );
  XOR2X2 U385 ( .IN1(b[5]), .IN2(n455), .Q(n528) );
  XOR2X2 U386 ( .IN1(b[5]), .IN2(n453), .Q(n517) );
  XOR2X2 U387 ( .IN1(b[5]), .IN2(n451), .Q(n507) );
  XOR2X2 U388 ( .IN1(b[5]), .IN2(a[1]), .Q(n495) );
  XOR3X1 U389 ( .IN1(n37), .IN2(n34), .IN3(n8), .Q(product[18]) );
  XOR3X1 U390 ( .IN1(n76), .IN2(n85), .IN3(n14), .Q(product[12]) );
  XNOR2X1 U391 ( .IN1(n66), .IN2(n75), .Q(n423) );
  INVX0 U392 ( .INP(n25), .ZN(n461) );
  INVX0 U393 ( .INP(n3), .ZN(product[23]) );
  INVX0 U394 ( .INP(n55), .ZN(n467) );
  XNOR2X1 U395 ( .IN1(n33), .IN2(n30), .Q(n424) );
  XOR2X1 U396 ( .IN1(n413), .IN2(a[1]), .Q(n493) );
  XOR2X1 U397 ( .IN1(n413), .IN2(n451), .Q(n505) );
  XOR2X1 U398 ( .IN1(n413), .IN2(n453), .Q(n515) );
  INVX0 U399 ( .INP(n73), .ZN(n469) );
  XOR2X1 U400 ( .IN1(n413), .IN2(n455), .Q(n526) );
  XOR2X1 U401 ( .IN1(n413), .IN2(n457), .Q(n537) );
  INVX0 U402 ( .INP(n41), .ZN(n465) );
  INVX0 U403 ( .INP(n31), .ZN(n463) );
  XOR2X1 U404 ( .IN1(n413), .IN2(n459), .Q(n548) );
  XOR2X1 U405 ( .IN1(n444), .IN2(a[1]), .Q(n492) );
  INVX0 U406 ( .INP(n511), .ZN(n468) );
  INVX0 U407 ( .INP(n522), .ZN(n466) );
  INVX0 U408 ( .INP(n533), .ZN(n464) );
  INVX0 U409 ( .INP(n501), .ZN(n470) );
  AND2X1 U410 ( .IN1(a[1]), .IN2(n450), .Q(n476) );
  XNOR2X1 U411 ( .IN1(n425), .IN2(n132), .Q(product[4]) );
  XNOR2X1 U412 ( .IN1(n133), .IN2(n22), .Q(n425) );
  INVX0 U413 ( .INP(n544), .ZN(n462) );
  NBUFFX2 U414 ( .INP(a[5]), .Z(n454) );
  FADDX1 U415 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  NBUFFX2 U416 ( .INP(a[3]), .Z(n452) );
  AND2X1 U417 ( .IN1(n501), .IN2(n556), .Q(n474) );
  AND2X1 U418 ( .IN1(n522), .IN2(n560), .Q(n483) );
  AND2X1 U419 ( .IN1(n511), .IN2(n558), .Q(n480) );
  AND2X1 U420 ( .IN1(n533), .IN2(n562), .Q(n486) );
  AND2X1 U421 ( .IN1(n544), .IN2(n564), .Q(n489) );
  NBUFFX2 U422 ( .INP(a[7]), .Z(n456) );
  NBUFFX2 U423 ( .INP(a[9]), .Z(n458) );
  NAND2X0 U424 ( .IN1(n37), .IN2(n34), .QN(n426) );
  NAND2X0 U425 ( .IN1(n37), .IN2(n8), .QN(n427) );
  NAND2X0 U426 ( .IN1(n34), .IN2(n8), .QN(n428) );
  NAND3X0 U427 ( .IN1(n428), .IN2(n427), .IN3(n426), .QN(n7) );
  NAND2X0 U428 ( .IN1(n33), .IN2(n30), .QN(n429) );
  NAND2X0 U429 ( .IN1(n33), .IN2(n7), .QN(n430) );
  NAND2X0 U430 ( .IN1(n30), .IN2(n7), .QN(n431) );
  NAND3X0 U431 ( .IN1(n429), .IN2(n430), .IN3(n431), .QN(n6) );
  NAND2X0 U432 ( .IN1(n76), .IN2(n85), .QN(n432) );
  NAND2X0 U433 ( .IN1(n76), .IN2(n14), .QN(n433) );
  NAND2X0 U434 ( .IN1(n85), .IN2(n14), .QN(n434) );
  NAND3X0 U435 ( .IN1(n434), .IN2(n433), .IN3(n432), .QN(n13) );
  NAND2X0 U436 ( .IN1(n66), .IN2(n75), .QN(n435) );
  NAND2X0 U437 ( .IN1(n66), .IN2(n13), .QN(n436) );
  NAND2X0 U438 ( .IN1(n75), .IN2(n13), .QN(n437) );
  NAND3X0 U439 ( .IN1(n437), .IN2(n436), .IN3(n435), .QN(n12) );
  XOR3X1 U440 ( .IN1(n221), .IN2(n200), .IN3(n210), .Q(n132) );
  NAND2X0 U441 ( .IN1(n221), .IN2(n200), .QN(n438) );
  NAND2X0 U442 ( .IN1(n221), .IN2(n210), .QN(n439) );
  NAND2X0 U443 ( .IN1(n200), .IN2(n210), .QN(n440) );
  NAND3X0 U444 ( .IN1(n438), .IN2(n439), .IN3(n440), .QN(n131) );
  NAND2X0 U445 ( .IN1(n133), .IN2(n22), .QN(n441) );
  NAND2X0 U446 ( .IN1(n133), .IN2(n132), .QN(n442) );
  NAND2X0 U447 ( .IN1(n22), .IN2(n132), .QN(n443) );
  NAND3X0 U448 ( .IN1(n441), .IN2(n442), .IN3(n443), .QN(n21) );
  DELLN1X2 U449 ( .INP(a[11]), .Z(n459) );
  INVX0 U450 ( .INP(n448), .ZN(n445) );
  INVX0 U451 ( .INP(b[0]), .ZN(n446) );
  INVX0 U452 ( .INP(b[0]), .ZN(n447) );
  INVX0 U453 ( .INP(b[0]), .ZN(n448) );
  INVX0 U454 ( .INP(n450), .ZN(n449) );
  INVX0 U455 ( .INP(a[0]), .ZN(n450) );
  DELLN1X2 U456 ( .INP(a[3]), .Z(n451) );
  DELLN1X2 U457 ( .INP(a[5]), .Z(n453) );
  DELLN1X2 U458 ( .INP(a[7]), .Z(n455) );
  DELLN1X2 U459 ( .INP(a[9]), .Z(n457) );
  NOR2X0 U460 ( .IN1(n450), .IN2(n447), .QN(product[0]) );
  XNOR2X1 U461 ( .IN1(n471), .IN2(n472), .Q(n84) );
  NAND2X0 U462 ( .IN1(n472), .IN2(n471), .QN(n83) );
  AOI22X1 U463 ( .IN1(n473), .IN2(n470), .IN3(n474), .IN4(n475), .QN(n471) );
  OA21X1 U464 ( .IN1(n476), .IN2(n449), .IN3(n477), .Q(n472) );
  AO22X1 U465 ( .IN1(n478), .IN2(n470), .IN3(n474), .IN4(n473), .Q(n73) );
  AO22X1 U466 ( .IN1(n479), .IN2(n468), .IN3(n480), .IN4(n481), .Q(n55) );
  AO22X1 U467 ( .IN1(n482), .IN2(n466), .IN3(n483), .IN4(n484), .Q(n41) );
  AO22X1 U468 ( .IN1(n485), .IN2(n464), .IN3(n486), .IN4(n487), .Q(n31) );
  AO22X1 U469 ( .IN1(n488), .IN2(n462), .IN3(n489), .IN4(n490), .Q(n25) );
  AO22X1 U470 ( .IN1(n449), .IN2(n491), .IN3(n476), .IN4(n448), .Q(n224) );
  AO22X1 U471 ( .IN1(n449), .IN2(n492), .IN3(n476), .IN4(n491), .Q(n223) );
  AO22X1 U472 ( .IN1(n449), .IN2(n493), .IN3(n476), .IN4(n492), .Q(n222) );
  AO22X1 U473 ( .IN1(n449), .IN2(n494), .IN3(n476), .IN4(n493), .Q(n221) );
  AO22X1 U474 ( .IN1(n449), .IN2(n495), .IN3(n476), .IN4(n494), .Q(n220) );
  AO22X1 U475 ( .IN1(n449), .IN2(n496), .IN3(n495), .IN4(n476), .Q(n219) );
  AO22X1 U476 ( .IN1(n449), .IN2(n497), .IN3(n476), .IN4(n496), .Q(n218) );
  AO22X1 U477 ( .IN1(n449), .IN2(n498), .IN3(n476), .IN4(n497), .Q(n217) );
  AO22X1 U478 ( .IN1(n449), .IN2(n500), .IN3(n476), .IN4(n499), .Q(n215) );
  AO22X1 U479 ( .IN1(n449), .IN2(n477), .IN3(n476), .IN4(n500), .Q(n214) );
  XOR2X1 U480 ( .IN1(b[11]), .IN2(a[1]), .Q(n477) );
  NOR2X0 U481 ( .IN1(n501), .IN2(n447), .QN(n212) );
  AO22X1 U482 ( .IN1(n502), .IN2(n470), .IN3(n474), .IN4(n503), .Q(n211) );
  XOR2X1 U483 ( .IN1(n445), .IN2(n451), .Q(n503) );
  AO22X1 U484 ( .IN1(n504), .IN2(n470), .IN3(n474), .IN4(n502), .Q(n210) );
  AO22X1 U485 ( .IN1(n505), .IN2(n470), .IN3(n474), .IN4(n504), .Q(n209) );
  XOR2X1 U486 ( .IN1(n444), .IN2(n451), .Q(n504) );
  AO22X1 U487 ( .IN1(n506), .IN2(n470), .IN3(n474), .IN4(n505), .Q(n208) );
  AO22X1 U488 ( .IN1(n507), .IN2(n470), .IN3(n474), .IN4(n506), .Q(n207) );
  AO22X1 U489 ( .IN1(n508), .IN2(n470), .IN3(n474), .IN4(n507), .Q(n206) );
  AO22X1 U490 ( .IN1(n509), .IN2(n470), .IN3(n474), .IN4(n508), .Q(n205) );
  AO22X1 U491 ( .IN1(n510), .IN2(n470), .IN3(n474), .IN4(n509), .Q(n204) );
  AO22X1 U492 ( .IN1(n475), .IN2(n470), .IN3(n474), .IN4(n510), .Q(n203) );
  OAI21X1 U493 ( .IN1(n470), .IN2(n474), .IN3(n478), .QN(n201) );
  XOR2X1 U494 ( .IN1(b[11]), .IN2(n451), .Q(n478) );
  NOR2X0 U495 ( .IN1(n511), .IN2(n447), .QN(n200) );
  AO22X1 U496 ( .IN1(n512), .IN2(n468), .IN3(n480), .IN4(n513), .Q(n199) );
  XOR2X1 U497 ( .IN1(n445), .IN2(n453), .Q(n513) );
  AO22X1 U498 ( .IN1(n514), .IN2(n468), .IN3(n480), .IN4(n512), .Q(n198) );
  AO22X1 U499 ( .IN1(n515), .IN2(n468), .IN3(n480), .IN4(n514), .Q(n197) );
  XOR2X1 U500 ( .IN1(n444), .IN2(n453), .Q(n514) );
  AO22X1 U501 ( .IN1(n516), .IN2(n468), .IN3(n480), .IN4(n515), .Q(n196) );
  AO22X1 U502 ( .IN1(n517), .IN2(n468), .IN3(n480), .IN4(n516), .Q(n195) );
  AO22X1 U503 ( .IN1(n518), .IN2(n468), .IN3(n480), .IN4(n517), .Q(n194) );
  AO22X1 U504 ( .IN1(n519), .IN2(n468), .IN3(n480), .IN4(n518), .Q(n193) );
  AO22X1 U505 ( .IN1(n520), .IN2(n468), .IN3(n480), .IN4(n519), .Q(n192) );
  AO22X1 U506 ( .IN1(n521), .IN2(n468), .IN3(n480), .IN4(n520), .Q(n191) );
  AO22X1 U507 ( .IN1(n481), .IN2(n468), .IN3(n480), .IN4(n521), .Q(n190) );
  OAI21X1 U508 ( .IN1(n468), .IN2(n480), .IN3(n479), .QN(n189) );
  XOR2X1 U509 ( .IN1(b[11]), .IN2(n453), .Q(n479) );
  NOR2X0 U510 ( .IN1(n522), .IN2(n446), .QN(n188) );
  AO22X1 U511 ( .IN1(n523), .IN2(n466), .IN3(n483), .IN4(n524), .Q(n187) );
  XOR2X1 U512 ( .IN1(n445), .IN2(n455), .Q(n524) );
  AO22X1 U513 ( .IN1(n525), .IN2(n466), .IN3(n483), .IN4(n523), .Q(n186) );
  AO22X1 U514 ( .IN1(n526), .IN2(n466), .IN3(n483), .IN4(n525), .Q(n185) );
  XOR2X1 U515 ( .IN1(n444), .IN2(n455), .Q(n525) );
  AO22X1 U516 ( .IN1(n527), .IN2(n466), .IN3(n483), .IN4(n526), .Q(n184) );
  AO22X1 U517 ( .IN1(n528), .IN2(n466), .IN3(n483), .IN4(n527), .Q(n183) );
  AO22X1 U518 ( .IN1(n529), .IN2(n466), .IN3(n483), .IN4(n528), .Q(n182) );
  AO22X1 U519 ( .IN1(n530), .IN2(n466), .IN3(n483), .IN4(n529), .Q(n181) );
  AO22X1 U520 ( .IN1(n531), .IN2(n466), .IN3(n483), .IN4(n530), .Q(n180) );
  AO22X1 U521 ( .IN1(n532), .IN2(n466), .IN3(n483), .IN4(n531), .Q(n179) );
  AO22X1 U522 ( .IN1(n484), .IN2(n466), .IN3(n483), .IN4(n532), .Q(n178) );
  OAI21X1 U523 ( .IN1(n466), .IN2(n483), .IN3(n482), .QN(n177) );
  XOR2X1 U524 ( .IN1(b[11]), .IN2(n455), .Q(n482) );
  NOR2X0 U525 ( .IN1(n533), .IN2(n446), .QN(n176) );
  AO22X1 U526 ( .IN1(n534), .IN2(n464), .IN3(n486), .IN4(n535), .Q(n175) );
  XOR2X1 U527 ( .IN1(n445), .IN2(n457), .Q(n535) );
  AO22X1 U528 ( .IN1(n536), .IN2(n464), .IN3(n486), .IN4(n534), .Q(n174) );
  AO22X1 U529 ( .IN1(n537), .IN2(n464), .IN3(n486), .IN4(n536), .Q(n173) );
  XOR2X1 U530 ( .IN1(n444), .IN2(n457), .Q(n536) );
  AO22X1 U531 ( .IN1(n538), .IN2(n464), .IN3(n486), .IN4(n537), .Q(n172) );
  AO22X1 U532 ( .IN1(n539), .IN2(n464), .IN3(n486), .IN4(n538), .Q(n171) );
  AO22X1 U533 ( .IN1(n540), .IN2(n464), .IN3(n486), .IN4(n539), .Q(n170) );
  AO22X1 U534 ( .IN1(n541), .IN2(n464), .IN3(n486), .IN4(n540), .Q(n169) );
  AO22X1 U535 ( .IN1(n542), .IN2(n464), .IN3(n486), .IN4(n541), .Q(n168) );
  AO22X1 U536 ( .IN1(n543), .IN2(n464), .IN3(n486), .IN4(n542), .Q(n167) );
  AO22X1 U537 ( .IN1(n487), .IN2(n464), .IN3(n486), .IN4(n543), .Q(n166) );
  OAI21X1 U538 ( .IN1(n464), .IN2(n486), .IN3(n485), .QN(n165) );
  XOR2X1 U539 ( .IN1(b[11]), .IN2(n457), .Q(n485) );
  NOR2X0 U540 ( .IN1(n544), .IN2(n446), .QN(n164) );
  AO22X1 U541 ( .IN1(n545), .IN2(n462), .IN3(n489), .IN4(n546), .Q(n163) );
  XOR2X1 U542 ( .IN1(n445), .IN2(n459), .Q(n546) );
  AO22X1 U543 ( .IN1(n547), .IN2(n462), .IN3(n489), .IN4(n545), .Q(n162) );
  AO22X1 U544 ( .IN1(n548), .IN2(n462), .IN3(n489), .IN4(n547), .Q(n161) );
  XOR2X1 U545 ( .IN1(n444), .IN2(n459), .Q(n547) );
  AO22X1 U546 ( .IN1(n549), .IN2(n462), .IN3(n489), .IN4(n548), .Q(n160) );
  AO22X1 U547 ( .IN1(n550), .IN2(n462), .IN3(n489), .IN4(n549), .Q(n159) );
  AO22X1 U548 ( .IN1(n551), .IN2(n462), .IN3(n489), .IN4(n550), .Q(n158) );
  AO22X1 U549 ( .IN1(n552), .IN2(n462), .IN3(n489), .IN4(n551), .Q(n157) );
  AO22X1 U550 ( .IN1(n553), .IN2(n462), .IN3(n489), .IN4(n552), .Q(n156) );
  AO22X1 U551 ( .IN1(n554), .IN2(n462), .IN3(n489), .IN4(n553), .Q(n155) );
  AO22X1 U552 ( .IN1(n490), .IN2(n462), .IN3(n489), .IN4(n554), .Q(n154) );
  OAI21X1 U553 ( .IN1(n462), .IN2(n489), .IN3(n488), .QN(n153) );
  XOR2X1 U554 ( .IN1(b[11]), .IN2(n459), .Q(n488) );
  AO21X1 U555 ( .IN1(a[1]), .IN2(n448), .IN3(n476), .Q(n152) );
  AO22X1 U556 ( .IN1(n555), .IN2(n452), .IN3(n474), .IN4(n452), .Q(n151) );
  XOR2X1 U557 ( .IN1(n451), .IN2(a[2]), .Q(n556) );
  NOR2X0 U558 ( .IN1(n445), .IN2(n501), .QN(n555) );
  XNOR2X1 U559 ( .IN1(a[2]), .IN2(a[1]), .Q(n501) );
  AO22X1 U560 ( .IN1(n557), .IN2(n454), .IN3(n480), .IN4(n454), .Q(n150) );
  XOR2X1 U561 ( .IN1(n453), .IN2(a[4]), .Q(n558) );
  NOR2X0 U562 ( .IN1(n445), .IN2(n511), .QN(n557) );
  XNOR2X1 U563 ( .IN1(a[4]), .IN2(n451), .Q(n511) );
  AO22X1 U564 ( .IN1(n559), .IN2(n456), .IN3(n483), .IN4(n456), .Q(n149) );
  XOR2X1 U565 ( .IN1(n455), .IN2(a[6]), .Q(n560) );
  NOR2X0 U566 ( .IN1(n445), .IN2(n522), .QN(n559) );
  XNOR2X1 U567 ( .IN1(a[6]), .IN2(n453), .Q(n522) );
  AO22X1 U568 ( .IN1(n561), .IN2(n458), .IN3(n486), .IN4(n458), .Q(n148) );
  XOR2X1 U569 ( .IN1(n457), .IN2(a[8]), .Q(n562) );
  NOR2X0 U570 ( .IN1(n445), .IN2(n533), .QN(n561) );
  XNOR2X1 U571 ( .IN1(a[8]), .IN2(n455), .Q(n533) );
  AO22X1 U572 ( .IN1(n563), .IN2(n459), .IN3(n489), .IN4(n459), .Q(n147) );
  XOR2X1 U573 ( .IN1(n459), .IN2(a[10]), .Q(n564) );
  NOR2X0 U574 ( .IN1(n445), .IN2(n544), .QN(n563) );
  XNOR2X1 U575 ( .IN1(a[10]), .IN2(n457), .Q(n544) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_9 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_9_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_8_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n449), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n451), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n453), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n455), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n457), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  DELLN1X2 U311 ( .INP(b[8]), .Z(n408) );
  XOR2X1 U312 ( .IN1(n433), .IN2(n439), .Q(n491) );
  INVX0 U313 ( .INP(b[1]), .ZN(n409) );
  INVX0 U314 ( .INP(n409), .ZN(n410) );
  INVX0 U315 ( .INP(b[6]), .ZN(n411) );
  INVX0 U316 ( .INP(n411), .ZN(n412) );
  INVX0 U317 ( .INP(n436), .ZN(n413) );
  INVX0 U318 ( .INP(n436), .ZN(n414) );
  DELLN2X2 U319 ( .INP(n9), .Z(n415) );
  XOR2X2 U320 ( .IN1(n413), .IN2(n447), .Q(n534) );
  XOR2X2 U321 ( .IN1(n413), .IN2(n445), .Q(n523) );
  XOR2X2 U322 ( .IN1(n414), .IN2(n443), .Q(n512) );
  XOR2X2 U323 ( .IN1(n413), .IN2(n441), .Q(n501) );
  DELLN2X2 U324 ( .INP(n15), .Z(n416) );
  INVX0 U325 ( .INP(b[3]), .ZN(n417) );
  INVX0 U326 ( .INP(n417), .ZN(n418) );
  XOR2X2 U327 ( .IN1(b[2]), .IN2(n447), .Q(n535) );
  XOR2X2 U328 ( .IN1(b[2]), .IN2(n445), .Q(n524) );
  XOR2X2 U329 ( .IN1(b[2]), .IN2(n443), .Q(n513) );
  XOR2X2 U330 ( .IN1(b[2]), .IN2(n441), .Q(n502) );
  XOR2X2 U331 ( .IN1(b[2]), .IN2(n439), .Q(n492) );
  XOR2X2 U332 ( .IN1(b[2]), .IN2(a[1]), .Q(n480) );
  XOR2X2 U333 ( .IN1(b[10]), .IN2(n447), .Q(n478) );
  XOR2X2 U334 ( .IN1(b[10]), .IN2(n445), .Q(n475) );
  XOR2X2 U335 ( .IN1(b[10]), .IN2(n443), .Q(n472) );
  XOR2X2 U336 ( .IN1(b[10]), .IN2(n441), .Q(n469) );
  XOR2X2 U337 ( .IN1(b[10]), .IN2(n439), .Q(n461) );
  XOR2X2 U338 ( .IN1(b[10]), .IN2(a[1]), .Q(n488) );
  XOR2X2 U339 ( .IN1(b[9]), .IN2(n447), .Q(n542) );
  XOR2X2 U340 ( .IN1(b[9]), .IN2(n445), .Q(n531) );
  XOR2X2 U341 ( .IN1(b[9]), .IN2(n443), .Q(n520) );
  XOR2X2 U342 ( .IN1(b[9]), .IN2(n441), .Q(n509) );
  XOR2X2 U343 ( .IN1(b[9]), .IN2(n439), .Q(n463) );
  XOR2X2 U344 ( .IN1(b[9]), .IN2(a[1]), .Q(n487) );
  XOR2X2 U345 ( .IN1(n408), .IN2(n447), .Q(n541) );
  XOR2X2 U346 ( .IN1(n408), .IN2(n445), .Q(n530) );
  XOR2X2 U347 ( .IN1(n408), .IN2(n443), .Q(n519) );
  XOR2X2 U348 ( .IN1(n408), .IN2(n441), .Q(n508) );
  XOR2X2 U349 ( .IN1(n408), .IN2(n439), .Q(n498) );
  XOR2X2 U350 ( .IN1(n408), .IN2(a[1]), .Q(n486) );
  XOR2X2 U351 ( .IN1(n412), .IN2(n447), .Q(n539) );
  XOR2X2 U352 ( .IN1(n412), .IN2(n445), .Q(n528) );
  XOR2X2 U353 ( .IN1(n412), .IN2(n443), .Q(n517) );
  XOR2X2 U354 ( .IN1(n412), .IN2(n441), .Q(n506) );
  XOR2X2 U355 ( .IN1(n412), .IN2(n439), .Q(n496) );
  XOR2X2 U356 ( .IN1(n412), .IN2(a[1]), .Q(n484) );
  XOR2X2 U357 ( .IN1(n410), .IN2(n447), .Q(n533) );
  XOR2X2 U358 ( .IN1(n410), .IN2(n445), .Q(n522) );
  XOR2X2 U359 ( .IN1(n410), .IN2(n443), .Q(n511) );
  XOR2X2 U360 ( .IN1(n410), .IN2(n441), .Q(n500) );
  XOR2X2 U361 ( .IN1(n410), .IN2(n439), .Q(n490) );
  XOR2X2 U362 ( .IN1(n410), .IN2(a[1]), .Q(n479) );
  FADDX1 U363 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U364 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  XNOR2X1 U365 ( .IN1(n419), .IN2(n415), .Q(product[17]) );
  XNOR2X1 U366 ( .IN1(n43), .IN2(n38), .Q(n419) );
  XOR3X1 U367 ( .IN1(n49), .IN2(n44), .IN3(n10), .Q(product[16]) );
  XOR3X1 U368 ( .IN1(n96), .IN2(n103), .IN3(n16), .Q(product[10]) );
  XNOR2X1 U369 ( .IN1(n420), .IN2(n416), .Q(product[11]) );
  XNOR2X1 U370 ( .IN1(n86), .IN2(n95), .Q(n420) );
  INVX0 U371 ( .INP(n25), .ZN(n449) );
  FADDX1 U372 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  INVX0 U373 ( .INP(n3), .ZN(product[23]) );
  INVX0 U374 ( .INP(n55), .ZN(n455) );
  FADDX1 U375 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U376 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X1 U377 ( .IN1(n418), .IN2(a[1]), .Q(n481) );
  XOR2X1 U378 ( .IN1(n418), .IN2(n439), .Q(n493) );
  XOR2X1 U379 ( .IN1(n418), .IN2(n441), .Q(n503) );
  INVX0 U380 ( .INP(n73), .ZN(n457) );
  XOR2X1 U381 ( .IN1(n418), .IN2(n443), .Q(n514) );
  XOR2X1 U382 ( .IN1(n418), .IN2(n445), .Q(n525) );
  INVX0 U383 ( .INP(n31), .ZN(n451) );
  INVX0 U384 ( .INP(n41), .ZN(n453) );
  XOR2X1 U385 ( .IN1(n418), .IN2(n447), .Q(n536) );
  INVX0 U386 ( .INP(n489), .ZN(n458) );
  INVX0 U387 ( .INP(n499), .ZN(n456) );
  INVX0 U388 ( .INP(n510), .ZN(n454) );
  INVX0 U389 ( .INP(n521), .ZN(n452) );
  AND2X1 U390 ( .IN1(a[1]), .IN2(n438), .Q(n464) );
  INVX0 U391 ( .INP(n532), .ZN(n450) );
  FADDX1 U392 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  NBUFFX2 U393 ( .INP(a[3]), .Z(n440) );
  NBUFFX2 U394 ( .INP(a[9]), .Z(n446) );
  NBUFFX2 U395 ( .INP(a[7]), .Z(n444) );
  NAND2X0 U396 ( .IN1(n49), .IN2(n44), .QN(n421) );
  NAND2X0 U397 ( .IN1(n49), .IN2(n10), .QN(n422) );
  NAND2X0 U398 ( .IN1(n44), .IN2(n10), .QN(n423) );
  NAND3X0 U399 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n9) );
  NAND2X0 U400 ( .IN1(n43), .IN2(n38), .QN(n424) );
  NAND2X0 U401 ( .IN1(n43), .IN2(n9), .QN(n425) );
  NAND2X0 U402 ( .IN1(n38), .IN2(n9), .QN(n426) );
  NAND3X0 U403 ( .IN1(n426), .IN2(n425), .IN3(n424), .QN(n8) );
  NAND2X0 U404 ( .IN1(n96), .IN2(n103), .QN(n427) );
  NAND2X0 U405 ( .IN1(n96), .IN2(n16), .QN(n428) );
  NAND2X0 U406 ( .IN1(n103), .IN2(n16), .QN(n429) );
  NAND3X0 U407 ( .IN1(n427), .IN2(n428), .IN3(n429), .QN(n15) );
  NAND2X0 U408 ( .IN1(n86), .IN2(n95), .QN(n430) );
  NAND2X0 U409 ( .IN1(n86), .IN2(n15), .QN(n431) );
  NAND2X0 U410 ( .IN1(n95), .IN2(n15), .QN(n432) );
  NAND3X0 U411 ( .IN1(n432), .IN2(n431), .IN3(n430), .QN(n14) );
  DELLN1X2 U412 ( .INP(a[11]), .Z(n447) );
  AND2X2 U413 ( .IN1(n489), .IN2(n544), .Q(n462) );
  AND2X2 U414 ( .IN1(n499), .IN2(n546), .Q(n468) );
  AND2X2 U415 ( .IN1(n510), .IN2(n548), .Q(n471) );
  AND2X2 U416 ( .IN1(n521), .IN2(n550), .Q(n474) );
  AND2X2 U417 ( .IN1(n532), .IN2(n552), .Q(n477) );
  INVX0 U418 ( .INP(n436), .ZN(n433) );
  INVX0 U419 ( .INP(b[0]), .ZN(n434) );
  INVX0 U420 ( .INP(b[0]), .ZN(n435) );
  INVX0 U421 ( .INP(b[0]), .ZN(n436) );
  INVX0 U422 ( .INP(n438), .ZN(n437) );
  INVX0 U423 ( .INP(a[0]), .ZN(n438) );
  DELLN1X2 U424 ( .INP(a[3]), .Z(n439) );
  DELLN1X2 U425 ( .INP(a[5]), .Z(n441) );
  DELLN1X2 U426 ( .INP(a[5]), .Z(n442) );
  DELLN1X2 U427 ( .INP(a[7]), .Z(n443) );
  DELLN1X2 U428 ( .INP(a[9]), .Z(n445) );
  NOR2X0 U429 ( .IN1(n438), .IN2(n435), .QN(product[0]) );
  XNOR2X1 U430 ( .IN1(n459), .IN2(n460), .Q(n84) );
  NAND2X0 U431 ( .IN1(n460), .IN2(n459), .QN(n83) );
  AOI22X1 U432 ( .IN1(n461), .IN2(n458), .IN3(n462), .IN4(n463), .QN(n459) );
  OA21X1 U433 ( .IN1(n464), .IN2(n437), .IN3(n465), .Q(n460) );
  AO22X1 U434 ( .IN1(n466), .IN2(n458), .IN3(n462), .IN4(n461), .Q(n73) );
  AO22X1 U435 ( .IN1(n467), .IN2(n456), .IN3(n468), .IN4(n469), .Q(n55) );
  AO22X1 U436 ( .IN1(n470), .IN2(n454), .IN3(n471), .IN4(n472), .Q(n41) );
  AO22X1 U437 ( .IN1(n473), .IN2(n452), .IN3(n474), .IN4(n475), .Q(n31) );
  AO22X1 U438 ( .IN1(n476), .IN2(n450), .IN3(n477), .IN4(n478), .Q(n25) );
  AO22X1 U439 ( .IN1(n437), .IN2(n479), .IN3(n464), .IN4(n436), .Q(n224) );
  AO22X1 U440 ( .IN1(n437), .IN2(n480), .IN3(n464), .IN4(n479), .Q(n223) );
  AO22X1 U441 ( .IN1(n437), .IN2(n481), .IN3(n464), .IN4(n480), .Q(n222) );
  AO22X1 U442 ( .IN1(n437), .IN2(n482), .IN3(n464), .IN4(n481), .Q(n221) );
  AO22X1 U443 ( .IN1(n437), .IN2(n483), .IN3(n464), .IN4(n482), .Q(n220) );
  XOR2X1 U444 ( .IN1(b[4]), .IN2(a[1]), .Q(n482) );
  AO22X1 U445 ( .IN1(n437), .IN2(n484), .IN3(n464), .IN4(n483), .Q(n219) );
  XOR2X1 U446 ( .IN1(b[5]), .IN2(a[1]), .Q(n483) );
  AO22X1 U447 ( .IN1(n437), .IN2(n485), .IN3(n464), .IN4(n484), .Q(n218) );
  AO22X1 U448 ( .IN1(n437), .IN2(n486), .IN3(n464), .IN4(n485), .Q(n217) );
  XOR2X1 U449 ( .IN1(b[7]), .IN2(a[1]), .Q(n485) );
  AO22X1 U450 ( .IN1(n437), .IN2(n487), .IN3(n464), .IN4(n486), .Q(n216) );
  AO22X1 U451 ( .IN1(n437), .IN2(n488), .IN3(n464), .IN4(n487), .Q(n215) );
  AO22X1 U452 ( .IN1(n437), .IN2(n465), .IN3(n464), .IN4(n488), .Q(n214) );
  XOR2X1 U453 ( .IN1(b[11]), .IN2(a[1]), .Q(n465) );
  NOR2X0 U454 ( .IN1(n489), .IN2(n435), .QN(n212) );
  AO22X1 U455 ( .IN1(n490), .IN2(n458), .IN3(n462), .IN4(n491), .Q(n211) );
  AO22X1 U456 ( .IN1(n492), .IN2(n458), .IN3(n462), .IN4(n490), .Q(n210) );
  AO22X1 U457 ( .IN1(n493), .IN2(n458), .IN3(n462), .IN4(n492), .Q(n209) );
  AO22X1 U458 ( .IN1(n494), .IN2(n458), .IN3(n462), .IN4(n493), .Q(n208) );
  AO22X1 U459 ( .IN1(n495), .IN2(n458), .IN3(n462), .IN4(n494), .Q(n207) );
  XOR2X1 U460 ( .IN1(b[4]), .IN2(n439), .Q(n494) );
  AO22X1 U461 ( .IN1(n496), .IN2(n458), .IN3(n462), .IN4(n495), .Q(n206) );
  XOR2X1 U462 ( .IN1(b[5]), .IN2(n439), .Q(n495) );
  AO22X1 U463 ( .IN1(n497), .IN2(n458), .IN3(n462), .IN4(n496), .Q(n205) );
  AO22X1 U464 ( .IN1(n498), .IN2(n458), .IN3(n462), .IN4(n497), .Q(n204) );
  XOR2X1 U465 ( .IN1(b[7]), .IN2(n439), .Q(n497) );
  AO22X1 U466 ( .IN1(n463), .IN2(n458), .IN3(n462), .IN4(n498), .Q(n203) );
  OAI21X1 U467 ( .IN1(n458), .IN2(n462), .IN3(n466), .QN(n201) );
  XOR2X1 U468 ( .IN1(b[11]), .IN2(n439), .Q(n466) );
  NOR2X0 U469 ( .IN1(n499), .IN2(n435), .QN(n200) );
  AO22X1 U470 ( .IN1(n500), .IN2(n456), .IN3(n468), .IN4(n501), .Q(n199) );
  AO22X1 U471 ( .IN1(n502), .IN2(n456), .IN3(n468), .IN4(n500), .Q(n198) );
  AO22X1 U472 ( .IN1(n503), .IN2(n456), .IN3(n468), .IN4(n502), .Q(n197) );
  AO22X1 U473 ( .IN1(n504), .IN2(n456), .IN3(n468), .IN4(n503), .Q(n196) );
  AO22X1 U474 ( .IN1(n505), .IN2(n456), .IN3(n468), .IN4(n504), .Q(n195) );
  XOR2X1 U475 ( .IN1(b[4]), .IN2(n441), .Q(n504) );
  AO22X1 U476 ( .IN1(n506), .IN2(n456), .IN3(n468), .IN4(n505), .Q(n194) );
  XOR2X1 U477 ( .IN1(b[5]), .IN2(n441), .Q(n505) );
  AO22X1 U478 ( .IN1(n507), .IN2(n456), .IN3(n468), .IN4(n506), .Q(n193) );
  AO22X1 U479 ( .IN1(n508), .IN2(n456), .IN3(n468), .IN4(n507), .Q(n192) );
  XOR2X1 U480 ( .IN1(b[7]), .IN2(n441), .Q(n507) );
  AO22X1 U481 ( .IN1(n509), .IN2(n456), .IN3(n468), .IN4(n508), .Q(n191) );
  AO22X1 U482 ( .IN1(n469), .IN2(n456), .IN3(n468), .IN4(n509), .Q(n190) );
  OAI21X1 U483 ( .IN1(n456), .IN2(n468), .IN3(n467), .QN(n189) );
  XOR2X1 U484 ( .IN1(b[11]), .IN2(n441), .Q(n467) );
  NOR2X0 U485 ( .IN1(n510), .IN2(n434), .QN(n188) );
  AO22X1 U486 ( .IN1(n511), .IN2(n454), .IN3(n471), .IN4(n512), .Q(n187) );
  AO22X1 U487 ( .IN1(n513), .IN2(n454), .IN3(n471), .IN4(n511), .Q(n186) );
  AO22X1 U488 ( .IN1(n514), .IN2(n454), .IN3(n471), .IN4(n513), .Q(n185) );
  AO22X1 U489 ( .IN1(n515), .IN2(n454), .IN3(n471), .IN4(n514), .Q(n184) );
  AO22X1 U490 ( .IN1(n516), .IN2(n454), .IN3(n471), .IN4(n515), .Q(n183) );
  XOR2X1 U491 ( .IN1(b[4]), .IN2(n443), .Q(n515) );
  AO22X1 U492 ( .IN1(n517), .IN2(n454), .IN3(n471), .IN4(n516), .Q(n182) );
  XOR2X1 U493 ( .IN1(b[5]), .IN2(n443), .Q(n516) );
  AO22X1 U494 ( .IN1(n518), .IN2(n454), .IN3(n471), .IN4(n517), .Q(n181) );
  AO22X1 U495 ( .IN1(n519), .IN2(n454), .IN3(n471), .IN4(n518), .Q(n180) );
  XOR2X1 U496 ( .IN1(b[7]), .IN2(n443), .Q(n518) );
  AO22X1 U497 ( .IN1(n520), .IN2(n454), .IN3(n471), .IN4(n519), .Q(n179) );
  AO22X1 U498 ( .IN1(n472), .IN2(n454), .IN3(n471), .IN4(n520), .Q(n178) );
  OAI21X1 U499 ( .IN1(n454), .IN2(n471), .IN3(n470), .QN(n177) );
  XOR2X1 U500 ( .IN1(b[11]), .IN2(n443), .Q(n470) );
  NOR2X0 U501 ( .IN1(n521), .IN2(n434), .QN(n176) );
  AO22X1 U502 ( .IN1(n522), .IN2(n452), .IN3(n474), .IN4(n523), .Q(n175) );
  AO22X1 U503 ( .IN1(n524), .IN2(n452), .IN3(n474), .IN4(n522), .Q(n174) );
  AO22X1 U504 ( .IN1(n525), .IN2(n452), .IN3(n474), .IN4(n524), .Q(n173) );
  AO22X1 U505 ( .IN1(n526), .IN2(n452), .IN3(n474), .IN4(n525), .Q(n172) );
  AO22X1 U506 ( .IN1(n527), .IN2(n452), .IN3(n474), .IN4(n526), .Q(n171) );
  XOR2X1 U507 ( .IN1(b[4]), .IN2(n445), .Q(n526) );
  AO22X1 U508 ( .IN1(n528), .IN2(n452), .IN3(n474), .IN4(n527), .Q(n170) );
  XOR2X1 U509 ( .IN1(b[5]), .IN2(n445), .Q(n527) );
  AO22X1 U510 ( .IN1(n529), .IN2(n452), .IN3(n474), .IN4(n528), .Q(n169) );
  AO22X1 U511 ( .IN1(n530), .IN2(n452), .IN3(n474), .IN4(n529), .Q(n168) );
  XOR2X1 U512 ( .IN1(b[7]), .IN2(n445), .Q(n529) );
  AO22X1 U513 ( .IN1(n531), .IN2(n452), .IN3(n474), .IN4(n530), .Q(n167) );
  AO22X1 U514 ( .IN1(n475), .IN2(n452), .IN3(n474), .IN4(n531), .Q(n166) );
  OAI21X1 U515 ( .IN1(n452), .IN2(n474), .IN3(n473), .QN(n165) );
  XOR2X1 U516 ( .IN1(b[11]), .IN2(n445), .Q(n473) );
  NOR2X0 U517 ( .IN1(n532), .IN2(n434), .QN(n164) );
  AO22X1 U518 ( .IN1(n533), .IN2(n450), .IN3(n477), .IN4(n534), .Q(n163) );
  AO22X1 U519 ( .IN1(n535), .IN2(n450), .IN3(n477), .IN4(n533), .Q(n162) );
  AO22X1 U520 ( .IN1(n536), .IN2(n450), .IN3(n477), .IN4(n535), .Q(n161) );
  AO22X1 U521 ( .IN1(n537), .IN2(n450), .IN3(n477), .IN4(n536), .Q(n160) );
  AO22X1 U522 ( .IN1(n538), .IN2(n450), .IN3(n477), .IN4(n537), .Q(n159) );
  XOR2X1 U523 ( .IN1(b[4]), .IN2(n447), .Q(n537) );
  AO22X1 U524 ( .IN1(n539), .IN2(n450), .IN3(n477), .IN4(n538), .Q(n158) );
  XOR2X1 U525 ( .IN1(b[5]), .IN2(n447), .Q(n538) );
  AO22X1 U526 ( .IN1(n540), .IN2(n450), .IN3(n477), .IN4(n539), .Q(n157) );
  AO22X1 U527 ( .IN1(n541), .IN2(n450), .IN3(n477), .IN4(n540), .Q(n156) );
  XOR2X1 U528 ( .IN1(b[7]), .IN2(n447), .Q(n540) );
  AO22X1 U529 ( .IN1(n542), .IN2(n450), .IN3(n477), .IN4(n541), .Q(n155) );
  AO22X1 U530 ( .IN1(n478), .IN2(n450), .IN3(n477), .IN4(n542), .Q(n154) );
  OAI21X1 U531 ( .IN1(n450), .IN2(n477), .IN3(n476), .QN(n153) );
  XOR2X1 U532 ( .IN1(b[11]), .IN2(n447), .Q(n476) );
  AO21X1 U533 ( .IN1(a[1]), .IN2(n436), .IN3(n464), .Q(n152) );
  AO22X1 U534 ( .IN1(n543), .IN2(n440), .IN3(n462), .IN4(n440), .Q(n151) );
  XOR2X1 U535 ( .IN1(n439), .IN2(a[2]), .Q(n544) );
  NOR2X0 U536 ( .IN1(n414), .IN2(n489), .QN(n543) );
  XNOR2X1 U537 ( .IN1(a[2]), .IN2(a[1]), .Q(n489) );
  AO22X1 U538 ( .IN1(n545), .IN2(n442), .IN3(n468), .IN4(n442), .Q(n150) );
  XOR2X1 U539 ( .IN1(n441), .IN2(a[4]), .Q(n546) );
  NOR2X0 U540 ( .IN1(n414), .IN2(n499), .QN(n545) );
  XNOR2X1 U541 ( .IN1(a[4]), .IN2(n439), .Q(n499) );
  AO22X1 U542 ( .IN1(n547), .IN2(n444), .IN3(n471), .IN4(n444), .Q(n149) );
  XOR2X1 U543 ( .IN1(n443), .IN2(a[6]), .Q(n548) );
  NOR2X0 U544 ( .IN1(n413), .IN2(n510), .QN(n547) );
  XNOR2X1 U545 ( .IN1(a[6]), .IN2(n441), .Q(n510) );
  AO22X1 U546 ( .IN1(n549), .IN2(n446), .IN3(n474), .IN4(n446), .Q(n148) );
  XOR2X1 U547 ( .IN1(n445), .IN2(a[8]), .Q(n550) );
  NOR2X0 U548 ( .IN1(n414), .IN2(n521), .QN(n549) );
  XNOR2X1 U549 ( .IN1(a[8]), .IN2(n443), .Q(n521) );
  AO22X1 U550 ( .IN1(n551), .IN2(n447), .IN3(n477), .IN4(n447), .Q(n147) );
  XOR2X1 U551 ( .IN1(n447), .IN2(a[10]), .Q(n552) );
  NOR2X0 U552 ( .IN1(n414), .IN2(n532), .QN(n551) );
  XNOR2X1 U553 ( .IN1(a[10]), .IN2(n445), .Q(n532) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_8 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;
  wire   n1, n2;
  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_8_DW_mult_tc_0 mult_30 ( .a(in_a), .b({
        in_b[11:5], n2, in_b[3:0]}), .product(pre_out) );
  INVX0 U3 ( .INP(in_b[4]), .ZN(n1) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_2_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [24:0] carry;

  FADDX1 U2_22 ( .A(A[22]), .B(n7), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n8), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n9), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n10), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n11), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n12), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n13), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n18), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n21), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n22), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XNOR3X1 U1 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(DIFF[23]) );
  INVX0 U2 ( .INP(B[21]), .ZN(n8) );
  INVX0 U3 ( .INP(B[20]), .ZN(n9) );
  INVX0 U4 ( .INP(B[22]), .ZN(n7) );
  INVX0 U5 ( .INP(B[19]), .ZN(n10) );
  INVX0 U6 ( .INP(B[18]), .ZN(n11) );
  INVX0 U7 ( .INP(B[17]), .ZN(n12) );
  INVX0 U8 ( .INP(B[16]), .ZN(n13) );
  INVX0 U9 ( .INP(B[15]), .ZN(n14) );
  INVX0 U10 ( .INP(B[14]), .ZN(n15) );
  INVX0 U11 ( .INP(B[13]), .ZN(n16) );
  INVX0 U12 ( .INP(B[12]), .ZN(n17) );
  INVX0 U13 ( .INP(B[11]), .ZN(n18) );
  INVX0 U14 ( .INP(B[10]), .ZN(n19) );
  INVX0 U15 ( .INP(B[9]), .ZN(n20) );
  INVX0 U16 ( .INP(B[8]), .ZN(n21) );
  INVX0 U17 ( .INP(B[7]), .ZN(n22) );
  INVX0 U18 ( .INP(A[3]), .ZN(n4) );
  INVX0 U19 ( .INP(A[1]), .ZN(n6) );
  INVX0 U20 ( .INP(A[5]), .ZN(n2) );
  INVX0 U21 ( .INP(A[2]), .ZN(n5) );
  INVX0 U22 ( .INP(B[0]), .ZN(n23) );
  INVX0 U23 ( .INP(A[4]), .ZN(n3) );
  INVX0 U24 ( .INP(A[6]), .ZN(n1) );
  OAI22X1 U25 ( .IN1(n24), .IN2(n1), .IN3(B[6]), .IN4(n25), .QN(carry[7]) );
  AND2X1 U26 ( .IN1(n1), .IN2(n24), .Q(n25) );
  OA22X1 U27 ( .IN1(n26), .IN2(n2), .IN3(B[5]), .IN4(n27), .Q(n24) );
  AND2X1 U28 ( .IN1(n2), .IN2(n26), .Q(n27) );
  OA22X1 U29 ( .IN1(n28), .IN2(n3), .IN3(B[4]), .IN4(n29), .Q(n26) );
  AND2X1 U30 ( .IN1(n3), .IN2(n28), .Q(n29) );
  OA22X1 U31 ( .IN1(n30), .IN2(n4), .IN3(B[3]), .IN4(n31), .Q(n28) );
  AND2X1 U32 ( .IN1(n4), .IN2(n30), .Q(n31) );
  OA22X1 U33 ( .IN1(n32), .IN2(n5), .IN3(B[2]), .IN4(n33), .Q(n30) );
  AND2X1 U34 ( .IN1(n5), .IN2(n32), .Q(n33) );
  OA22X1 U35 ( .IN1(n34), .IN2(n6), .IN3(B[1]), .IN4(n35), .Q(n32) );
  AND2X1 U36 ( .IN1(n6), .IN2(n34), .Q(n35) );
  NOR2X0 U37 ( .IN1(n23), .IN2(A[0]), .QN(n34) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_2 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_2_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(\output ) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_2_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AO22X1 U1 ( .IN1(A[6]), .IN2(n1), .IN3(B[6]), .IN4(n2), .Q(carry[7]) );
  OR2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AO22X1 U3 ( .IN1(A[5]), .IN2(n3), .IN3(B[5]), .IN4(n4), .Q(n1) );
  OR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AO22X1 U5 ( .IN1(A[4]), .IN2(n5), .IN3(B[4]), .IN4(n6), .Q(n3) );
  OR2X1 U6 ( .IN1(n5), .IN2(A[4]), .Q(n6) );
  AO22X1 U7 ( .IN1(A[3]), .IN2(n7), .IN3(B[3]), .IN4(n8), .Q(n5) );
  OR2X1 U8 ( .IN1(n7), .IN2(A[3]), .Q(n8) );
  AO22X1 U9 ( .IN1(A[2]), .IN2(n9), .IN3(B[2]), .IN4(n10), .Q(n7) );
  OR2X1 U10 ( .IN1(n9), .IN2(A[2]), .Q(n10) );
  AO22X1 U11 ( .IN1(B[1]), .IN2(A[1]), .IN3(n11), .IN4(B[0]), .Q(n9) );
  OA21X1 U12 ( .IN1(A[1]), .IN2(B[1]), .IN3(A[0]), .Q(n11) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_2 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_2_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(\output ) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2 ( a_r, a_i, b_r, b_i, out_r, 
        out_i, clk );
  input [11:0] a_r;
  input [11:0] a_i;
  input [11:0] b_r;
  input [11:0] b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44;
  wire   [23:0] mult1_out;
  wire   [23:0] mult2_out;
  wire   [23:0] mult3_out;
  wire   [23:0] mult4_out;
  wire   [23:7] pre_out_r;
  wire   [23:7] pre_out_i;
  wire   [11:0] rnd_out_r;
  wire   [11:0] rnd_out_i;
  wire   [11:0] pos_out_r;
  wire   [11:0] pos_out_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFFX1 \out_r_reg_reg[11]  ( .D(pos_out_r[11]), .CLK(clk), .Q(out_r[11]) );
  DFFX1 \out_r_reg_reg[10]  ( .D(pos_out_r[10]), .CLK(clk), .Q(out_r[10]) );
  DFFX1 \out_r_reg_reg[9]  ( .D(pos_out_r[9]), .CLK(clk), .Q(out_r[9]) );
  DFFX1 \out_r_reg_reg[8]  ( .D(pos_out_r[8]), .CLK(clk), .Q(out_r[8]) );
  DFFX1 \out_r_reg_reg[7]  ( .D(pos_out_r[7]), .CLK(clk), .Q(out_r[7]) );
  DFFX1 \out_r_reg_reg[6]  ( .D(pos_out_r[6]), .CLK(clk), .Q(out_r[6]) );
  DFFX1 \out_r_reg_reg[5]  ( .D(pos_out_r[5]), .CLK(clk), .Q(out_r[5]) );
  DFFX1 \out_r_reg_reg[4]  ( .D(pos_out_r[4]), .CLK(clk), .Q(out_r[4]) );
  DFFX1 \out_r_reg_reg[3]  ( .D(pos_out_r[3]), .CLK(clk), .Q(out_r[3]) );
  DFFX1 \out_r_reg_reg[2]  ( .D(pos_out_r[2]), .CLK(clk), .Q(out_r[2]) );
  DFFX1 \out_r_reg_reg[1]  ( .D(pos_out_r[1]), .CLK(clk), .Q(out_r[1]) );
  DFFX1 \out_r_reg_reg[0]  ( .D(pos_out_r[0]), .CLK(clk), .Q(out_r[0]) );
  DFFX1 \out_i_reg_reg[11]  ( .D(pos_out_i[11]), .CLK(clk), .Q(out_i[11]) );
  DFFX1 \out_i_reg_reg[10]  ( .D(pos_out_i[10]), .CLK(clk), .Q(out_i[10]) );
  DFFX1 \out_i_reg_reg[9]  ( .D(pos_out_i[9]), .CLK(clk), .Q(out_i[9]) );
  DFFX1 \out_i_reg_reg[8]  ( .D(pos_out_i[8]), .CLK(clk), .Q(out_i[8]) );
  DFFX1 \out_i_reg_reg[7]  ( .D(pos_out_i[7]), .CLK(clk), .Q(out_i[7]) );
  DFFX1 \out_i_reg_reg[6]  ( .D(pos_out_i[6]), .CLK(clk), .Q(out_i[6]) );
  DFFX1 \out_i_reg_reg[5]  ( .D(pos_out_i[5]), .CLK(clk), .Q(out_i[5]) );
  DFFX1 \out_i_reg_reg[4]  ( .D(pos_out_i[4]), .CLK(clk), .Q(out_i[4]) );
  DFFX1 \out_i_reg_reg[3]  ( .D(pos_out_i[3]), .CLK(clk), .Q(out_i[3]) );
  DFFX1 \out_i_reg_reg[2]  ( .D(pos_out_i[2]), .CLK(clk), .Q(out_i[2]) );
  DFFX1 \out_i_reg_reg[1]  ( .D(pos_out_i[1]), .CLK(clk), .Q(out_i[1]) );
  DFFX1 \out_i_reg_reg[0]  ( .D(pos_out_i[0]), .CLK(clk), .Q(out_i[0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_11 mult1 ( .in_a({a_r[11:2], n14, a_r[0]}), 
        .in_b({b_r[11:8], n11, b_r[6:3], n12, b_r[1], n1}), .clk(clk), 
        .\output (mult1_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_10 mult2 ( .in_a({a_i[11:2], n13, a_i[0]}), 
        .in_b({b_i[11:8], n2, n4, b_i[5:2], n6, b_i[0]}), .clk(clk), 
        .\output (mult2_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_9 mult3 ( .in_a({a_r[11:2], n14, a_r[0]}), 
        .in_b({b_i[11:8], n2, n4, b_i[5:2], n6, b_i[0]}), .clk(clk), 
        .\output (mult3_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_8 mult4 ( .in_a({a_i[11:2], n13, a_i[0]}), 
        .in_b({b_r[11:8], n11, b_r[6:3], n12, b_r[1], n1}), .clk(clk), 
        .\output (mult4_out) );
  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_2 sub ( .a(mult1_out), .b(mult2_out), .\output ({pre_out_r, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_2 add ( .a(mult3_out), .b(mult4_out), .\output ({pre_out_i, SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_DW01_inc_0 add_154_round ( .A(
        pre_out_i[19:7]), .SUM({rnd_out_i, SYNOPSYS_UNCONNECTED__14}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2_DW01_inc_1 add_140_round ( .A(
        pre_out_r[19:7]), .SUM({rnd_out_r, SYNOPSYS_UNCONNECTED__15}) );
  DELLN2X2 U3 ( .INP(b_r[0]), .Z(n1) );
  DELLN1X2 U4 ( .INP(b_r[2]), .Z(n12) );
  DELLN2X2 U5 ( .INP(b_i[7]), .Z(n2) );
  INVX0 U6 ( .INP(b_i[6]), .ZN(n3) );
  INVX1 U7 ( .INP(n3), .ZN(n4) );
  INVX0 U8 ( .INP(b_i[1]), .ZN(n5) );
  INVX1 U9 ( .INP(n5), .ZN(n6) );
  INVX0 U10 ( .INP(pre_out_r[23]), .ZN(n37) );
  INVX0 U11 ( .INP(pre_out_i[23]), .ZN(n22) );
  INVX0 U12 ( .INP(n38), .ZN(n40) );
  INVX0 U13 ( .INP(n23), .ZN(n25) );
  AND2X1 U14 ( .IN1(n24), .IN2(n26), .Q(n7) );
  AND2X1 U15 ( .IN1(n39), .IN2(n41), .Q(n8) );
  AND2X1 U16 ( .IN1(n25), .IN2(n26), .Q(n9) );
  AND2X1 U17 ( .IN1(n40), .IN2(n41), .Q(n10) );
  NOR2X0 U18 ( .IN1(pre_out_r[21]), .IN2(pre_out_r[22]), .QN(n30) );
  NOR2X0 U19 ( .IN1(pre_out_i[21]), .IN2(pre_out_i[22]), .QN(n15) );
  NAND2X0 U20 ( .IN1(n31), .IN2(n30), .QN(n33) );
  NOR2X0 U21 ( .IN1(pre_out_r[19]), .IN2(pre_out_r[20]), .QN(n31) );
  NAND2X0 U22 ( .IN1(n16), .IN2(n15), .QN(n18) );
  NOR2X0 U23 ( .IN1(pre_out_i[19]), .IN2(pre_out_i[20]), .QN(n16) );
  INVX0 U24 ( .INP(n28), .ZN(n21) );
  INVX0 U25 ( .INP(n26), .ZN(n27) );
  INVX0 U26 ( .INP(n41), .ZN(n42) );
  INVX0 U27 ( .INP(n43), .ZN(n36) );
  DELLN1X2 U28 ( .INP(b_r[7]), .Z(n11) );
  XNOR2X1 U29 ( .IN1(mult3_out[23]), .IN2(mult4_out[23]), .Q(n20) );
  NAND2X0 U30 ( .IN1(n35), .IN2(n34), .QN(n43) );
  DELLN1X2 U31 ( .INP(a_i[1]), .Z(n13) );
  DELLN1X2 U32 ( .INP(a_r[1]), .Z(n14) );
  NAND4X0 U33 ( .IN1(pre_out_i[22]), .IN2(pre_out_i[21]), .IN3(pre_out_i[20]), 
        .IN4(pre_out_i[19]), .QN(n17) );
  MUX21X1 U34 ( .IN1(n18), .IN2(n17), .S(pre_out_i[23]), .Q(n23) );
  XOR2X1 U35 ( .IN1(pre_out_i[23]), .IN2(mult3_out[23]), .Q(n19) );
  NAND2X1 U36 ( .IN1(n20), .IN2(n19), .QN(n28) );
  NAND2X1 U37 ( .IN1(mult3_out[23]), .IN2(n21), .QN(n26) );
  AO21X1 U38 ( .IN1(n23), .IN2(n22), .IN3(n21), .Q(n24) );
  AO21X1 U39 ( .IN1(rnd_out_i[0]), .IN2(n9), .IN3(n7), .Q(pos_out_i[0]) );
  AO21X1 U40 ( .IN1(rnd_out_i[1]), .IN2(n9), .IN3(n7), .Q(pos_out_i[1]) );
  AO21X1 U41 ( .IN1(rnd_out_i[2]), .IN2(n9), .IN3(n7), .Q(pos_out_i[2]) );
  AO21X1 U42 ( .IN1(rnd_out_i[3]), .IN2(n9), .IN3(n7), .Q(pos_out_i[3]) );
  AO21X1 U43 ( .IN1(rnd_out_i[4]), .IN2(n9), .IN3(n7), .Q(pos_out_i[4]) );
  AO21X1 U44 ( .IN1(rnd_out_i[5]), .IN2(n9), .IN3(n7), .Q(pos_out_i[5]) );
  AO21X1 U45 ( .IN1(rnd_out_i[6]), .IN2(n9), .IN3(n7), .Q(pos_out_i[6]) );
  AO21X1 U46 ( .IN1(rnd_out_i[7]), .IN2(n9), .IN3(n7), .Q(pos_out_i[7]) );
  AO21X1 U47 ( .IN1(rnd_out_i[8]), .IN2(n9), .IN3(n7), .Q(pos_out_i[8]) );
  AO21X1 U48 ( .IN1(rnd_out_i[9]), .IN2(n9), .IN3(n7), .Q(pos_out_i[9]) );
  AO21X1 U49 ( .IN1(rnd_out_i[10]), .IN2(n9), .IN3(n7), .Q(pos_out_i[10]) );
  MUX21X1 U50 ( .IN1(pre_out_i[23]), .IN2(rnd_out_i[11]), .S(n25), .Q(n29) );
  AO21X1 U51 ( .IN1(n29), .IN2(n28), .IN3(n27), .Q(pos_out_i[11]) );
  NAND4X0 U52 ( .IN1(pre_out_r[22]), .IN2(pre_out_r[21]), .IN3(pre_out_r[20]), 
        .IN4(pre_out_r[19]), .QN(n32) );
  MUX21X1 U53 ( .IN1(n33), .IN2(n32), .S(pre_out_r[23]), .Q(n38) );
  XOR2X1 U54 ( .IN1(mult2_out[23]), .IN2(mult1_out[23]), .Q(n35) );
  XOR2X1 U55 ( .IN1(pre_out_r[23]), .IN2(mult1_out[23]), .Q(n34) );
  NAND2X1 U56 ( .IN1(mult1_out[23]), .IN2(n36), .QN(n41) );
  AO21X1 U57 ( .IN1(n38), .IN2(n37), .IN3(n36), .Q(n39) );
  AO21X1 U58 ( .IN1(rnd_out_r[0]), .IN2(n10), .IN3(n8), .Q(pos_out_r[0]) );
  AO21X1 U59 ( .IN1(rnd_out_r[1]), .IN2(n10), .IN3(n8), .Q(pos_out_r[1]) );
  AO21X1 U60 ( .IN1(rnd_out_r[2]), .IN2(n10), .IN3(n8), .Q(pos_out_r[2]) );
  AO21X1 U61 ( .IN1(rnd_out_r[3]), .IN2(n10), .IN3(n8), .Q(pos_out_r[3]) );
  AO21X1 U62 ( .IN1(rnd_out_r[4]), .IN2(n10), .IN3(n8), .Q(pos_out_r[4]) );
  AO21X1 U63 ( .IN1(rnd_out_r[5]), .IN2(n10), .IN3(n8), .Q(pos_out_r[5]) );
  AO21X1 U64 ( .IN1(rnd_out_r[6]), .IN2(n10), .IN3(n8), .Q(pos_out_r[6]) );
  AO21X1 U65 ( .IN1(rnd_out_r[7]), .IN2(n10), .IN3(n8), .Q(pos_out_r[7]) );
  AO21X1 U66 ( .IN1(rnd_out_r[8]), .IN2(n10), .IN3(n8), .Q(pos_out_r[8]) );
  AO21X1 U67 ( .IN1(rnd_out_r[9]), .IN2(n10), .IN3(n8), .Q(pos_out_r[9]) );
  AO21X1 U68 ( .IN1(rnd_out_r[10]), .IN2(n10), .IN3(n8), .Q(pos_out_r[10]) );
  MUX21X1 U69 ( .IN1(pre_out_r[23]), .IN2(rnd_out_r[11]), .S(n40), .Q(n44) );
  AO21X1 U70 ( .IN1(n44), .IN2(n43), .IN3(n42), .Q(pos_out_r[11]) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_7_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n452), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n454), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n456), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n458), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n460), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  FADDX1 U311 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U312 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  XOR2X2 U313 ( .IN1(n437), .IN2(n450), .Q(n537) );
  XOR2X2 U314 ( .IN1(n437), .IN2(n448), .Q(n526) );
  XOR2X2 U315 ( .IN1(n437), .IN2(n446), .Q(n515) );
  XOR2X2 U316 ( .IN1(n437), .IN2(n444), .Q(n504) );
  INVX0 U317 ( .INP(b[2]), .ZN(n408) );
  INVX0 U318 ( .INP(n408), .ZN(n409) );
  DELLN2X2 U319 ( .INP(n15), .Z(n410) );
  INVX0 U320 ( .INP(b[1]), .ZN(n411) );
  INVX0 U321 ( .INP(n411), .ZN(n412) );
  DELLN2X2 U322 ( .INP(n7), .Z(n413) );
  DELLN2X2 U323 ( .INP(n11), .Z(n414) );
  XOR2X2 U324 ( .IN1(n409), .IN2(n450), .Q(n538) );
  XOR2X2 U325 ( .IN1(n409), .IN2(n448), .Q(n527) );
  XOR2X2 U326 ( .IN1(n409), .IN2(n446), .Q(n516) );
  XOR2X2 U327 ( .IN1(n409), .IN2(n444), .Q(n505) );
  XOR2X2 U328 ( .IN1(n409), .IN2(n442), .Q(n495) );
  XOR2X2 U329 ( .IN1(n409), .IN2(n436), .Q(n483) );
  XOR2X2 U330 ( .IN1(b[8]), .IN2(n450), .Q(n544) );
  XOR2X2 U331 ( .IN1(b[8]), .IN2(n448), .Q(n533) );
  XOR2X2 U332 ( .IN1(b[8]), .IN2(n446), .Q(n522) );
  XOR2X2 U333 ( .IN1(b[8]), .IN2(n444), .Q(n511) );
  XOR2X2 U334 ( .IN1(b[8]), .IN2(n442), .Q(n501) );
  XOR2X2 U335 ( .IN1(b[8]), .IN2(n436), .Q(n489) );
  XOR3X2 U336 ( .IN1(n65), .IN2(n58), .IN3(n12), .Q(product[14]) );
  NAND2X0 U337 ( .IN1(n65), .IN2(n58), .QN(n415) );
  NAND2X0 U338 ( .IN1(n65), .IN2(n12), .QN(n416) );
  NAND2X0 U339 ( .IN1(n58), .IN2(n12), .QN(n417) );
  NAND3X0 U340 ( .IN1(n415), .IN2(n416), .IN3(n417), .QN(n11) );
  XOR2X1 U341 ( .IN1(n57), .IN2(n50), .Q(n418) );
  XOR2X1 U342 ( .IN1(n418), .IN2(n414), .Q(product[15]) );
  NAND2X0 U343 ( .IN1(n57), .IN2(n50), .QN(n419) );
  NAND2X0 U344 ( .IN1(n57), .IN2(n11), .QN(n420) );
  NAND2X0 U345 ( .IN1(n50), .IN2(n11), .QN(n421) );
  NAND3X0 U346 ( .IN1(n421), .IN2(n420), .IN3(n419), .QN(n10) );
  XOR2X2 U347 ( .IN1(b[6]), .IN2(n450), .Q(n542) );
  XOR2X2 U348 ( .IN1(b[6]), .IN2(n448), .Q(n531) );
  XOR2X2 U349 ( .IN1(b[6]), .IN2(n446), .Q(n520) );
  XOR2X2 U350 ( .IN1(b[6]), .IN2(n444), .Q(n509) );
  XOR2X2 U351 ( .IN1(b[6]), .IN2(n442), .Q(n499) );
  XOR2X2 U352 ( .IN1(b[6]), .IN2(n436), .Q(n487) );
  XOR2X2 U353 ( .IN1(b[4]), .IN2(n450), .Q(n540) );
  XOR2X2 U354 ( .IN1(b[4]), .IN2(n448), .Q(n529) );
  XOR2X2 U355 ( .IN1(b[4]), .IN2(n446), .Q(n518) );
  XOR2X2 U356 ( .IN1(b[4]), .IN2(n444), .Q(n507) );
  XOR2X2 U357 ( .IN1(b[4]), .IN2(n442), .Q(n497) );
  XOR2X2 U358 ( .IN1(b[4]), .IN2(n436), .Q(n485) );
  XOR2X2 U359 ( .IN1(b[3]), .IN2(n450), .Q(n539) );
  XOR2X2 U360 ( .IN1(b[3]), .IN2(n448), .Q(n528) );
  XOR2X2 U361 ( .IN1(b[3]), .IN2(n446), .Q(n517) );
  XOR2X2 U362 ( .IN1(b[3]), .IN2(n444), .Q(n506) );
  XOR2X2 U363 ( .IN1(b[3]), .IN2(n442), .Q(n496) );
  XOR2X2 U364 ( .IN1(b[3]), .IN2(n436), .Q(n484) );
  XOR2X2 U365 ( .IN1(b[5]), .IN2(n450), .Q(n541) );
  XOR2X2 U366 ( .IN1(b[5]), .IN2(n448), .Q(n530) );
  XOR2X2 U367 ( .IN1(b[5]), .IN2(n446), .Q(n519) );
  XOR2X2 U368 ( .IN1(b[5]), .IN2(n444), .Q(n508) );
  XOR2X2 U369 ( .IN1(b[5]), .IN2(n442), .Q(n498) );
  XOR2X2 U370 ( .IN1(b[5]), .IN2(n436), .Q(n486) );
  XOR2X2 U371 ( .IN1(n412), .IN2(n450), .Q(n536) );
  XOR2X2 U372 ( .IN1(n412), .IN2(n448), .Q(n525) );
  XOR2X2 U373 ( .IN1(n412), .IN2(n446), .Q(n514) );
  XOR2X2 U374 ( .IN1(n412), .IN2(n444), .Q(n503) );
  XOR2X2 U375 ( .IN1(n412), .IN2(n442), .Q(n493) );
  XOR2X2 U376 ( .IN1(n412), .IN2(n436), .Q(n482) );
  XOR3X1 U377 ( .IN1(n37), .IN2(n34), .IN3(n8), .Q(product[18]) );
  XOR3X1 U378 ( .IN1(n96), .IN2(n103), .IN3(n16), .Q(product[10]) );
  XNOR2X1 U379 ( .IN1(n422), .IN2(n410), .Q(product[11]) );
  XNOR2X1 U380 ( .IN1(n86), .IN2(n95), .Q(n422) );
  INVX0 U381 ( .INP(n25), .ZN(n452) );
  INVX0 U382 ( .INP(n3), .ZN(product[23]) );
  INVX0 U383 ( .INP(n55), .ZN(n458) );
  XNOR2X1 U384 ( .IN1(n413), .IN2(n423), .Q(product[19]) );
  XNOR2X1 U385 ( .IN1(n33), .IN2(n30), .Q(n423) );
  INVX0 U386 ( .INP(n73), .ZN(n460) );
  FADDX1 U387 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U388 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  INVX0 U389 ( .INP(n41), .ZN(n456) );
  INVX0 U390 ( .INP(n31), .ZN(n454) );
  NBUFFX2 U391 ( .INP(a[1]), .Z(n436) );
  INVX0 U392 ( .INP(n492), .ZN(n461) );
  AND2X1 U393 ( .IN1(n436), .IN2(n441), .Q(n467) );
  INVX0 U394 ( .INP(n502), .ZN(n459) );
  INVX0 U395 ( .INP(n513), .ZN(n457) );
  INVX0 U396 ( .INP(n524), .ZN(n455) );
  INVX0 U397 ( .INP(n535), .ZN(n453) );
  NBUFFX2 U398 ( .INP(a[5]), .Z(n445) );
  NBUFFX2 U399 ( .INP(a[3]), .Z(n443) );
  XOR2X1 U400 ( .IN1(b[7]), .IN2(n436), .Q(n488) );
  AND2X1 U401 ( .IN1(n492), .IN2(n547), .Q(n465) );
  AND2X1 U402 ( .IN1(n513), .IN2(n551), .Q(n474) );
  AND2X1 U403 ( .IN1(n502), .IN2(n549), .Q(n471) );
  AND2X1 U404 ( .IN1(n524), .IN2(n553), .Q(n477) );
  AND2X1 U405 ( .IN1(n535), .IN2(n555), .Q(n480) );
  NBUFFX2 U406 ( .INP(a[7]), .Z(n447) );
  NBUFFX2 U407 ( .INP(a[9]), .Z(n449) );
  NAND2X0 U408 ( .IN1(n37), .IN2(n34), .QN(n424) );
  NAND2X0 U409 ( .IN1(n37), .IN2(n8), .QN(n425) );
  NAND2X0 U410 ( .IN1(n34), .IN2(n8), .QN(n426) );
  NAND3X0 U411 ( .IN1(n424), .IN2(n425), .IN3(n426), .QN(n7) );
  NAND2X0 U412 ( .IN1(n33), .IN2(n30), .QN(n427) );
  NAND2X0 U413 ( .IN1(n33), .IN2(n7), .QN(n428) );
  NAND2X0 U414 ( .IN1(n30), .IN2(n7), .QN(n429) );
  NAND3X0 U415 ( .IN1(n429), .IN2(n428), .IN3(n427), .QN(n6) );
  NAND2X0 U416 ( .IN1(n96), .IN2(n103), .QN(n430) );
  NAND2X0 U417 ( .IN1(n96), .IN2(n16), .QN(n431) );
  NAND2X0 U418 ( .IN1(n103), .IN2(n16), .QN(n432) );
  NAND3X0 U419 ( .IN1(n432), .IN2(n431), .IN3(n430), .QN(n15) );
  NAND2X0 U420 ( .IN1(n86), .IN2(n95), .QN(n433) );
  NAND2X0 U421 ( .IN1(n86), .IN2(n15), .QN(n434) );
  NAND2X0 U422 ( .IN1(n95), .IN2(n15), .QN(n435) );
  NAND3X0 U423 ( .IN1(n435), .IN2(n434), .IN3(n433), .QN(n14) );
  DELLN1X2 U424 ( .INP(a[11]), .Z(n450) );
  INVX0 U425 ( .INP(n439), .ZN(n437) );
  INVX0 U426 ( .INP(b[0]), .ZN(n438) );
  INVX0 U427 ( .INP(b[0]), .ZN(n439) );
  INVX0 U428 ( .INP(n441), .ZN(n440) );
  INVX0 U429 ( .INP(a[0]), .ZN(n441) );
  DELLN1X2 U430 ( .INP(a[3]), .Z(n442) );
  DELLN1X2 U431 ( .INP(a[5]), .Z(n444) );
  DELLN1X2 U432 ( .INP(a[7]), .Z(n446) );
  DELLN1X2 U433 ( .INP(a[9]), .Z(n448) );
  NOR2X0 U434 ( .IN1(n441), .IN2(n438), .QN(product[0]) );
  XNOR2X1 U435 ( .IN1(n462), .IN2(n463), .Q(n84) );
  NAND2X0 U436 ( .IN1(n463), .IN2(n462), .QN(n83) );
  AOI22X1 U437 ( .IN1(n464), .IN2(n461), .IN3(n465), .IN4(n466), .QN(n462) );
  OA21X1 U438 ( .IN1(n467), .IN2(n440), .IN3(n468), .Q(n463) );
  AO22X1 U439 ( .IN1(n469), .IN2(n461), .IN3(n465), .IN4(n464), .Q(n73) );
  XOR2X1 U440 ( .IN1(b[10]), .IN2(n442), .Q(n464) );
  AO22X1 U441 ( .IN1(n470), .IN2(n459), .IN3(n471), .IN4(n472), .Q(n55) );
  AO22X1 U442 ( .IN1(n473), .IN2(n457), .IN3(n474), .IN4(n475), .Q(n41) );
  AO22X1 U443 ( .IN1(n476), .IN2(n455), .IN3(n477), .IN4(n478), .Q(n31) );
  AO22X1 U444 ( .IN1(n479), .IN2(n453), .IN3(n480), .IN4(n481), .Q(n25) );
  AO22X1 U445 ( .IN1(n440), .IN2(n482), .IN3(n467), .IN4(n439), .Q(n224) );
  AO22X1 U446 ( .IN1(n440), .IN2(n483), .IN3(n467), .IN4(n482), .Q(n223) );
  AO22X1 U447 ( .IN1(n440), .IN2(n484), .IN3(n467), .IN4(n483), .Q(n222) );
  AO22X1 U448 ( .IN1(n440), .IN2(n485), .IN3(n467), .IN4(n484), .Q(n221) );
  AO22X1 U449 ( .IN1(n440), .IN2(n486), .IN3(n467), .IN4(n485), .Q(n220) );
  AO22X1 U450 ( .IN1(n440), .IN2(n487), .IN3(n467), .IN4(n486), .Q(n219) );
  AO22X1 U451 ( .IN1(n440), .IN2(n488), .IN3(n467), .IN4(n487), .Q(n218) );
  AO22X1 U452 ( .IN1(n440), .IN2(n489), .IN3(n467), .IN4(n488), .Q(n217) );
  AO22X1 U453 ( .IN1(n440), .IN2(n490), .IN3(n467), .IN4(n489), .Q(n216) );
  AO22X1 U454 ( .IN1(n440), .IN2(n491), .IN3(n467), .IN4(n490), .Q(n215) );
  XOR2X1 U455 ( .IN1(b[9]), .IN2(n436), .Q(n490) );
  AO22X1 U456 ( .IN1(n440), .IN2(n468), .IN3(n467), .IN4(n491), .Q(n214) );
  XOR2X1 U457 ( .IN1(b[10]), .IN2(n436), .Q(n491) );
  XOR2X1 U458 ( .IN1(b[11]), .IN2(n436), .Q(n468) );
  NOR2X0 U459 ( .IN1(n492), .IN2(n438), .QN(n212) );
  AO22X1 U460 ( .IN1(n493), .IN2(n461), .IN3(n465), .IN4(n494), .Q(n211) );
  XOR2X1 U461 ( .IN1(n437), .IN2(n442), .Q(n494) );
  AO22X1 U462 ( .IN1(n495), .IN2(n461), .IN3(n465), .IN4(n493), .Q(n210) );
  AO22X1 U463 ( .IN1(n496), .IN2(n461), .IN3(n465), .IN4(n495), .Q(n209) );
  AO22X1 U464 ( .IN1(n497), .IN2(n461), .IN3(n465), .IN4(n496), .Q(n208) );
  AO22X1 U465 ( .IN1(n498), .IN2(n461), .IN3(n465), .IN4(n497), .Q(n207) );
  AO22X1 U466 ( .IN1(n499), .IN2(n461), .IN3(n465), .IN4(n498), .Q(n206) );
  AO22X1 U467 ( .IN1(n500), .IN2(n461), .IN3(n465), .IN4(n499), .Q(n205) );
  AO22X1 U468 ( .IN1(n501), .IN2(n461), .IN3(n465), .IN4(n500), .Q(n204) );
  XOR2X1 U469 ( .IN1(b[7]), .IN2(n442), .Q(n500) );
  AO22X1 U470 ( .IN1(n466), .IN2(n461), .IN3(n465), .IN4(n501), .Q(n203) );
  XOR2X1 U471 ( .IN1(b[9]), .IN2(n442), .Q(n466) );
  OAI21X1 U472 ( .IN1(n461), .IN2(n465), .IN3(n469), .QN(n201) );
  XOR2X1 U473 ( .IN1(b[11]), .IN2(n442), .Q(n469) );
  NOR2X0 U474 ( .IN1(n502), .IN2(n438), .QN(n200) );
  AO22X1 U475 ( .IN1(n503), .IN2(n459), .IN3(n471), .IN4(n504), .Q(n199) );
  AO22X1 U476 ( .IN1(n505), .IN2(n459), .IN3(n471), .IN4(n503), .Q(n198) );
  AO22X1 U477 ( .IN1(n506), .IN2(n459), .IN3(n471), .IN4(n505), .Q(n197) );
  AO22X1 U478 ( .IN1(n507), .IN2(n459), .IN3(n471), .IN4(n506), .Q(n196) );
  AO22X1 U479 ( .IN1(n508), .IN2(n459), .IN3(n471), .IN4(n507), .Q(n195) );
  AO22X1 U480 ( .IN1(n509), .IN2(n459), .IN3(n471), .IN4(n508), .Q(n194) );
  AO22X1 U481 ( .IN1(n510), .IN2(n459), .IN3(n471), .IN4(n509), .Q(n193) );
  AO22X1 U482 ( .IN1(n511), .IN2(n459), .IN3(n471), .IN4(n510), .Q(n192) );
  XOR2X1 U483 ( .IN1(b[7]), .IN2(n444), .Q(n510) );
  AO22X1 U484 ( .IN1(n512), .IN2(n459), .IN3(n471), .IN4(n511), .Q(n191) );
  AO22X1 U485 ( .IN1(n472), .IN2(n459), .IN3(n471), .IN4(n512), .Q(n190) );
  XOR2X1 U486 ( .IN1(b[9]), .IN2(n444), .Q(n512) );
  XOR2X1 U487 ( .IN1(b[10]), .IN2(n444), .Q(n472) );
  OAI21X1 U488 ( .IN1(n459), .IN2(n471), .IN3(n470), .QN(n189) );
  XOR2X1 U489 ( .IN1(b[11]), .IN2(n444), .Q(n470) );
  NOR2X0 U490 ( .IN1(n513), .IN2(n438), .QN(n188) );
  AO22X1 U491 ( .IN1(n514), .IN2(n457), .IN3(n474), .IN4(n515), .Q(n187) );
  AO22X1 U492 ( .IN1(n516), .IN2(n457), .IN3(n474), .IN4(n514), .Q(n186) );
  AO22X1 U493 ( .IN1(n517), .IN2(n457), .IN3(n474), .IN4(n516), .Q(n185) );
  AO22X1 U494 ( .IN1(n518), .IN2(n457), .IN3(n474), .IN4(n517), .Q(n184) );
  AO22X1 U495 ( .IN1(n519), .IN2(n457), .IN3(n474), .IN4(n518), .Q(n183) );
  AO22X1 U496 ( .IN1(n520), .IN2(n457), .IN3(n474), .IN4(n519), .Q(n182) );
  AO22X1 U497 ( .IN1(n521), .IN2(n457), .IN3(n474), .IN4(n520), .Q(n181) );
  AO22X1 U498 ( .IN1(n522), .IN2(n457), .IN3(n474), .IN4(n521), .Q(n180) );
  XOR2X1 U499 ( .IN1(b[7]), .IN2(n446), .Q(n521) );
  AO22X1 U500 ( .IN1(n523), .IN2(n457), .IN3(n474), .IN4(n522), .Q(n179) );
  AO22X1 U501 ( .IN1(n475), .IN2(n457), .IN3(n474), .IN4(n523), .Q(n178) );
  XOR2X1 U502 ( .IN1(b[9]), .IN2(n446), .Q(n523) );
  XOR2X1 U503 ( .IN1(b[10]), .IN2(n446), .Q(n475) );
  OAI21X1 U504 ( .IN1(n457), .IN2(n474), .IN3(n473), .QN(n177) );
  XOR2X1 U505 ( .IN1(b[11]), .IN2(n446), .Q(n473) );
  NOR2X0 U506 ( .IN1(n524), .IN2(n438), .QN(n176) );
  AO22X1 U507 ( .IN1(n525), .IN2(n455), .IN3(n477), .IN4(n526), .Q(n175) );
  AO22X1 U508 ( .IN1(n527), .IN2(n455), .IN3(n477), .IN4(n525), .Q(n174) );
  AO22X1 U509 ( .IN1(n528), .IN2(n455), .IN3(n477), .IN4(n527), .Q(n173) );
  AO22X1 U510 ( .IN1(n529), .IN2(n455), .IN3(n477), .IN4(n528), .Q(n172) );
  AO22X1 U511 ( .IN1(n530), .IN2(n455), .IN3(n477), .IN4(n529), .Q(n171) );
  AO22X1 U512 ( .IN1(n531), .IN2(n455), .IN3(n477), .IN4(n530), .Q(n170) );
  AO22X1 U513 ( .IN1(n532), .IN2(n455), .IN3(n477), .IN4(n531), .Q(n169) );
  AO22X1 U514 ( .IN1(n533), .IN2(n455), .IN3(n477), .IN4(n532), .Q(n168) );
  XOR2X1 U515 ( .IN1(b[7]), .IN2(n448), .Q(n532) );
  AO22X1 U516 ( .IN1(n534), .IN2(n455), .IN3(n477), .IN4(n533), .Q(n167) );
  AO22X1 U517 ( .IN1(n478), .IN2(n455), .IN3(n477), .IN4(n534), .Q(n166) );
  XOR2X1 U518 ( .IN1(b[9]), .IN2(n448), .Q(n534) );
  XOR2X1 U519 ( .IN1(b[10]), .IN2(n448), .Q(n478) );
  OAI21X1 U520 ( .IN1(n455), .IN2(n477), .IN3(n476), .QN(n165) );
  XOR2X1 U521 ( .IN1(b[11]), .IN2(n448), .Q(n476) );
  NOR2X0 U522 ( .IN1(n535), .IN2(n438), .QN(n164) );
  AO22X1 U523 ( .IN1(n536), .IN2(n453), .IN3(n480), .IN4(n537), .Q(n163) );
  AO22X1 U524 ( .IN1(n538), .IN2(n453), .IN3(n480), .IN4(n536), .Q(n162) );
  AO22X1 U525 ( .IN1(n539), .IN2(n453), .IN3(n480), .IN4(n538), .Q(n161) );
  AO22X1 U526 ( .IN1(n540), .IN2(n453), .IN3(n480), .IN4(n539), .Q(n160) );
  AO22X1 U527 ( .IN1(n541), .IN2(n453), .IN3(n480), .IN4(n540), .Q(n159) );
  AO22X1 U528 ( .IN1(n542), .IN2(n453), .IN3(n480), .IN4(n541), .Q(n158) );
  AO22X1 U529 ( .IN1(n543), .IN2(n453), .IN3(n480), .IN4(n542), .Q(n157) );
  AO22X1 U530 ( .IN1(n544), .IN2(n453), .IN3(n480), .IN4(n543), .Q(n156) );
  XOR2X1 U531 ( .IN1(b[7]), .IN2(n450), .Q(n543) );
  AO22X1 U532 ( .IN1(n545), .IN2(n453), .IN3(n480), .IN4(n544), .Q(n155) );
  AO22X1 U533 ( .IN1(n481), .IN2(n453), .IN3(n480), .IN4(n545), .Q(n154) );
  XOR2X1 U534 ( .IN1(b[9]), .IN2(n450), .Q(n545) );
  XOR2X1 U535 ( .IN1(b[10]), .IN2(n450), .Q(n481) );
  OAI21X1 U536 ( .IN1(n453), .IN2(n480), .IN3(n479), .QN(n153) );
  XOR2X1 U537 ( .IN1(b[11]), .IN2(n450), .Q(n479) );
  AO21X1 U538 ( .IN1(n436), .IN2(n439), .IN3(n467), .Q(n152) );
  AO22X1 U539 ( .IN1(n546), .IN2(n443), .IN3(n465), .IN4(n443), .Q(n151) );
  XOR2X1 U540 ( .IN1(n442), .IN2(a[2]), .Q(n547) );
  NOR2X0 U541 ( .IN1(n437), .IN2(n492), .QN(n546) );
  XNOR2X1 U542 ( .IN1(a[2]), .IN2(n436), .Q(n492) );
  AO22X1 U543 ( .IN1(n548), .IN2(n445), .IN3(n471), .IN4(n445), .Q(n150) );
  XOR2X1 U544 ( .IN1(n444), .IN2(a[4]), .Q(n549) );
  NOR2X0 U545 ( .IN1(n437), .IN2(n502), .QN(n548) );
  XNOR2X1 U546 ( .IN1(a[4]), .IN2(n442), .Q(n502) );
  AO22X1 U547 ( .IN1(n550), .IN2(n447), .IN3(n474), .IN4(n447), .Q(n149) );
  XOR2X1 U548 ( .IN1(n446), .IN2(a[6]), .Q(n551) );
  NOR2X0 U549 ( .IN1(n437), .IN2(n513), .QN(n550) );
  XNOR2X1 U550 ( .IN1(a[6]), .IN2(n444), .Q(n513) );
  AO22X1 U551 ( .IN1(n552), .IN2(n449), .IN3(n477), .IN4(n449), .Q(n148) );
  XOR2X1 U552 ( .IN1(n448), .IN2(a[8]), .Q(n553) );
  NOR2X0 U553 ( .IN1(n437), .IN2(n524), .QN(n552) );
  XNOR2X1 U554 ( .IN1(a[8]), .IN2(n446), .Q(n524) );
  AO22X1 U555 ( .IN1(n554), .IN2(n450), .IN3(n480), .IN4(n450), .Q(n147) );
  XOR2X1 U556 ( .IN1(n450), .IN2(a[10]), .Q(n555) );
  NOR2X0 U557 ( .IN1(n437), .IN2(n535), .QN(n554) );
  XNOR2X1 U558 ( .IN1(a[10]), .IN2(n448), .Q(n535) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_7 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_7_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_6_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n459), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n461), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n463), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n465), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n467), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  FADDX1 U311 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U312 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  XOR2X2 U313 ( .IN1(n445), .IN2(n457), .Q(n544) );
  XOR2X2 U314 ( .IN1(n445), .IN2(n455), .Q(n533) );
  XOR2X2 U315 ( .IN1(n445), .IN2(n453), .Q(n522) );
  XOR2X2 U316 ( .IN1(n445), .IN2(n451), .Q(n511) );
  INVX0 U317 ( .INP(b[3]), .ZN(n408) );
  INVX0 U318 ( .INP(n408), .ZN(n409) );
  INVX0 U319 ( .INP(b[1]), .ZN(n410) );
  INVX0 U320 ( .INP(n410), .ZN(n411) );
  XOR3X2 U321 ( .IN1(n124), .IN2(n127), .IN3(n20), .Q(product[6]) );
  NAND2X0 U322 ( .IN1(n124), .IN2(n127), .QN(n412) );
  NAND2X0 U323 ( .IN1(n124), .IN2(n20), .QN(n413) );
  NAND2X0 U324 ( .IN1(n127), .IN2(n20), .QN(n414) );
  NAND3X0 U325 ( .IN1(n412), .IN2(n413), .IN3(n414), .QN(n19) );
  XOR2X1 U326 ( .IN1(n118), .IN2(n123), .Q(n415) );
  XOR2X1 U327 ( .IN1(n415), .IN2(n19), .Q(product[7]) );
  NAND2X0 U328 ( .IN1(n118), .IN2(n123), .QN(n416) );
  NAND2X0 U329 ( .IN1(n118), .IN2(n19), .QN(n417) );
  NAND2X0 U330 ( .IN1(n123), .IN2(n19), .QN(n418) );
  NAND3X0 U331 ( .IN1(n416), .IN2(n417), .IN3(n418), .QN(n18) );
  INVX0 U332 ( .INP(n14), .ZN(n419) );
  INVX0 U333 ( .INP(n419), .ZN(n420) );
  XOR2X2 U334 ( .IN1(b[4]), .IN2(n457), .Q(n547) );
  XOR2X2 U335 ( .IN1(b[4]), .IN2(n455), .Q(n536) );
  XOR2X2 U336 ( .IN1(b[4]), .IN2(n453), .Q(n525) );
  XOR2X2 U337 ( .IN1(b[4]), .IN2(n451), .Q(n514) );
  XOR2X2 U338 ( .IN1(b[4]), .IN2(n449), .Q(n504) );
  XOR2X2 U339 ( .IN1(b[4]), .IN2(n444), .Q(n492) );
  XOR2X2 U340 ( .IN1(n409), .IN2(n457), .Q(n546) );
  XOR2X2 U341 ( .IN1(n409), .IN2(n455), .Q(n535) );
  XOR2X2 U342 ( .IN1(n409), .IN2(n453), .Q(n524) );
  XOR2X2 U343 ( .IN1(n409), .IN2(n451), .Q(n513) );
  XOR2X2 U344 ( .IN1(n409), .IN2(n449), .Q(n503) );
  XOR2X2 U345 ( .IN1(n409), .IN2(n444), .Q(n491) );
  XNOR2X1 U346 ( .IN1(n421), .IN2(n420), .Q(product[12]) );
  NAND2X0 U347 ( .IN1(n221), .IN2(n200), .QN(n437) );
  XOR3X1 U348 ( .IN1(n37), .IN2(n34), .IN3(n8), .Q(product[18]) );
  XOR3X1 U349 ( .IN1(n86), .IN2(n95), .IN3(n15), .Q(product[11]) );
  XNOR2X1 U350 ( .IN1(n76), .IN2(n85), .Q(n421) );
  INVX0 U351 ( .INP(n25), .ZN(n459) );
  INVX0 U352 ( .INP(n3), .ZN(product[23]) );
  INVX0 U353 ( .INP(n55), .ZN(n465) );
  XNOR2X1 U354 ( .IN1(n7), .IN2(n422), .Q(product[19]) );
  XNOR2X1 U355 ( .IN1(n33), .IN2(n30), .Q(n422) );
  XOR2X1 U356 ( .IN1(n443), .IN2(n444), .Q(n490) );
  XOR2X1 U357 ( .IN1(n411), .IN2(n444), .Q(n489) );
  XOR2X1 U358 ( .IN1(n411), .IN2(n449), .Q(n500) );
  XOR2X1 U359 ( .IN1(n411), .IN2(n451), .Q(n510) );
  XOR2X1 U360 ( .IN1(n411), .IN2(n453), .Q(n521) );
  INVX0 U361 ( .INP(n73), .ZN(n467) );
  FADDX1 U362 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X1 U363 ( .IN1(n411), .IN2(n455), .Q(n532) );
  XOR2X1 U364 ( .IN1(n411), .IN2(n457), .Q(n543) );
  INVX0 U365 ( .INP(n41), .ZN(n463) );
  INVX0 U366 ( .INP(n31), .ZN(n461) );
  NBUFFX2 U367 ( .INP(b[7]), .Z(n430) );
  NBUFFX2 U368 ( .INP(b[2]), .Z(n443) );
  NBUFFX2 U369 ( .INP(a[1]), .Z(n444) );
  INVX0 U370 ( .INP(n499), .ZN(n468) );
  AND2X1 U371 ( .IN1(n444), .IN2(n448), .Q(n474) );
  XOR2X1 U372 ( .IN1(b[6]), .IN2(n444), .Q(n494) );
  INVX0 U373 ( .INP(n509), .ZN(n466) );
  INVX0 U374 ( .INP(n520), .ZN(n464) );
  INVX0 U375 ( .INP(n531), .ZN(n462) );
  XNOR2X1 U376 ( .IN1(n423), .IN2(n132), .Q(product[4]) );
  XNOR2X1 U377 ( .IN1(n133), .IN2(n22), .Q(n423) );
  INVX0 U378 ( .INP(n542), .ZN(n460) );
  NBUFFX2 U379 ( .INP(a[5]), .Z(n452) );
  NBUFFX2 U380 ( .INP(a[3]), .Z(n450) );
  XOR2X1 U381 ( .IN1(b[5]), .IN2(n444), .Q(n493) );
  AND2X1 U382 ( .IN1(n499), .IN2(n554), .Q(n472) );
  AND2X1 U383 ( .IN1(n520), .IN2(n558), .Q(n481) );
  AND2X1 U384 ( .IN1(n509), .IN2(n556), .Q(n478) );
  AND2X1 U385 ( .IN1(n531), .IN2(n560), .Q(n484) );
  AND2X1 U386 ( .IN1(n542), .IN2(n562), .Q(n487) );
  NBUFFX2 U387 ( .INP(a[7]), .Z(n454) );
  NBUFFX2 U388 ( .INP(a[9]), .Z(n456) );
  NAND2X0 U389 ( .IN1(n37), .IN2(n34), .QN(n424) );
  NAND2X0 U390 ( .IN1(n37), .IN2(n8), .QN(n425) );
  NAND2X0 U391 ( .IN1(n34), .IN2(n8), .QN(n426) );
  NAND3X0 U392 ( .IN1(n426), .IN2(n425), .IN3(n424), .QN(n7) );
  NAND2X0 U393 ( .IN1(n33), .IN2(n30), .QN(n427) );
  NAND2X0 U394 ( .IN1(n33), .IN2(n7), .QN(n428) );
  NAND2X0 U395 ( .IN1(n30), .IN2(n7), .QN(n429) );
  NAND3X0 U396 ( .IN1(n429), .IN2(n428), .IN3(n427), .QN(n6) );
  NAND2X0 U397 ( .IN1(n86), .IN2(n95), .QN(n431) );
  NAND2X0 U398 ( .IN1(n86), .IN2(n15), .QN(n432) );
  NAND2X0 U399 ( .IN1(n95), .IN2(n15), .QN(n433) );
  NAND3X0 U400 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(n14) );
  NAND2X0 U401 ( .IN1(n76), .IN2(n85), .QN(n434) );
  NAND2X0 U402 ( .IN1(n76), .IN2(n14), .QN(n435) );
  NAND2X0 U403 ( .IN1(n85), .IN2(n14), .QN(n436) );
  NAND3X0 U404 ( .IN1(n436), .IN2(n435), .IN3(n434), .QN(n13) );
  XOR3X1 U405 ( .IN1(n221), .IN2(n200), .IN3(n210), .Q(n132) );
  NAND2X0 U406 ( .IN1(n221), .IN2(n210), .QN(n438) );
  NAND2X0 U407 ( .IN1(n200), .IN2(n210), .QN(n439) );
  NAND3X0 U408 ( .IN1(n437), .IN2(n438), .IN3(n439), .QN(n131) );
  NAND2X0 U409 ( .IN1(n133), .IN2(n22), .QN(n440) );
  NAND2X0 U410 ( .IN1(n133), .IN2(n132), .QN(n441) );
  NAND2X0 U411 ( .IN1(n22), .IN2(n132), .QN(n442) );
  NAND3X0 U412 ( .IN1(n440), .IN2(n441), .IN3(n442), .QN(n21) );
  DELLN1X2 U413 ( .INP(a[11]), .Z(n457) );
  INVX0 U414 ( .INP(n446), .ZN(n445) );
  INVX0 U415 ( .INP(b[0]), .ZN(n446) );
  INVX0 U416 ( .INP(n448), .ZN(n447) );
  INVX0 U417 ( .INP(a[0]), .ZN(n448) );
  DELLN1X2 U418 ( .INP(a[3]), .Z(n449) );
  DELLN1X2 U419 ( .INP(a[5]), .Z(n451) );
  DELLN1X2 U420 ( .INP(a[7]), .Z(n453) );
  DELLN1X2 U421 ( .INP(a[9]), .Z(n455) );
  NOR2X0 U422 ( .IN1(n448), .IN2(n446), .QN(product[0]) );
  XNOR2X1 U423 ( .IN1(n469), .IN2(n470), .Q(n84) );
  NAND2X0 U424 ( .IN1(n470), .IN2(n469), .QN(n83) );
  AOI22X1 U425 ( .IN1(n471), .IN2(n468), .IN3(n472), .IN4(n473), .QN(n469) );
  OA21X1 U426 ( .IN1(n474), .IN2(n447), .IN3(n475), .Q(n470) );
  AO22X1 U427 ( .IN1(n476), .IN2(n468), .IN3(n472), .IN4(n471), .Q(n73) );
  XOR2X1 U428 ( .IN1(b[10]), .IN2(n449), .Q(n471) );
  AO22X1 U429 ( .IN1(n477), .IN2(n466), .IN3(n478), .IN4(n479), .Q(n55) );
  AO22X1 U430 ( .IN1(n480), .IN2(n464), .IN3(n481), .IN4(n482), .Q(n41) );
  AO22X1 U431 ( .IN1(n483), .IN2(n462), .IN3(n484), .IN4(n485), .Q(n31) );
  AO22X1 U432 ( .IN1(n486), .IN2(n460), .IN3(n487), .IN4(n488), .Q(n25) );
  AO22X1 U433 ( .IN1(n447), .IN2(n489), .IN3(n474), .IN4(n446), .Q(n224) );
  AO22X1 U434 ( .IN1(n447), .IN2(n490), .IN3(n474), .IN4(n489), .Q(n223) );
  AO22X1 U435 ( .IN1(n447), .IN2(n491), .IN3(n474), .IN4(n490), .Q(n222) );
  AO22X1 U436 ( .IN1(n447), .IN2(n492), .IN3(n474), .IN4(n491), .Q(n221) );
  AO22X1 U437 ( .IN1(n447), .IN2(n493), .IN3(n474), .IN4(n492), .Q(n220) );
  AO22X1 U438 ( .IN1(n447), .IN2(n494), .IN3(n474), .IN4(n493), .Q(n219) );
  AO22X1 U439 ( .IN1(n447), .IN2(n495), .IN3(n474), .IN4(n494), .Q(n218) );
  AO22X1 U440 ( .IN1(n447), .IN2(n496), .IN3(n474), .IN4(n495), .Q(n217) );
  XOR2X1 U441 ( .IN1(n430), .IN2(n444), .Q(n495) );
  AO22X1 U442 ( .IN1(n447), .IN2(n497), .IN3(n474), .IN4(n496), .Q(n216) );
  XOR2X1 U443 ( .IN1(b[8]), .IN2(n444), .Q(n496) );
  AO22X1 U444 ( .IN1(n447), .IN2(n498), .IN3(n474), .IN4(n497), .Q(n215) );
  XOR2X1 U445 ( .IN1(b[9]), .IN2(n444), .Q(n497) );
  AO22X1 U446 ( .IN1(n447), .IN2(n475), .IN3(n474), .IN4(n498), .Q(n214) );
  XOR2X1 U447 ( .IN1(b[10]), .IN2(n444), .Q(n498) );
  XOR2X1 U448 ( .IN1(b[11]), .IN2(n444), .Q(n475) );
  NOR2X0 U449 ( .IN1(n499), .IN2(n446), .QN(n212) );
  AO22X1 U450 ( .IN1(n500), .IN2(n468), .IN3(n472), .IN4(n501), .Q(n211) );
  XOR2X1 U451 ( .IN1(n445), .IN2(n449), .Q(n501) );
  AO22X1 U452 ( .IN1(n502), .IN2(n468), .IN3(n472), .IN4(n500), .Q(n210) );
  AO22X1 U453 ( .IN1(n503), .IN2(n468), .IN3(n472), .IN4(n502), .Q(n209) );
  XOR2X1 U454 ( .IN1(n443), .IN2(n449), .Q(n502) );
  AO22X1 U455 ( .IN1(n504), .IN2(n468), .IN3(n472), .IN4(n503), .Q(n208) );
  AO22X1 U456 ( .IN1(n505), .IN2(n468), .IN3(n472), .IN4(n504), .Q(n207) );
  AO22X1 U457 ( .IN1(n506), .IN2(n468), .IN3(n472), .IN4(n505), .Q(n206) );
  XOR2X1 U458 ( .IN1(b[5]), .IN2(n449), .Q(n505) );
  AO22X1 U459 ( .IN1(n507), .IN2(n468), .IN3(n472), .IN4(n506), .Q(n205) );
  XOR2X1 U460 ( .IN1(b[6]), .IN2(n449), .Q(n506) );
  AO22X1 U461 ( .IN1(n508), .IN2(n468), .IN3(n472), .IN4(n507), .Q(n204) );
  XOR2X1 U462 ( .IN1(n430), .IN2(n449), .Q(n507) );
  AO22X1 U463 ( .IN1(n473), .IN2(n468), .IN3(n472), .IN4(n508), .Q(n203) );
  XOR2X1 U464 ( .IN1(b[8]), .IN2(n449), .Q(n508) );
  XOR2X1 U465 ( .IN1(b[9]), .IN2(n449), .Q(n473) );
  OAI21X1 U466 ( .IN1(n468), .IN2(n472), .IN3(n476), .QN(n201) );
  XOR2X1 U467 ( .IN1(b[11]), .IN2(n449), .Q(n476) );
  NOR2X0 U468 ( .IN1(n509), .IN2(n446), .QN(n200) );
  AO22X1 U469 ( .IN1(n510), .IN2(n466), .IN3(n478), .IN4(n511), .Q(n199) );
  AO22X1 U470 ( .IN1(n512), .IN2(n466), .IN3(n478), .IN4(n510), .Q(n198) );
  AO22X1 U471 ( .IN1(n513), .IN2(n466), .IN3(n478), .IN4(n512), .Q(n197) );
  XOR2X1 U472 ( .IN1(n443), .IN2(n451), .Q(n512) );
  AO22X1 U473 ( .IN1(n514), .IN2(n466), .IN3(n478), .IN4(n513), .Q(n196) );
  AO22X1 U474 ( .IN1(n515), .IN2(n466), .IN3(n478), .IN4(n514), .Q(n195) );
  AO22X1 U475 ( .IN1(n516), .IN2(n466), .IN3(n478), .IN4(n515), .Q(n194) );
  XOR2X1 U476 ( .IN1(b[5]), .IN2(n451), .Q(n515) );
  AO22X1 U477 ( .IN1(n517), .IN2(n466), .IN3(n478), .IN4(n516), .Q(n193) );
  XOR2X1 U478 ( .IN1(b[6]), .IN2(n451), .Q(n516) );
  AO22X1 U479 ( .IN1(n518), .IN2(n466), .IN3(n478), .IN4(n517), .Q(n192) );
  XOR2X1 U480 ( .IN1(n430), .IN2(n451), .Q(n517) );
  AO22X1 U481 ( .IN1(n519), .IN2(n466), .IN3(n478), .IN4(n518), .Q(n191) );
  XOR2X1 U482 ( .IN1(b[8]), .IN2(n451), .Q(n518) );
  AO22X1 U483 ( .IN1(n479), .IN2(n466), .IN3(n478), .IN4(n519), .Q(n190) );
  XOR2X1 U484 ( .IN1(b[9]), .IN2(n451), .Q(n519) );
  XOR2X1 U485 ( .IN1(b[10]), .IN2(n451), .Q(n479) );
  OAI21X1 U486 ( .IN1(n466), .IN2(n478), .IN3(n477), .QN(n189) );
  XOR2X1 U487 ( .IN1(b[11]), .IN2(n451), .Q(n477) );
  NOR2X0 U488 ( .IN1(n520), .IN2(n446), .QN(n188) );
  AO22X1 U489 ( .IN1(n521), .IN2(n464), .IN3(n481), .IN4(n522), .Q(n187) );
  AO22X1 U490 ( .IN1(n523), .IN2(n464), .IN3(n481), .IN4(n521), .Q(n186) );
  AO22X1 U491 ( .IN1(n524), .IN2(n464), .IN3(n481), .IN4(n523), .Q(n185) );
  XOR2X1 U492 ( .IN1(n443), .IN2(n453), .Q(n523) );
  AO22X1 U493 ( .IN1(n525), .IN2(n464), .IN3(n481), .IN4(n524), .Q(n184) );
  AO22X1 U494 ( .IN1(n526), .IN2(n464), .IN3(n481), .IN4(n525), .Q(n183) );
  AO22X1 U495 ( .IN1(n527), .IN2(n464), .IN3(n481), .IN4(n526), .Q(n182) );
  XOR2X1 U496 ( .IN1(b[5]), .IN2(n453), .Q(n526) );
  AO22X1 U497 ( .IN1(n528), .IN2(n464), .IN3(n481), .IN4(n527), .Q(n181) );
  XOR2X1 U498 ( .IN1(b[6]), .IN2(n453), .Q(n527) );
  AO22X1 U499 ( .IN1(n529), .IN2(n464), .IN3(n481), .IN4(n528), .Q(n180) );
  XOR2X1 U500 ( .IN1(n430), .IN2(n453), .Q(n528) );
  AO22X1 U501 ( .IN1(n530), .IN2(n464), .IN3(n481), .IN4(n529), .Q(n179) );
  XOR2X1 U502 ( .IN1(b[8]), .IN2(n453), .Q(n529) );
  AO22X1 U503 ( .IN1(n482), .IN2(n464), .IN3(n481), .IN4(n530), .Q(n178) );
  XOR2X1 U504 ( .IN1(b[9]), .IN2(n453), .Q(n530) );
  XOR2X1 U505 ( .IN1(b[10]), .IN2(n453), .Q(n482) );
  OAI21X1 U506 ( .IN1(n464), .IN2(n481), .IN3(n480), .QN(n177) );
  XOR2X1 U507 ( .IN1(b[11]), .IN2(n453), .Q(n480) );
  NOR2X0 U508 ( .IN1(n531), .IN2(n446), .QN(n176) );
  AO22X1 U509 ( .IN1(n532), .IN2(n462), .IN3(n484), .IN4(n533), .Q(n175) );
  AO22X1 U510 ( .IN1(n534), .IN2(n462), .IN3(n484), .IN4(n532), .Q(n174) );
  AO22X1 U511 ( .IN1(n535), .IN2(n462), .IN3(n484), .IN4(n534), .Q(n173) );
  XOR2X1 U512 ( .IN1(n443), .IN2(n455), .Q(n534) );
  AO22X1 U513 ( .IN1(n536), .IN2(n462), .IN3(n484), .IN4(n535), .Q(n172) );
  AO22X1 U514 ( .IN1(n537), .IN2(n462), .IN3(n484), .IN4(n536), .Q(n171) );
  AO22X1 U515 ( .IN1(n538), .IN2(n462), .IN3(n484), .IN4(n537), .Q(n170) );
  XOR2X1 U516 ( .IN1(b[5]), .IN2(n455), .Q(n537) );
  AO22X1 U517 ( .IN1(n539), .IN2(n462), .IN3(n484), .IN4(n538), .Q(n169) );
  XOR2X1 U518 ( .IN1(b[6]), .IN2(n455), .Q(n538) );
  AO22X1 U519 ( .IN1(n540), .IN2(n462), .IN3(n484), .IN4(n539), .Q(n168) );
  XOR2X1 U520 ( .IN1(n430), .IN2(n455), .Q(n539) );
  AO22X1 U521 ( .IN1(n541), .IN2(n462), .IN3(n484), .IN4(n540), .Q(n167) );
  XOR2X1 U522 ( .IN1(b[8]), .IN2(n455), .Q(n540) );
  AO22X1 U523 ( .IN1(n485), .IN2(n462), .IN3(n484), .IN4(n541), .Q(n166) );
  XOR2X1 U524 ( .IN1(b[9]), .IN2(n455), .Q(n541) );
  XOR2X1 U525 ( .IN1(b[10]), .IN2(n455), .Q(n485) );
  OAI21X1 U526 ( .IN1(n462), .IN2(n484), .IN3(n483), .QN(n165) );
  XOR2X1 U527 ( .IN1(b[11]), .IN2(n455), .Q(n483) );
  NOR2X0 U528 ( .IN1(n542), .IN2(n446), .QN(n164) );
  AO22X1 U529 ( .IN1(n543), .IN2(n460), .IN3(n487), .IN4(n544), .Q(n163) );
  AO22X1 U530 ( .IN1(n545), .IN2(n460), .IN3(n487), .IN4(n543), .Q(n162) );
  AO22X1 U531 ( .IN1(n546), .IN2(n460), .IN3(n487), .IN4(n545), .Q(n161) );
  XOR2X1 U532 ( .IN1(n443), .IN2(n457), .Q(n545) );
  AO22X1 U533 ( .IN1(n547), .IN2(n460), .IN3(n487), .IN4(n546), .Q(n160) );
  AO22X1 U534 ( .IN1(n548), .IN2(n460), .IN3(n487), .IN4(n547), .Q(n159) );
  AO22X1 U535 ( .IN1(n549), .IN2(n460), .IN3(n487), .IN4(n548), .Q(n158) );
  XOR2X1 U536 ( .IN1(b[5]), .IN2(n457), .Q(n548) );
  AO22X1 U537 ( .IN1(n550), .IN2(n460), .IN3(n487), .IN4(n549), .Q(n157) );
  XOR2X1 U538 ( .IN1(b[6]), .IN2(n457), .Q(n549) );
  AO22X1 U539 ( .IN1(n551), .IN2(n460), .IN3(n487), .IN4(n550), .Q(n156) );
  XOR2X1 U540 ( .IN1(n430), .IN2(n457), .Q(n550) );
  AO22X1 U541 ( .IN1(n552), .IN2(n460), .IN3(n487), .IN4(n551), .Q(n155) );
  XOR2X1 U542 ( .IN1(b[8]), .IN2(n457), .Q(n551) );
  AO22X1 U543 ( .IN1(n488), .IN2(n460), .IN3(n487), .IN4(n552), .Q(n154) );
  XOR2X1 U544 ( .IN1(b[9]), .IN2(n457), .Q(n552) );
  XOR2X1 U545 ( .IN1(b[10]), .IN2(n457), .Q(n488) );
  OAI21X1 U546 ( .IN1(n460), .IN2(n487), .IN3(n486), .QN(n153) );
  XOR2X1 U547 ( .IN1(b[11]), .IN2(n457), .Q(n486) );
  AO21X1 U548 ( .IN1(n444), .IN2(n446), .IN3(n474), .Q(n152) );
  AO22X1 U549 ( .IN1(n553), .IN2(n450), .IN3(n472), .IN4(n450), .Q(n151) );
  XOR2X1 U550 ( .IN1(n449), .IN2(a[2]), .Q(n554) );
  NOR2X0 U551 ( .IN1(n445), .IN2(n499), .QN(n553) );
  XNOR2X1 U552 ( .IN1(a[2]), .IN2(n444), .Q(n499) );
  AO22X1 U553 ( .IN1(n555), .IN2(n452), .IN3(n478), .IN4(n452), .Q(n150) );
  XOR2X1 U554 ( .IN1(n451), .IN2(a[4]), .Q(n556) );
  NOR2X0 U555 ( .IN1(n445), .IN2(n509), .QN(n555) );
  XNOR2X1 U556 ( .IN1(a[4]), .IN2(n449), .Q(n509) );
  AO22X1 U557 ( .IN1(n557), .IN2(n454), .IN3(n481), .IN4(n454), .Q(n149) );
  XOR2X1 U558 ( .IN1(n453), .IN2(a[6]), .Q(n558) );
  NOR2X0 U559 ( .IN1(n445), .IN2(n520), .QN(n557) );
  XNOR2X1 U560 ( .IN1(a[6]), .IN2(n451), .Q(n520) );
  AO22X1 U561 ( .IN1(n559), .IN2(n456), .IN3(n484), .IN4(n456), .Q(n148) );
  XOR2X1 U562 ( .IN1(n455), .IN2(a[8]), .Q(n560) );
  NOR2X0 U563 ( .IN1(n445), .IN2(n531), .QN(n559) );
  XNOR2X1 U564 ( .IN1(a[8]), .IN2(n453), .Q(n531) );
  AO22X1 U565 ( .IN1(n561), .IN2(n457), .IN3(n487), .IN4(n457), .Q(n147) );
  XOR2X1 U566 ( .IN1(n457), .IN2(a[10]), .Q(n562) );
  NOR2X0 U567 ( .IN1(n445), .IN2(n542), .QN(n561) );
  XNOR2X1 U568 ( .IN1(a[10]), .IN2(n455), .Q(n542) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_6 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_6_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_5_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553;

  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n452), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n454), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n456), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n458), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  AO22X1 U311 ( .IN1(n439), .IN2(n484), .IN3(n465), .IN4(n483), .Q(n220) );
  FADDX1 U312 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U313 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U314 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U315 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U316 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U317 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U318 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U319 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  AND3X1 U320 ( .IN1(n413), .IN2(n414), .IN3(n415), .Q(product[23]) );
  XOR3X2 U321 ( .IN1(n27), .IN2(n450), .IN3(n5), .Q(product[21]) );
  NAND2X0 U322 ( .IN1(n27), .IN2(n450), .QN(n409) );
  NAND2X0 U323 ( .IN1(n27), .IN2(n5), .QN(n410) );
  NAND2X0 U324 ( .IN1(n450), .IN2(n5), .QN(n411) );
  NAND3X0 U325 ( .IN1(n409), .IN2(n410), .IN3(n411), .QN(n4) );
  XOR2X2 U326 ( .IN1(n25), .IN2(n153), .Q(n412) );
  XOR2X1 U327 ( .IN1(n412), .IN2(n4), .Q(product[22]) );
  NAND2X0 U328 ( .IN1(n25), .IN2(n153), .QN(n413) );
  NAND2X0 U329 ( .IN1(n25), .IN2(n4), .QN(n414) );
  NAND2X0 U330 ( .IN1(n153), .IN2(n4), .QN(n415) );
  DELLN2X2 U331 ( .INP(n13), .Z(n416) );
  HADDX2 U332 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  XOR2X2 U333 ( .IN1(b[4]), .IN2(n449), .Q(n538) );
  XOR2X2 U334 ( .IN1(b[4]), .IN2(n447), .Q(n527) );
  XOR2X2 U335 ( .IN1(b[4]), .IN2(n445), .Q(n516) );
  XOR2X2 U336 ( .IN1(b[4]), .IN2(n443), .Q(n505) );
  XOR2X2 U337 ( .IN1(b[4]), .IN2(n441), .Q(n495) );
  XOR2X2 U338 ( .IN1(b[4]), .IN2(a[1]), .Q(n483) );
  XOR2X2 U339 ( .IN1(b[3]), .IN2(n449), .Q(n537) );
  XOR2X2 U340 ( .IN1(b[3]), .IN2(n447), .Q(n526) );
  XOR2X2 U341 ( .IN1(b[3]), .IN2(n445), .Q(n515) );
  XOR2X2 U342 ( .IN1(b[3]), .IN2(n443), .Q(n504) );
  XOR2X2 U343 ( .IN1(b[3]), .IN2(n441), .Q(n494) );
  XOR2X2 U344 ( .IN1(b[3]), .IN2(a[1]), .Q(n482) );
  XOR3X2 U345 ( .IN1(n57), .IN2(n50), .IN3(n11), .Q(product[15]) );
  NAND2X0 U346 ( .IN1(n57), .IN2(n50), .QN(n417) );
  NAND2X0 U347 ( .IN1(n57), .IN2(n11), .QN(n418) );
  NAND2X0 U348 ( .IN1(n50), .IN2(n11), .QN(n419) );
  NAND3X0 U349 ( .IN1(n417), .IN2(n418), .IN3(n419), .QN(n10) );
  XOR2X1 U350 ( .IN1(n49), .IN2(n44), .Q(n420) );
  XOR2X1 U351 ( .IN1(n420), .IN2(n10), .Q(product[16]) );
  NAND2X0 U352 ( .IN1(n49), .IN2(n44), .QN(n421) );
  NAND2X0 U353 ( .IN1(n49), .IN2(n10), .QN(n422) );
  NAND2X0 U354 ( .IN1(n44), .IN2(n10), .QN(n423) );
  NAND3X0 U355 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n9) );
  FADDX1 U356 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  XOR3X1 U357 ( .IN1(n76), .IN2(n85), .IN3(n14), .Q(product[12]) );
  XNOR2X1 U358 ( .IN1(n424), .IN2(n416), .Q(product[13]) );
  XNOR2X1 U359 ( .IN1(n66), .IN2(n75), .Q(n424) );
  XNOR2X1 U360 ( .IN1(n425), .IN2(n15), .Q(product[11]) );
  XNOR2X1 U361 ( .IN1(n95), .IN2(n86), .Q(n425) );
  INVX0 U362 ( .INP(n25), .ZN(n450) );
  FADDX1 U363 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U364 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  INVX0 U365 ( .INP(n55), .ZN(n456) );
  XOR2X1 U366 ( .IN1(b[1]), .IN2(a[1]), .Q(n480) );
  XOR2X1 U367 ( .IN1(b[1]), .IN2(n441), .Q(n491) );
  XOR2X1 U368 ( .IN1(b[1]), .IN2(n443), .Q(n501) );
  XOR2X1 U369 ( .IN1(b[1]), .IN2(n445), .Q(n512) );
  INVX0 U370 ( .INP(n73), .ZN(n458) );
  XOR2X1 U371 ( .IN1(b[1]), .IN2(n447), .Q(n523) );
  XOR2X1 U372 ( .IN1(b[1]), .IN2(n449), .Q(n534) );
  INVX0 U373 ( .INP(n31), .ZN(n452) );
  INVX0 U374 ( .INP(n41), .ZN(n454) );
  XOR2X1 U375 ( .IN1(b[2]), .IN2(a[1]), .Q(n481) );
  INVX0 U376 ( .INP(n490), .ZN(n459) );
  INVX0 U377 ( .INP(n500), .ZN(n457) );
  INVX0 U378 ( .INP(n511), .ZN(n455) );
  INVX0 U379 ( .INP(n522), .ZN(n453) );
  AND2X1 U380 ( .IN1(a[1]), .IN2(n440), .Q(n465) );
  INVX0 U381 ( .INP(n533), .ZN(n451) );
  NBUFFX2 U382 ( .INP(a[3]), .Z(n442) );
  NBUFFX2 U383 ( .INP(a[5]), .Z(n444) );
  NBUFFX2 U384 ( .INP(b[5]), .Z(n435) );
  AND2X1 U385 ( .IN1(n490), .IN2(n545), .Q(n463) );
  AND2X1 U386 ( .IN1(n511), .IN2(n549), .Q(n472) );
  AND2X1 U387 ( .IN1(n500), .IN2(n547), .Q(n469) );
  AND2X1 U388 ( .IN1(n522), .IN2(n551), .Q(n475) );
  AND2X1 U389 ( .IN1(n533), .IN2(n553), .Q(n478) );
  NBUFFX2 U390 ( .INP(a[7]), .Z(n446) );
  NBUFFX2 U391 ( .INP(a[9]), .Z(n448) );
  NAND2X0 U392 ( .IN1(n76), .IN2(n85), .QN(n426) );
  NAND2X0 U393 ( .IN1(n76), .IN2(n14), .QN(n427) );
  NAND2X0 U394 ( .IN1(n85), .IN2(n14), .QN(n428) );
  NAND3X0 U395 ( .IN1(n428), .IN2(n427), .IN3(n426), .QN(n13) );
  NAND2X0 U396 ( .IN1(n66), .IN2(n75), .QN(n429) );
  NAND2X0 U397 ( .IN1(n66), .IN2(n13), .QN(n430) );
  NAND2X0 U398 ( .IN1(n75), .IN2(n13), .QN(n431) );
  NAND3X0 U399 ( .IN1(n431), .IN2(n430), .IN3(n429), .QN(n12) );
  NAND2X0 U400 ( .IN1(n86), .IN2(n15), .QN(n432) );
  NAND2X0 U401 ( .IN1(n95), .IN2(n15), .QN(n433) );
  NAND2X0 U402 ( .IN1(n95), .IN2(n86), .QN(n434) );
  NAND3X0 U403 ( .IN1(n432), .IN2(n434), .IN3(n433), .QN(n14) );
  DELLN1X2 U404 ( .INP(a[11]), .Z(n449) );
  INVX0 U405 ( .INP(n438), .ZN(n436) );
  INVX0 U406 ( .INP(b[0]), .ZN(n437) );
  INVX0 U407 ( .INP(b[0]), .ZN(n438) );
  INVX0 U408 ( .INP(n440), .ZN(n439) );
  INVX0 U409 ( .INP(a[0]), .ZN(n440) );
  DELLN1X2 U410 ( .INP(a[3]), .Z(n441) );
  DELLN1X2 U411 ( .INP(a[5]), .Z(n443) );
  DELLN1X2 U412 ( .INP(a[7]), .Z(n445) );
  DELLN1X2 U413 ( .INP(a[9]), .Z(n447) );
  NOR2X0 U414 ( .IN1(n440), .IN2(n438), .QN(product[0]) );
  XNOR2X1 U415 ( .IN1(n460), .IN2(n461), .Q(n84) );
  NAND2X0 U416 ( .IN1(n461), .IN2(n460), .QN(n83) );
  AOI22X1 U417 ( .IN1(n462), .IN2(n459), .IN3(n463), .IN4(n464), .QN(n460) );
  OA21X1 U418 ( .IN1(n465), .IN2(n439), .IN3(n466), .Q(n461) );
  AO22X1 U419 ( .IN1(n467), .IN2(n459), .IN3(n463), .IN4(n462), .Q(n73) );
  XOR2X1 U420 ( .IN1(b[10]), .IN2(n441), .Q(n462) );
  AO22X1 U421 ( .IN1(n468), .IN2(n457), .IN3(n469), .IN4(n470), .Q(n55) );
  AO22X1 U422 ( .IN1(n471), .IN2(n455), .IN3(n472), .IN4(n473), .Q(n41) );
  AO22X1 U423 ( .IN1(n474), .IN2(n453), .IN3(n475), .IN4(n476), .Q(n31) );
  AO22X1 U424 ( .IN1(n477), .IN2(n451), .IN3(n478), .IN4(n479), .Q(n25) );
  AO22X1 U425 ( .IN1(n439), .IN2(n480), .IN3(n465), .IN4(n437), .Q(n224) );
  AO22X1 U426 ( .IN1(n439), .IN2(n481), .IN3(n465), .IN4(n480), .Q(n223) );
  AO22X1 U427 ( .IN1(n439), .IN2(n482), .IN3(n465), .IN4(n481), .Q(n222) );
  AO22X1 U428 ( .IN1(n439), .IN2(n483), .IN3(n465), .IN4(n482), .Q(n221) );
  AO22X1 U429 ( .IN1(n439), .IN2(n485), .IN3(n465), .IN4(n484), .Q(n219) );
  XOR2X1 U430 ( .IN1(n435), .IN2(a[1]), .Q(n484) );
  AO22X1 U431 ( .IN1(n439), .IN2(n486), .IN3(n465), .IN4(n485), .Q(n218) );
  XOR2X1 U432 ( .IN1(b[6]), .IN2(a[1]), .Q(n485) );
  AO22X1 U433 ( .IN1(n439), .IN2(n487), .IN3(n465), .IN4(n486), .Q(n217) );
  XOR2X1 U434 ( .IN1(b[7]), .IN2(a[1]), .Q(n486) );
  AO22X1 U435 ( .IN1(n439), .IN2(n488), .IN3(n465), .IN4(n487), .Q(n216) );
  XOR2X1 U436 ( .IN1(b[8]), .IN2(a[1]), .Q(n487) );
  AO22X1 U437 ( .IN1(n439), .IN2(n489), .IN3(n465), .IN4(n488), .Q(n215) );
  XOR2X1 U438 ( .IN1(b[9]), .IN2(a[1]), .Q(n488) );
  AO22X1 U439 ( .IN1(n439), .IN2(n466), .IN3(n465), .IN4(n489), .Q(n214) );
  XOR2X1 U440 ( .IN1(b[10]), .IN2(a[1]), .Q(n489) );
  XOR2X1 U441 ( .IN1(b[11]), .IN2(a[1]), .Q(n466) );
  NOR2X0 U442 ( .IN1(n490), .IN2(n438), .QN(n212) );
  AO22X1 U443 ( .IN1(n491), .IN2(n459), .IN3(n463), .IN4(n492), .Q(n211) );
  XOR2X1 U444 ( .IN1(n436), .IN2(n441), .Q(n492) );
  AO22X1 U445 ( .IN1(n493), .IN2(n459), .IN3(n463), .IN4(n491), .Q(n210) );
  AO22X1 U446 ( .IN1(n494), .IN2(n459), .IN3(n463), .IN4(n493), .Q(n209) );
  XOR2X1 U447 ( .IN1(b[2]), .IN2(n441), .Q(n493) );
  AO22X1 U448 ( .IN1(n495), .IN2(n459), .IN3(n463), .IN4(n494), .Q(n208) );
  AO22X1 U449 ( .IN1(n496), .IN2(n459), .IN3(n463), .IN4(n495), .Q(n207) );
  AO22X1 U450 ( .IN1(n497), .IN2(n459), .IN3(n463), .IN4(n496), .Q(n206) );
  XOR2X1 U451 ( .IN1(n435), .IN2(n441), .Q(n496) );
  AO22X1 U452 ( .IN1(n498), .IN2(n459), .IN3(n463), .IN4(n497), .Q(n205) );
  XOR2X1 U453 ( .IN1(b[6]), .IN2(n441), .Q(n497) );
  AO22X1 U454 ( .IN1(n499), .IN2(n459), .IN3(n463), .IN4(n498), .Q(n204) );
  XOR2X1 U455 ( .IN1(b[7]), .IN2(n441), .Q(n498) );
  AO22X1 U456 ( .IN1(n464), .IN2(n459), .IN3(n463), .IN4(n499), .Q(n203) );
  XOR2X1 U457 ( .IN1(b[8]), .IN2(n441), .Q(n499) );
  XOR2X1 U458 ( .IN1(b[9]), .IN2(n441), .Q(n464) );
  OAI21X1 U459 ( .IN1(n459), .IN2(n463), .IN3(n467), .QN(n201) );
  XOR2X1 U460 ( .IN1(b[11]), .IN2(n441), .Q(n467) );
  NOR2X0 U461 ( .IN1(n500), .IN2(n438), .QN(n200) );
  AO22X1 U462 ( .IN1(n501), .IN2(n457), .IN3(n469), .IN4(n502), .Q(n199) );
  XOR2X1 U463 ( .IN1(n436), .IN2(n443), .Q(n502) );
  AO22X1 U464 ( .IN1(n503), .IN2(n457), .IN3(n469), .IN4(n501), .Q(n198) );
  AO22X1 U465 ( .IN1(n504), .IN2(n457), .IN3(n469), .IN4(n503), .Q(n197) );
  XOR2X1 U466 ( .IN1(b[2]), .IN2(n443), .Q(n503) );
  AO22X1 U467 ( .IN1(n505), .IN2(n457), .IN3(n469), .IN4(n504), .Q(n196) );
  AO22X1 U468 ( .IN1(n506), .IN2(n457), .IN3(n469), .IN4(n505), .Q(n195) );
  AO22X1 U469 ( .IN1(n507), .IN2(n457), .IN3(n469), .IN4(n506), .Q(n194) );
  XOR2X1 U470 ( .IN1(n435), .IN2(n443), .Q(n506) );
  AO22X1 U471 ( .IN1(n508), .IN2(n457), .IN3(n469), .IN4(n507), .Q(n193) );
  XOR2X1 U472 ( .IN1(b[6]), .IN2(n443), .Q(n507) );
  AO22X1 U473 ( .IN1(n509), .IN2(n457), .IN3(n469), .IN4(n508), .Q(n192) );
  XOR2X1 U474 ( .IN1(b[7]), .IN2(n443), .Q(n508) );
  AO22X1 U475 ( .IN1(n510), .IN2(n457), .IN3(n469), .IN4(n509), .Q(n191) );
  XOR2X1 U476 ( .IN1(b[8]), .IN2(n443), .Q(n509) );
  AO22X1 U477 ( .IN1(n470), .IN2(n457), .IN3(n469), .IN4(n510), .Q(n190) );
  XOR2X1 U478 ( .IN1(b[9]), .IN2(n443), .Q(n510) );
  XOR2X1 U479 ( .IN1(b[10]), .IN2(n443), .Q(n470) );
  OAI21X1 U480 ( .IN1(n457), .IN2(n469), .IN3(n468), .QN(n189) );
  XOR2X1 U481 ( .IN1(b[11]), .IN2(n443), .Q(n468) );
  NOR2X0 U482 ( .IN1(n511), .IN2(n437), .QN(n188) );
  AO22X1 U483 ( .IN1(n512), .IN2(n455), .IN3(n472), .IN4(n513), .Q(n187) );
  XOR2X1 U484 ( .IN1(n436), .IN2(n445), .Q(n513) );
  AO22X1 U485 ( .IN1(n514), .IN2(n455), .IN3(n472), .IN4(n512), .Q(n186) );
  AO22X1 U486 ( .IN1(n515), .IN2(n455), .IN3(n472), .IN4(n514), .Q(n185) );
  XOR2X1 U487 ( .IN1(b[2]), .IN2(n445), .Q(n514) );
  AO22X1 U488 ( .IN1(n516), .IN2(n455), .IN3(n472), .IN4(n515), .Q(n184) );
  AO22X1 U489 ( .IN1(n517), .IN2(n455), .IN3(n472), .IN4(n516), .Q(n183) );
  AO22X1 U490 ( .IN1(n518), .IN2(n455), .IN3(n472), .IN4(n517), .Q(n182) );
  XOR2X1 U491 ( .IN1(n435), .IN2(n445), .Q(n517) );
  AO22X1 U492 ( .IN1(n519), .IN2(n455), .IN3(n472), .IN4(n518), .Q(n181) );
  XOR2X1 U493 ( .IN1(b[6]), .IN2(n445), .Q(n518) );
  AO22X1 U494 ( .IN1(n520), .IN2(n455), .IN3(n472), .IN4(n519), .Q(n180) );
  XOR2X1 U495 ( .IN1(b[7]), .IN2(n445), .Q(n519) );
  AO22X1 U496 ( .IN1(n521), .IN2(n455), .IN3(n472), .IN4(n520), .Q(n179) );
  XOR2X1 U497 ( .IN1(b[8]), .IN2(n445), .Q(n520) );
  AO22X1 U498 ( .IN1(n473), .IN2(n455), .IN3(n472), .IN4(n521), .Q(n178) );
  XOR2X1 U499 ( .IN1(b[9]), .IN2(n445), .Q(n521) );
  XOR2X1 U500 ( .IN1(b[10]), .IN2(n445), .Q(n473) );
  OAI21X1 U501 ( .IN1(n455), .IN2(n472), .IN3(n471), .QN(n177) );
  XOR2X1 U502 ( .IN1(b[11]), .IN2(n445), .Q(n471) );
  NOR2X0 U503 ( .IN1(n522), .IN2(n437), .QN(n176) );
  AO22X1 U504 ( .IN1(n523), .IN2(n453), .IN3(n475), .IN4(n524), .Q(n175) );
  XOR2X1 U505 ( .IN1(n436), .IN2(n447), .Q(n524) );
  AO22X1 U506 ( .IN1(n525), .IN2(n453), .IN3(n475), .IN4(n523), .Q(n174) );
  AO22X1 U507 ( .IN1(n526), .IN2(n453), .IN3(n475), .IN4(n525), .Q(n173) );
  XOR2X1 U508 ( .IN1(b[2]), .IN2(n447), .Q(n525) );
  AO22X1 U509 ( .IN1(n527), .IN2(n453), .IN3(n475), .IN4(n526), .Q(n172) );
  AO22X1 U510 ( .IN1(n528), .IN2(n453), .IN3(n475), .IN4(n527), .Q(n171) );
  AO22X1 U511 ( .IN1(n529), .IN2(n453), .IN3(n475), .IN4(n528), .Q(n170) );
  XOR2X1 U512 ( .IN1(n435), .IN2(n447), .Q(n528) );
  AO22X1 U513 ( .IN1(n530), .IN2(n453), .IN3(n475), .IN4(n529), .Q(n169) );
  XOR2X1 U514 ( .IN1(b[6]), .IN2(n447), .Q(n529) );
  AO22X1 U515 ( .IN1(n531), .IN2(n453), .IN3(n475), .IN4(n530), .Q(n168) );
  XOR2X1 U516 ( .IN1(b[7]), .IN2(n447), .Q(n530) );
  AO22X1 U517 ( .IN1(n532), .IN2(n453), .IN3(n475), .IN4(n531), .Q(n167) );
  XOR2X1 U518 ( .IN1(b[8]), .IN2(n447), .Q(n531) );
  AO22X1 U519 ( .IN1(n476), .IN2(n453), .IN3(n475), .IN4(n532), .Q(n166) );
  XOR2X1 U520 ( .IN1(b[9]), .IN2(n447), .Q(n532) );
  XOR2X1 U521 ( .IN1(b[10]), .IN2(n447), .Q(n476) );
  OAI21X1 U522 ( .IN1(n453), .IN2(n475), .IN3(n474), .QN(n165) );
  XOR2X1 U523 ( .IN1(b[11]), .IN2(n447), .Q(n474) );
  NOR2X0 U524 ( .IN1(n533), .IN2(n437), .QN(n164) );
  AO22X1 U525 ( .IN1(n534), .IN2(n451), .IN3(n478), .IN4(n535), .Q(n163) );
  XOR2X1 U526 ( .IN1(n436), .IN2(n449), .Q(n535) );
  AO22X1 U527 ( .IN1(n536), .IN2(n451), .IN3(n478), .IN4(n534), .Q(n162) );
  AO22X1 U528 ( .IN1(n537), .IN2(n451), .IN3(n478), .IN4(n536), .Q(n161) );
  XOR2X1 U529 ( .IN1(b[2]), .IN2(n449), .Q(n536) );
  AO22X1 U530 ( .IN1(n538), .IN2(n451), .IN3(n478), .IN4(n537), .Q(n160) );
  AO22X1 U531 ( .IN1(n539), .IN2(n451), .IN3(n478), .IN4(n538), .Q(n159) );
  AO22X1 U532 ( .IN1(n540), .IN2(n451), .IN3(n478), .IN4(n539), .Q(n158) );
  XOR2X1 U533 ( .IN1(n435), .IN2(n449), .Q(n539) );
  AO22X1 U534 ( .IN1(n541), .IN2(n451), .IN3(n478), .IN4(n540), .Q(n157) );
  XOR2X1 U535 ( .IN1(b[6]), .IN2(n449), .Q(n540) );
  AO22X1 U536 ( .IN1(n542), .IN2(n451), .IN3(n478), .IN4(n541), .Q(n156) );
  XOR2X1 U537 ( .IN1(b[7]), .IN2(n449), .Q(n541) );
  AO22X1 U538 ( .IN1(n543), .IN2(n451), .IN3(n478), .IN4(n542), .Q(n155) );
  XOR2X1 U539 ( .IN1(b[8]), .IN2(n449), .Q(n542) );
  AO22X1 U540 ( .IN1(n479), .IN2(n451), .IN3(n478), .IN4(n543), .Q(n154) );
  XOR2X1 U541 ( .IN1(b[9]), .IN2(n449), .Q(n543) );
  XOR2X1 U542 ( .IN1(b[10]), .IN2(n449), .Q(n479) );
  OAI21X1 U543 ( .IN1(n451), .IN2(n478), .IN3(n477), .QN(n153) );
  XOR2X1 U544 ( .IN1(b[11]), .IN2(n449), .Q(n477) );
  AO21X1 U545 ( .IN1(a[1]), .IN2(n437), .IN3(n465), .Q(n152) );
  AO22X1 U546 ( .IN1(n544), .IN2(n442), .IN3(n463), .IN4(n442), .Q(n151) );
  XOR2X1 U547 ( .IN1(n441), .IN2(a[2]), .Q(n545) );
  NOR2X0 U548 ( .IN1(n436), .IN2(n490), .QN(n544) );
  XNOR2X1 U549 ( .IN1(a[2]), .IN2(a[1]), .Q(n490) );
  AO22X1 U550 ( .IN1(n546), .IN2(n444), .IN3(n469), .IN4(n444), .Q(n150) );
  XOR2X1 U551 ( .IN1(n443), .IN2(a[4]), .Q(n547) );
  NOR2X0 U552 ( .IN1(n436), .IN2(n500), .QN(n546) );
  XNOR2X1 U553 ( .IN1(a[4]), .IN2(n441), .Q(n500) );
  AO22X1 U554 ( .IN1(n548), .IN2(n446), .IN3(n472), .IN4(n446), .Q(n149) );
  XOR2X1 U555 ( .IN1(n445), .IN2(a[6]), .Q(n549) );
  NOR2X0 U556 ( .IN1(n436), .IN2(n511), .QN(n548) );
  XNOR2X1 U557 ( .IN1(a[6]), .IN2(n443), .Q(n511) );
  AO22X1 U558 ( .IN1(n550), .IN2(n448), .IN3(n475), .IN4(n448), .Q(n148) );
  XOR2X1 U559 ( .IN1(n447), .IN2(a[8]), .Q(n551) );
  NOR2X0 U560 ( .IN1(n436), .IN2(n522), .QN(n550) );
  XNOR2X1 U561 ( .IN1(a[8]), .IN2(n445), .Q(n522) );
  AO22X1 U562 ( .IN1(n552), .IN2(n449), .IN3(n478), .IN4(n449), .Q(n147) );
  XOR2X1 U563 ( .IN1(n449), .IN2(a[10]), .Q(n553) );
  NOR2X0 U564 ( .IN1(n436), .IN2(n533), .QN(n552) );
  XNOR2X1 U565 ( .IN1(a[10]), .IN2(n447), .Q(n533) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_5 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;
  wire   n1;
  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_5_DW_mult_tc_0 mult_30 ( .a(in_a), .b({
        in_b[11:2], n1, in_b[0]}), .product(pre_out) );
  DELLN1X2 U3 ( .INP(in_b[1]), .Z(n1) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_4_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n456), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n458), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n460), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n462), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  XOR3X1 U311 ( .IN1(n223), .IN2(n212), .IN3(n24), .Q(product[2]) );
  FADDX1 U312 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U313 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U314 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U315 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U316 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U317 ( .A(n27), .B(n454), .CI(n5), .CO(n4), .S(product[21]) );
  INVX0 U318 ( .INP(b[4]), .ZN(n408) );
  INVX0 U319 ( .INP(n408), .ZN(n409) );
  XOR2X2 U320 ( .IN1(b[2]), .IN2(n452), .Q(n540) );
  XOR2X2 U321 ( .IN1(b[2]), .IN2(n450), .Q(n529) );
  XOR2X2 U322 ( .IN1(b[2]), .IN2(n448), .Q(n518) );
  XOR2X2 U323 ( .IN1(b[2]), .IN2(n446), .Q(n507) );
  XOR2X2 U324 ( .IN1(b[2]), .IN2(n444), .Q(n497) );
  XOR2X2 U325 ( .IN1(b[2]), .IN2(a[1]), .Q(n485) );
  XOR2X2 U326 ( .IN1(b[8]), .IN2(n452), .Q(n546) );
  XOR2X2 U327 ( .IN1(b[8]), .IN2(n450), .Q(n535) );
  XOR2X2 U328 ( .IN1(b[8]), .IN2(n448), .Q(n524) );
  XOR2X2 U329 ( .IN1(b[8]), .IN2(n446), .Q(n513) );
  XOR2X2 U330 ( .IN1(b[8]), .IN2(n444), .Q(n503) );
  XOR2X2 U331 ( .IN1(b[8]), .IN2(a[1]), .Q(n491) );
  XOR2X2 U332 ( .IN1(b[6]), .IN2(n452), .Q(n544) );
  XOR2X2 U333 ( .IN1(b[6]), .IN2(n450), .Q(n533) );
  XOR2X2 U334 ( .IN1(b[6]), .IN2(n448), .Q(n522) );
  XOR2X2 U335 ( .IN1(b[6]), .IN2(n446), .Q(n511) );
  XOR2X2 U336 ( .IN1(b[6]), .IN2(n444), .Q(n501) );
  XOR3X2 U337 ( .IN1(n37), .IN2(n34), .IN3(n8), .Q(product[18]) );
  NAND2X0 U338 ( .IN1(n37), .IN2(n34), .QN(n410) );
  NAND2X0 U339 ( .IN1(n37), .IN2(n8), .QN(n411) );
  NAND2X0 U340 ( .IN1(n34), .IN2(n8), .QN(n412) );
  NAND3X0 U341 ( .IN1(n410), .IN2(n411), .IN3(n412), .QN(n7) );
  XOR2X1 U342 ( .IN1(n33), .IN2(n30), .Q(n413) );
  XOR2X1 U343 ( .IN1(n413), .IN2(n7), .Q(product[19]) );
  NAND2X0 U344 ( .IN1(n33), .IN2(n30), .QN(n414) );
  NAND2X0 U345 ( .IN1(n33), .IN2(n7), .QN(n415) );
  NAND2X0 U346 ( .IN1(n30), .IN2(n7), .QN(n416) );
  NAND3X0 U347 ( .IN1(n414), .IN2(n415), .IN3(n416), .QN(n6) );
  XOR3X2 U348 ( .IN1(n86), .IN2(n95), .IN3(n15), .Q(product[11]) );
  NAND2X0 U349 ( .IN1(n86), .IN2(n95), .QN(n417) );
  NAND2X0 U350 ( .IN1(n86), .IN2(n15), .QN(n418) );
  NAND2X0 U351 ( .IN1(n95), .IN2(n15), .QN(n419) );
  NAND3X0 U352 ( .IN1(n417), .IN2(n418), .IN3(n419), .QN(n14) );
  XOR2X1 U353 ( .IN1(n76), .IN2(n85), .Q(n420) );
  XOR2X1 U354 ( .IN1(n420), .IN2(n14), .Q(product[12]) );
  NAND2X0 U355 ( .IN1(n76), .IN2(n85), .QN(n421) );
  NAND2X0 U356 ( .IN1(n76), .IN2(n14), .QN(n422) );
  NAND2X0 U357 ( .IN1(n85), .IN2(n14), .QN(n423) );
  NAND3X0 U358 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n13) );
  NAND2X0 U359 ( .IN1(n223), .IN2(n212), .QN(n424) );
  NAND2X0 U360 ( .IN1(n223), .IN2(n24), .QN(n425) );
  NAND2X0 U361 ( .IN1(n212), .IN2(n24), .QN(n426) );
  NAND3X0 U362 ( .IN1(n424), .IN2(n425), .IN3(n426), .QN(n23) );
  XOR2X2 U363 ( .IN1(n134), .IN2(n151), .Q(n427) );
  XOR2X1 U364 ( .IN1(n427), .IN2(n23), .Q(product[3]) );
  NAND2X0 U365 ( .IN1(n134), .IN2(n151), .QN(n428) );
  NAND2X0 U366 ( .IN1(n134), .IN2(n23), .QN(n429) );
  NAND2X0 U367 ( .IN1(n151), .IN2(n23), .QN(n430) );
  NAND3X0 U368 ( .IN1(n428), .IN2(n429), .IN3(n430), .QN(n22) );
  XOR2X2 U369 ( .IN1(n409), .IN2(n452), .Q(n542) );
  XOR2X2 U370 ( .IN1(n409), .IN2(n450), .Q(n531) );
  XOR2X2 U371 ( .IN1(n409), .IN2(n448), .Q(n520) );
  XOR2X2 U372 ( .IN1(n409), .IN2(n446), .Q(n509) );
  XOR2X2 U373 ( .IN1(n409), .IN2(n444), .Q(n499) );
  DELLN2X2 U374 ( .INP(n12), .Z(n431) );
  FADDX1 U375 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  XOR2X2 U376 ( .IN1(b[3]), .IN2(n452), .Q(n541) );
  XOR2X2 U377 ( .IN1(b[3]), .IN2(n450), .Q(n530) );
  XOR2X2 U378 ( .IN1(b[3]), .IN2(n448), .Q(n519) );
  XOR2X2 U379 ( .IN1(b[3]), .IN2(n446), .Q(n508) );
  XOR2X2 U380 ( .IN1(b[3]), .IN2(n444), .Q(n498) );
  XOR2X2 U381 ( .IN1(b[3]), .IN2(a[1]), .Q(n486) );
  XOR2X2 U382 ( .IN1(b[5]), .IN2(n452), .Q(n543) );
  XOR2X2 U383 ( .IN1(b[5]), .IN2(n450), .Q(n532) );
  XOR2X2 U384 ( .IN1(b[5]), .IN2(n448), .Q(n521) );
  XOR2X2 U385 ( .IN1(b[5]), .IN2(n446), .Q(n510) );
  XOR2X2 U386 ( .IN1(b[5]), .IN2(n444), .Q(n500) );
  XOR2X2 U387 ( .IN1(b[1]), .IN2(n452), .Q(n538) );
  XOR2X2 U388 ( .IN1(b[1]), .IN2(n450), .Q(n527) );
  XOR2X2 U389 ( .IN1(b[1]), .IN2(n448), .Q(n516) );
  XOR2X2 U390 ( .IN1(b[1]), .IN2(n446), .Q(n505) );
  XOR2X2 U391 ( .IN1(b[1]), .IN2(n444), .Q(n495) );
  XOR2X2 U392 ( .IN1(b[1]), .IN2(a[1]), .Q(n484) );
  XOR3X1 U393 ( .IN1(n66), .IN2(n75), .IN3(n13), .Q(product[13]) );
  NAND2X0 U394 ( .IN1(n66), .IN2(n75), .QN(n432) );
  NAND2X0 U395 ( .IN1(n65), .IN2(n58), .QN(n436) );
  NAND2X0 U396 ( .IN1(n66), .IN2(n13), .QN(n433) );
  NAND2X0 U397 ( .IN1(n75), .IN2(n13), .QN(n434) );
  NAND3X0 U398 ( .IN1(n432), .IN2(n433), .IN3(n434), .QN(n12) );
  XOR2X1 U399 ( .IN1(n65), .IN2(n58), .Q(n435) );
  XOR2X1 U400 ( .IN1(n435), .IN2(n431), .Q(product[14]) );
  NAND2X0 U401 ( .IN1(n65), .IN2(n12), .QN(n437) );
  NAND2X0 U402 ( .IN1(n58), .IN2(n12), .QN(n438) );
  NAND3X0 U403 ( .IN1(n438), .IN2(n437), .IN3(n436), .QN(n11) );
  INVX0 U404 ( .INP(n25), .ZN(n454) );
  INVX0 U405 ( .INP(n3), .ZN(product[23]) );
  INVX0 U406 ( .INP(n55), .ZN(n460) );
  INVX0 U407 ( .INP(n73), .ZN(n462) );
  FADDX1 U408 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U409 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  INVX0 U410 ( .INP(n31), .ZN(n456) );
  INVX0 U411 ( .INP(n41), .ZN(n458) );
  INVX0 U412 ( .INP(n504), .ZN(n461) );
  INVX0 U413 ( .INP(n494), .ZN(n463) );
  AND2X1 U414 ( .IN1(a[1]), .IN2(n443), .Q(n469) );
  INVX0 U415 ( .INP(n526), .ZN(n457) );
  INVX0 U416 ( .INP(n515), .ZN(n459) );
  INVX0 U417 ( .INP(n537), .ZN(n455) );
  NBUFFX2 U418 ( .INP(a[5]), .Z(n447) );
  NBUFFX2 U419 ( .INP(a[3]), .Z(n445) );
  NBUFFX2 U420 ( .INP(a[9]), .Z(n451) );
  XOR2X2 U421 ( .IN1(b[6]), .IN2(a[1]), .Q(n489) );
  XOR2X2 U422 ( .IN1(b[5]), .IN2(a[1]), .Q(n488) );
  XOR2X2 U423 ( .IN1(n409), .IN2(a[1]), .Q(n487) );
  DELLN1X2 U424 ( .INP(a[11]), .Z(n452) );
  AND2X2 U425 ( .IN1(n494), .IN2(n549), .Q(n467) );
  AND2X2 U426 ( .IN1(n504), .IN2(n551), .Q(n473) );
  AND2X2 U427 ( .IN1(n515), .IN2(n553), .Q(n476) );
  AND2X2 U428 ( .IN1(n526), .IN2(n555), .Q(n479) );
  AND2X2 U429 ( .IN1(n537), .IN2(n557), .Q(n482) );
  INVX0 U430 ( .INP(n441), .ZN(n439) );
  INVX0 U431 ( .INP(b[0]), .ZN(n440) );
  INVX0 U432 ( .INP(b[0]), .ZN(n441) );
  INVX0 U433 ( .INP(n443), .ZN(n442) );
  INVX0 U434 ( .INP(a[0]), .ZN(n443) );
  DELLN1X2 U435 ( .INP(a[3]), .Z(n444) );
  DELLN1X2 U436 ( .INP(a[5]), .Z(n446) );
  DELLN1X2 U437 ( .INP(a[7]), .Z(n448) );
  DELLN1X2 U438 ( .INP(a[7]), .Z(n449) );
  DELLN1X2 U439 ( .INP(a[9]), .Z(n450) );
  NOR2X0 U440 ( .IN1(n443), .IN2(n440), .QN(product[0]) );
  XNOR2X1 U441 ( .IN1(n464), .IN2(n465), .Q(n84) );
  NAND2X0 U442 ( .IN1(n465), .IN2(n464), .QN(n83) );
  AOI22X1 U443 ( .IN1(n466), .IN2(n463), .IN3(n467), .IN4(n468), .QN(n464) );
  OA21X1 U444 ( .IN1(n469), .IN2(n442), .IN3(n470), .Q(n465) );
  AO22X1 U445 ( .IN1(n471), .IN2(n463), .IN3(n467), .IN4(n466), .Q(n73) );
  XOR2X1 U446 ( .IN1(b[10]), .IN2(n444), .Q(n466) );
  AO22X1 U447 ( .IN1(n472), .IN2(n461), .IN3(n473), .IN4(n474), .Q(n55) );
  AO22X1 U448 ( .IN1(n475), .IN2(n459), .IN3(n476), .IN4(n477), .Q(n41) );
  AO22X1 U449 ( .IN1(n478), .IN2(n457), .IN3(n479), .IN4(n480), .Q(n31) );
  AO22X1 U450 ( .IN1(n481), .IN2(n455), .IN3(n482), .IN4(n483), .Q(n25) );
  AO22X1 U451 ( .IN1(n442), .IN2(n484), .IN3(n469), .IN4(n441), .Q(n224) );
  AO22X1 U452 ( .IN1(n442), .IN2(n485), .IN3(n469), .IN4(n484), .Q(n223) );
  AO22X1 U453 ( .IN1(n442), .IN2(n486), .IN3(n469), .IN4(n485), .Q(n222) );
  AO22X1 U454 ( .IN1(n442), .IN2(n487), .IN3(n469), .IN4(n486), .Q(n221) );
  AO22X1 U455 ( .IN1(n442), .IN2(n488), .IN3(n469), .IN4(n487), .Q(n220) );
  AO22X1 U456 ( .IN1(n442), .IN2(n489), .IN3(n469), .IN4(n488), .Q(n219) );
  AO22X1 U457 ( .IN1(n442), .IN2(n490), .IN3(n469), .IN4(n489), .Q(n218) );
  AO22X1 U458 ( .IN1(n442), .IN2(n491), .IN3(n469), .IN4(n490), .Q(n217) );
  XOR2X1 U459 ( .IN1(b[7]), .IN2(a[1]), .Q(n490) );
  AO22X1 U460 ( .IN1(n442), .IN2(n492), .IN3(n469), .IN4(n491), .Q(n216) );
  AO22X1 U461 ( .IN1(n442), .IN2(n493), .IN3(n469), .IN4(n492), .Q(n215) );
  XOR2X1 U462 ( .IN1(b[9]), .IN2(a[1]), .Q(n492) );
  AO22X1 U463 ( .IN1(n442), .IN2(n470), .IN3(n469), .IN4(n493), .Q(n214) );
  XOR2X1 U464 ( .IN1(b[10]), .IN2(a[1]), .Q(n493) );
  XOR2X1 U465 ( .IN1(b[11]), .IN2(a[1]), .Q(n470) );
  NOR2X0 U466 ( .IN1(n494), .IN2(n440), .QN(n212) );
  AO22X1 U467 ( .IN1(n495), .IN2(n463), .IN3(n467), .IN4(n496), .Q(n211) );
  XOR2X1 U468 ( .IN1(n439), .IN2(n444), .Q(n496) );
  AO22X1 U469 ( .IN1(n497), .IN2(n463), .IN3(n467), .IN4(n495), .Q(n210) );
  AO22X1 U470 ( .IN1(n498), .IN2(n463), .IN3(n467), .IN4(n497), .Q(n209) );
  AO22X1 U471 ( .IN1(n499), .IN2(n463), .IN3(n467), .IN4(n498), .Q(n208) );
  AO22X1 U472 ( .IN1(n500), .IN2(n463), .IN3(n467), .IN4(n499), .Q(n207) );
  AO22X1 U473 ( .IN1(n501), .IN2(n463), .IN3(n467), .IN4(n500), .Q(n206) );
  AO22X1 U474 ( .IN1(n502), .IN2(n463), .IN3(n467), .IN4(n501), .Q(n205) );
  AO22X1 U475 ( .IN1(n503), .IN2(n463), .IN3(n467), .IN4(n502), .Q(n204) );
  XOR2X1 U476 ( .IN1(b[7]), .IN2(n444), .Q(n502) );
  AO22X1 U477 ( .IN1(n468), .IN2(n463), .IN3(n467), .IN4(n503), .Q(n203) );
  XOR2X1 U478 ( .IN1(b[9]), .IN2(n444), .Q(n468) );
  OAI21X1 U479 ( .IN1(n463), .IN2(n467), .IN3(n471), .QN(n201) );
  XOR2X1 U480 ( .IN1(b[11]), .IN2(n444), .Q(n471) );
  NOR2X0 U481 ( .IN1(n504), .IN2(n440), .QN(n200) );
  AO22X1 U482 ( .IN1(n505), .IN2(n461), .IN3(n473), .IN4(n506), .Q(n199) );
  XOR2X1 U483 ( .IN1(n439), .IN2(n446), .Q(n506) );
  AO22X1 U484 ( .IN1(n507), .IN2(n461), .IN3(n473), .IN4(n505), .Q(n198) );
  AO22X1 U485 ( .IN1(n508), .IN2(n461), .IN3(n473), .IN4(n507), .Q(n197) );
  AO22X1 U486 ( .IN1(n509), .IN2(n461), .IN3(n473), .IN4(n508), .Q(n196) );
  AO22X1 U487 ( .IN1(n510), .IN2(n461), .IN3(n473), .IN4(n509), .Q(n195) );
  AO22X1 U488 ( .IN1(n511), .IN2(n461), .IN3(n473), .IN4(n510), .Q(n194) );
  AO22X1 U489 ( .IN1(n512), .IN2(n461), .IN3(n473), .IN4(n511), .Q(n193) );
  AO22X1 U490 ( .IN1(n513), .IN2(n461), .IN3(n473), .IN4(n512), .Q(n192) );
  XOR2X1 U491 ( .IN1(b[7]), .IN2(n446), .Q(n512) );
  AO22X1 U492 ( .IN1(n514), .IN2(n461), .IN3(n473), .IN4(n513), .Q(n191) );
  AO22X1 U493 ( .IN1(n474), .IN2(n461), .IN3(n473), .IN4(n514), .Q(n190) );
  XOR2X1 U494 ( .IN1(b[9]), .IN2(n446), .Q(n514) );
  XOR2X1 U495 ( .IN1(b[10]), .IN2(n446), .Q(n474) );
  OAI21X1 U496 ( .IN1(n461), .IN2(n473), .IN3(n472), .QN(n189) );
  XOR2X1 U497 ( .IN1(b[11]), .IN2(n446), .Q(n472) );
  NOR2X0 U498 ( .IN1(n515), .IN2(n440), .QN(n188) );
  AO22X1 U499 ( .IN1(n516), .IN2(n459), .IN3(n476), .IN4(n517), .Q(n187) );
  XOR2X1 U500 ( .IN1(n439), .IN2(n448), .Q(n517) );
  AO22X1 U501 ( .IN1(n518), .IN2(n459), .IN3(n476), .IN4(n516), .Q(n186) );
  AO22X1 U502 ( .IN1(n519), .IN2(n459), .IN3(n476), .IN4(n518), .Q(n185) );
  AO22X1 U503 ( .IN1(n520), .IN2(n459), .IN3(n476), .IN4(n519), .Q(n184) );
  AO22X1 U504 ( .IN1(n521), .IN2(n459), .IN3(n476), .IN4(n520), .Q(n183) );
  AO22X1 U505 ( .IN1(n522), .IN2(n459), .IN3(n476), .IN4(n521), .Q(n182) );
  AO22X1 U506 ( .IN1(n523), .IN2(n459), .IN3(n476), .IN4(n522), .Q(n181) );
  AO22X1 U507 ( .IN1(n524), .IN2(n459), .IN3(n476), .IN4(n523), .Q(n180) );
  XOR2X1 U508 ( .IN1(b[7]), .IN2(n448), .Q(n523) );
  AO22X1 U509 ( .IN1(n525), .IN2(n459), .IN3(n476), .IN4(n524), .Q(n179) );
  AO22X1 U510 ( .IN1(n477), .IN2(n459), .IN3(n476), .IN4(n525), .Q(n178) );
  XOR2X1 U511 ( .IN1(b[9]), .IN2(n448), .Q(n525) );
  XOR2X1 U512 ( .IN1(b[10]), .IN2(n448), .Q(n477) );
  OAI21X1 U513 ( .IN1(n459), .IN2(n476), .IN3(n475), .QN(n177) );
  XOR2X1 U514 ( .IN1(b[11]), .IN2(n448), .Q(n475) );
  NOR2X0 U515 ( .IN1(n526), .IN2(n440), .QN(n176) );
  AO22X1 U516 ( .IN1(n527), .IN2(n457), .IN3(n479), .IN4(n528), .Q(n175) );
  XOR2X1 U517 ( .IN1(n439), .IN2(n450), .Q(n528) );
  AO22X1 U518 ( .IN1(n529), .IN2(n457), .IN3(n479), .IN4(n527), .Q(n174) );
  AO22X1 U519 ( .IN1(n530), .IN2(n457), .IN3(n479), .IN4(n529), .Q(n173) );
  AO22X1 U520 ( .IN1(n531), .IN2(n457), .IN3(n479), .IN4(n530), .Q(n172) );
  AO22X1 U521 ( .IN1(n532), .IN2(n457), .IN3(n479), .IN4(n531), .Q(n171) );
  AO22X1 U522 ( .IN1(n533), .IN2(n457), .IN3(n479), .IN4(n532), .Q(n170) );
  AO22X1 U523 ( .IN1(n534), .IN2(n457), .IN3(n479), .IN4(n533), .Q(n169) );
  AO22X1 U524 ( .IN1(n535), .IN2(n457), .IN3(n479), .IN4(n534), .Q(n168) );
  XOR2X1 U525 ( .IN1(b[7]), .IN2(n450), .Q(n534) );
  AO22X1 U526 ( .IN1(n536), .IN2(n457), .IN3(n479), .IN4(n535), .Q(n167) );
  AO22X1 U527 ( .IN1(n480), .IN2(n457), .IN3(n479), .IN4(n536), .Q(n166) );
  XOR2X1 U528 ( .IN1(b[9]), .IN2(n450), .Q(n536) );
  XOR2X1 U529 ( .IN1(b[10]), .IN2(n450), .Q(n480) );
  OAI21X1 U530 ( .IN1(n457), .IN2(n479), .IN3(n478), .QN(n165) );
  XOR2X1 U531 ( .IN1(b[11]), .IN2(n450), .Q(n478) );
  NOR2X0 U532 ( .IN1(n537), .IN2(n440), .QN(n164) );
  AO22X1 U533 ( .IN1(n538), .IN2(n455), .IN3(n482), .IN4(n539), .Q(n163) );
  XOR2X1 U534 ( .IN1(n439), .IN2(n452), .Q(n539) );
  AO22X1 U535 ( .IN1(n540), .IN2(n455), .IN3(n482), .IN4(n538), .Q(n162) );
  AO22X1 U536 ( .IN1(n541), .IN2(n455), .IN3(n482), .IN4(n540), .Q(n161) );
  AO22X1 U537 ( .IN1(n542), .IN2(n455), .IN3(n482), .IN4(n541), .Q(n160) );
  AO22X1 U538 ( .IN1(n543), .IN2(n455), .IN3(n482), .IN4(n542), .Q(n159) );
  AO22X1 U539 ( .IN1(n544), .IN2(n455), .IN3(n482), .IN4(n543), .Q(n158) );
  AO22X1 U540 ( .IN1(n545), .IN2(n455), .IN3(n482), .IN4(n544), .Q(n157) );
  AO22X1 U541 ( .IN1(n546), .IN2(n455), .IN3(n482), .IN4(n545), .Q(n156) );
  XOR2X1 U542 ( .IN1(b[7]), .IN2(n452), .Q(n545) );
  AO22X1 U543 ( .IN1(n547), .IN2(n455), .IN3(n482), .IN4(n546), .Q(n155) );
  AO22X1 U544 ( .IN1(n483), .IN2(n455), .IN3(n482), .IN4(n547), .Q(n154) );
  XOR2X1 U545 ( .IN1(b[9]), .IN2(n452), .Q(n547) );
  XOR2X1 U546 ( .IN1(b[10]), .IN2(n452), .Q(n483) );
  OAI21X1 U547 ( .IN1(n455), .IN2(n482), .IN3(n481), .QN(n153) );
  XOR2X1 U548 ( .IN1(b[11]), .IN2(n452), .Q(n481) );
  AO21X1 U549 ( .IN1(a[1]), .IN2(n441), .IN3(n469), .Q(n152) );
  AO22X1 U550 ( .IN1(n548), .IN2(n445), .IN3(n467), .IN4(n445), .Q(n151) );
  XOR2X1 U551 ( .IN1(n444), .IN2(a[2]), .Q(n549) );
  NOR2X0 U552 ( .IN1(n439), .IN2(n494), .QN(n548) );
  XNOR2X1 U553 ( .IN1(a[2]), .IN2(a[1]), .Q(n494) );
  AO22X1 U554 ( .IN1(n550), .IN2(n447), .IN3(n473), .IN4(n447), .Q(n150) );
  XOR2X1 U555 ( .IN1(n446), .IN2(a[4]), .Q(n551) );
  NOR2X0 U556 ( .IN1(n439), .IN2(n504), .QN(n550) );
  XNOR2X1 U557 ( .IN1(a[4]), .IN2(n444), .Q(n504) );
  AO22X1 U558 ( .IN1(n552), .IN2(n449), .IN3(n476), .IN4(n449), .Q(n149) );
  XOR2X1 U559 ( .IN1(n448), .IN2(a[6]), .Q(n553) );
  NOR2X0 U560 ( .IN1(n439), .IN2(n515), .QN(n552) );
  XNOR2X1 U561 ( .IN1(a[6]), .IN2(n446), .Q(n515) );
  AO22X1 U562 ( .IN1(n554), .IN2(n451), .IN3(n479), .IN4(n451), .Q(n148) );
  XOR2X1 U563 ( .IN1(n450), .IN2(a[8]), .Q(n555) );
  NOR2X0 U564 ( .IN1(n439), .IN2(n526), .QN(n554) );
  XNOR2X1 U565 ( .IN1(a[8]), .IN2(n448), .Q(n526) );
  AO22X1 U566 ( .IN1(n556), .IN2(n452), .IN3(n482), .IN4(n452), .Q(n147) );
  XOR2X1 U567 ( .IN1(n452), .IN2(a[10]), .Q(n557) );
  NOR2X0 U568 ( .IN1(n439), .IN2(n537), .QN(n556) );
  XNOR2X1 U569 ( .IN1(a[10]), .IN2(n450), .Q(n537) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_4 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;
  wire   n1, n2, n3;
  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_4_DW_mult_tc_0 mult_30 ( .a(in_a), .b({
        in_b[11:8], n3, in_b[6:2], n2, in_b[0]}), .product(pre_out) );
  INVX0 U3 ( .INP(in_b[1]), .ZN(n1) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  NBUFFX4 U5 ( .INP(in_b[7]), .Z(n3) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_1_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [24:0] carry;

  FADDX1 U2_22 ( .A(A[22]), .B(n7), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n8), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n9), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n10), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n11), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n12), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n13), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n18), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n21), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n22), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XNOR3X1 U1 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(DIFF[23]) );
  INVX0 U2 ( .INP(B[21]), .ZN(n8) );
  INVX0 U3 ( .INP(B[20]), .ZN(n9) );
  INVX0 U4 ( .INP(B[22]), .ZN(n7) );
  INVX0 U5 ( .INP(B[19]), .ZN(n10) );
  INVX0 U6 ( .INP(B[18]), .ZN(n11) );
  INVX0 U7 ( .INP(B[17]), .ZN(n12) );
  INVX0 U8 ( .INP(B[16]), .ZN(n13) );
  INVX0 U9 ( .INP(B[15]), .ZN(n14) );
  INVX0 U10 ( .INP(B[14]), .ZN(n15) );
  INVX0 U11 ( .INP(B[13]), .ZN(n16) );
  INVX0 U12 ( .INP(B[12]), .ZN(n17) );
  INVX0 U13 ( .INP(B[11]), .ZN(n18) );
  INVX0 U14 ( .INP(B[10]), .ZN(n19) );
  INVX0 U15 ( .INP(B[9]), .ZN(n20) );
  INVX0 U16 ( .INP(B[8]), .ZN(n21) );
  INVX0 U17 ( .INP(B[7]), .ZN(n22) );
  INVX0 U18 ( .INP(A[3]), .ZN(n4) );
  INVX0 U19 ( .INP(A[1]), .ZN(n6) );
  INVX0 U20 ( .INP(A[5]), .ZN(n2) );
  INVX0 U21 ( .INP(A[2]), .ZN(n5) );
  INVX0 U22 ( .INP(B[0]), .ZN(n23) );
  INVX0 U23 ( .INP(A[4]), .ZN(n3) );
  INVX0 U24 ( .INP(A[6]), .ZN(n1) );
  OAI22X1 U25 ( .IN1(n24), .IN2(n1), .IN3(B[6]), .IN4(n25), .QN(carry[7]) );
  AND2X1 U26 ( .IN1(n1), .IN2(n24), .Q(n25) );
  OA22X1 U27 ( .IN1(n26), .IN2(n2), .IN3(B[5]), .IN4(n27), .Q(n24) );
  AND2X1 U28 ( .IN1(n2), .IN2(n26), .Q(n27) );
  OA22X1 U29 ( .IN1(n28), .IN2(n3), .IN3(B[4]), .IN4(n29), .Q(n26) );
  AND2X1 U30 ( .IN1(n3), .IN2(n28), .Q(n29) );
  OA22X1 U31 ( .IN1(n30), .IN2(n4), .IN3(B[3]), .IN4(n31), .Q(n28) );
  AND2X1 U32 ( .IN1(n4), .IN2(n30), .Q(n31) );
  OA22X1 U33 ( .IN1(n32), .IN2(n5), .IN3(B[2]), .IN4(n33), .Q(n30) );
  AND2X1 U34 ( .IN1(n5), .IN2(n32), .Q(n33) );
  OA22X1 U35 ( .IN1(n34), .IN2(n6), .IN3(B[1]), .IN4(n35), .Q(n32) );
  AND2X1 U36 ( .IN1(n6), .IN2(n34), .Q(n35) );
  NOR2X0 U37 ( .IN1(n23), .IN2(A[0]), .QN(n34) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_1 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_1_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(\output ) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_1_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AO22X1 U1 ( .IN1(A[6]), .IN2(n1), .IN3(B[6]), .IN4(n2), .Q(carry[7]) );
  OR2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AO22X1 U3 ( .IN1(A[5]), .IN2(n3), .IN3(B[5]), .IN4(n4), .Q(n1) );
  OR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AO22X1 U5 ( .IN1(A[4]), .IN2(n5), .IN3(B[4]), .IN4(n6), .Q(n3) );
  OR2X1 U6 ( .IN1(n5), .IN2(A[4]), .Q(n6) );
  AO22X1 U7 ( .IN1(A[3]), .IN2(n7), .IN3(B[3]), .IN4(n8), .Q(n5) );
  OR2X1 U8 ( .IN1(n7), .IN2(A[3]), .Q(n8) );
  AO22X1 U9 ( .IN1(A[2]), .IN2(n9), .IN3(B[2]), .IN4(n10), .Q(n7) );
  OR2X1 U10 ( .IN1(n9), .IN2(A[2]), .Q(n10) );
  AO22X1 U11 ( .IN1(B[1]), .IN2(A[1]), .IN3(n11), .IN4(B[0]), .Q(n9) );
  OA21X1 U12 ( .IN1(A[1]), .IN2(B[1]), .IN3(A[0]), .Q(n11) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_1 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_1_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(\output ) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1 ( a_r, a_i, b_r, b_i, out_r, 
        out_i, clk );
  input [11:0] a_r;
  input [11:0] a_i;
  input [11:0] b_r;
  input [11:0] b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;
  wire   [23:0] mult1_out;
  wire   [23:0] mult2_out;
  wire   [23:0] mult3_out;
  wire   [23:0] mult4_out;
  wire   [23:7] pre_out_r;
  wire   [23:7] pre_out_i;
  wire   [11:0] rnd_out_r;
  wire   [11:0] rnd_out_i;
  wire   [11:0] pos_out_r;
  wire   [11:0] pos_out_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFFX1 \out_r_reg_reg[11]  ( .D(pos_out_r[11]), .CLK(clk), .Q(out_r[11]) );
  DFFX1 \out_r_reg_reg[10]  ( .D(pos_out_r[10]), .CLK(clk), .Q(out_r[10]) );
  DFFX1 \out_r_reg_reg[9]  ( .D(pos_out_r[9]), .CLK(clk), .Q(out_r[9]) );
  DFFX1 \out_r_reg_reg[8]  ( .D(pos_out_r[8]), .CLK(clk), .Q(out_r[8]) );
  DFFX1 \out_r_reg_reg[7]  ( .D(pos_out_r[7]), .CLK(clk), .Q(out_r[7]) );
  DFFX1 \out_r_reg_reg[6]  ( .D(pos_out_r[6]), .CLK(clk), .Q(out_r[6]) );
  DFFX1 \out_r_reg_reg[5]  ( .D(pos_out_r[5]), .CLK(clk), .Q(out_r[5]) );
  DFFX1 \out_r_reg_reg[4]  ( .D(pos_out_r[4]), .CLK(clk), .Q(out_r[4]) );
  DFFX1 \out_r_reg_reg[3]  ( .D(pos_out_r[3]), .CLK(clk), .Q(out_r[3]) );
  DFFX1 \out_r_reg_reg[2]  ( .D(pos_out_r[2]), .CLK(clk), .Q(out_r[2]) );
  DFFX1 \out_r_reg_reg[1]  ( .D(pos_out_r[1]), .CLK(clk), .Q(out_r[1]) );
  DFFX1 \out_r_reg_reg[0]  ( .D(pos_out_r[0]), .CLK(clk), .Q(out_r[0]) );
  DFFX1 \out_i_reg_reg[11]  ( .D(pos_out_i[11]), .CLK(clk), .Q(out_i[11]) );
  DFFX1 \out_i_reg_reg[10]  ( .D(pos_out_i[10]), .CLK(clk), .Q(out_i[10]) );
  DFFX1 \out_i_reg_reg[9]  ( .D(pos_out_i[9]), .CLK(clk), .Q(out_i[9]) );
  DFFX1 \out_i_reg_reg[8]  ( .D(pos_out_i[8]), .CLK(clk), .Q(out_i[8]) );
  DFFX1 \out_i_reg_reg[7]  ( .D(pos_out_i[7]), .CLK(clk), .Q(out_i[7]) );
  DFFX1 \out_i_reg_reg[6]  ( .D(pos_out_i[6]), .CLK(clk), .Q(out_i[6]) );
  DFFX1 \out_i_reg_reg[5]  ( .D(pos_out_i[5]), .CLK(clk), .Q(out_i[5]) );
  DFFX1 \out_i_reg_reg[4]  ( .D(pos_out_i[4]), .CLK(clk), .Q(out_i[4]) );
  DFFX1 \out_i_reg_reg[3]  ( .D(pos_out_i[3]), .CLK(clk), .Q(out_i[3]) );
  DFFX1 \out_i_reg_reg[2]  ( .D(pos_out_i[2]), .CLK(clk), .Q(out_i[2]) );
  DFFX1 \out_i_reg_reg[1]  ( .D(pos_out_i[1]), .CLK(clk), .Q(out_i[1]) );
  DFFX1 \out_i_reg_reg[0]  ( .D(pos_out_i[0]), .CLK(clk), .Q(out_i[0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_7 mult1 ( .in_a({a_r[11:2], n19, a_r[0]}), 
        .in_b({b_r[11], n15, b_r[9:6], n7, b_r[4], n6, b_r[2:1], n2}), .clk(
        clk), .\output (mult1_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_6 mult2 ( .in_a({a_i[11:2], n18, a_i[0]}), 
        .in_b({b_i[11], n12, b_i[9], n16, n14, n13, b_i[5], n4, b_i[3], n17, 
        b_i[1:0]}), .clk(clk), .\output (mult2_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_5 mult3 ( .in_a({a_r[11:2], n19, a_r[0]}), 
        .in_b({b_i[11], n12, b_i[9], n16, n14, n13, b_i[5], n4, b_i[3], n17, 
        b_i[1:0]}), .clk(clk), .\output (mult3_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_4 mult4 ( .in_a({a_i[11:2], n18, a_i[0]}), 
        .in_b({b_r[11], n15, b_r[9:6], n7, b_r[4], n6, b_r[2:1], n2}), .clk(
        clk), .\output (mult4_out) );
  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_1 sub ( .a(mult1_out), .b(mult2_out), .\output ({pre_out_r, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_1 add ( .a(mult3_out), .b(mult4_out), .\output ({pre_out_i, SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_DW01_inc_0 add_154_round ( .A(
        pre_out_i[19:7]), .SUM({rnd_out_i, SYNOPSYS_UNCONNECTED__14}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1_DW01_inc_1 add_140_round ( .A(
        pre_out_r[19:7]), .SUM({rnd_out_r, SYNOPSYS_UNCONNECTED__15}) );
  DELLN2X2 U3 ( .INP(b_r[10]), .Z(n15) );
  DELLN2X2 U4 ( .INP(b_i[6]), .Z(n13) );
  INVX0 U5 ( .INP(b_r[0]), .ZN(n1) );
  INVX0 U6 ( .INP(n1), .ZN(n2) );
  INVX0 U7 ( .INP(b_i[4]), .ZN(n3) );
  INVX1 U8 ( .INP(n3), .ZN(n4) );
  DELLN1X2 U9 ( .INP(b_i[2]), .Z(n17) );
  INVX0 U10 ( .INP(b_r[3]), .ZN(n5) );
  INVX1 U11 ( .INP(n5), .ZN(n6) );
  DELLN2X2 U12 ( .INP(b_r[5]), .Z(n7) );
  INVX0 U13 ( .INP(pre_out_r[23]), .ZN(n42) );
  INVX0 U14 ( .INP(pre_out_i[23]), .ZN(n27) );
  INVX0 U15 ( .INP(n43), .ZN(n45) );
  INVX0 U16 ( .INP(n28), .ZN(n30) );
  AND2X1 U17 ( .IN1(n29), .IN2(n31), .Q(n8) );
  AND2X1 U18 ( .IN1(n44), .IN2(n46), .Q(n9) );
  AND2X1 U19 ( .IN1(n30), .IN2(n31), .Q(n10) );
  AND2X1 U20 ( .IN1(n45), .IN2(n46), .Q(n11) );
  NOR2X0 U21 ( .IN1(pre_out_r[21]), .IN2(pre_out_r[22]), .QN(n35) );
  NOR2X0 U22 ( .IN1(pre_out_i[21]), .IN2(pre_out_i[22]), .QN(n20) );
  NAND2X0 U23 ( .IN1(n36), .IN2(n35), .QN(n38) );
  NOR2X0 U24 ( .IN1(pre_out_r[19]), .IN2(pre_out_r[20]), .QN(n36) );
  NAND2X0 U25 ( .IN1(n21), .IN2(n20), .QN(n23) );
  NOR2X0 U26 ( .IN1(pre_out_i[19]), .IN2(pre_out_i[20]), .QN(n21) );
  INVX0 U27 ( .INP(n33), .ZN(n26) );
  INVX0 U28 ( .INP(n31), .ZN(n32) );
  INVX0 U29 ( .INP(n46), .ZN(n47) );
  INVX0 U30 ( .INP(n48), .ZN(n41) );
  NBUFFX4 U31 ( .INP(b_i[7]), .Z(n14) );
  DELLN1X2 U32 ( .INP(b_i[8]), .Z(n16) );
  DELLN1X2 U33 ( .INP(b_i[10]), .Z(n12) );
  XNOR2X1 U34 ( .IN1(mult3_out[23]), .IN2(mult4_out[23]), .Q(n25) );
  NAND2X0 U35 ( .IN1(n40), .IN2(n39), .QN(n48) );
  DELLN1X2 U36 ( .INP(a_i[1]), .Z(n18) );
  DELLN1X2 U37 ( .INP(a_r[1]), .Z(n19) );
  NAND4X0 U38 ( .IN1(pre_out_i[22]), .IN2(pre_out_i[21]), .IN3(pre_out_i[20]), 
        .IN4(pre_out_i[19]), .QN(n22) );
  MUX21X1 U39 ( .IN1(n23), .IN2(n22), .S(pre_out_i[23]), .Q(n28) );
  XOR2X1 U40 ( .IN1(pre_out_i[23]), .IN2(mult3_out[23]), .Q(n24) );
  NAND2X1 U41 ( .IN1(n25), .IN2(n24), .QN(n33) );
  NAND2X1 U42 ( .IN1(mult3_out[23]), .IN2(n26), .QN(n31) );
  AO21X1 U43 ( .IN1(n28), .IN2(n27), .IN3(n26), .Q(n29) );
  AO21X1 U44 ( .IN1(rnd_out_i[0]), .IN2(n10), .IN3(n8), .Q(pos_out_i[0]) );
  AO21X1 U45 ( .IN1(rnd_out_i[1]), .IN2(n10), .IN3(n8), .Q(pos_out_i[1]) );
  AO21X1 U46 ( .IN1(rnd_out_i[2]), .IN2(n10), .IN3(n8), .Q(pos_out_i[2]) );
  AO21X1 U47 ( .IN1(rnd_out_i[3]), .IN2(n10), .IN3(n8), .Q(pos_out_i[3]) );
  AO21X1 U48 ( .IN1(rnd_out_i[4]), .IN2(n10), .IN3(n8), .Q(pos_out_i[4]) );
  AO21X1 U49 ( .IN1(rnd_out_i[5]), .IN2(n10), .IN3(n8), .Q(pos_out_i[5]) );
  AO21X1 U50 ( .IN1(rnd_out_i[6]), .IN2(n10), .IN3(n8), .Q(pos_out_i[6]) );
  AO21X1 U51 ( .IN1(rnd_out_i[7]), .IN2(n10), .IN3(n8), .Q(pos_out_i[7]) );
  AO21X1 U52 ( .IN1(rnd_out_i[8]), .IN2(n10), .IN3(n8), .Q(pos_out_i[8]) );
  AO21X1 U53 ( .IN1(rnd_out_i[9]), .IN2(n10), .IN3(n8), .Q(pos_out_i[9]) );
  AO21X1 U54 ( .IN1(rnd_out_i[10]), .IN2(n10), .IN3(n8), .Q(pos_out_i[10]) );
  MUX21X1 U55 ( .IN1(pre_out_i[23]), .IN2(rnd_out_i[11]), .S(n30), .Q(n34) );
  AO21X1 U56 ( .IN1(n34), .IN2(n33), .IN3(n32), .Q(pos_out_i[11]) );
  NAND4X0 U57 ( .IN1(pre_out_r[22]), .IN2(pre_out_r[21]), .IN3(pre_out_r[20]), 
        .IN4(pre_out_r[19]), .QN(n37) );
  MUX21X1 U58 ( .IN1(n38), .IN2(n37), .S(pre_out_r[23]), .Q(n43) );
  XOR2X1 U59 ( .IN1(mult2_out[23]), .IN2(mult1_out[23]), .Q(n40) );
  XOR2X1 U60 ( .IN1(pre_out_r[23]), .IN2(mult1_out[23]), .Q(n39) );
  NAND2X1 U61 ( .IN1(mult1_out[23]), .IN2(n41), .QN(n46) );
  AO21X1 U62 ( .IN1(n43), .IN2(n42), .IN3(n41), .Q(n44) );
  AO21X1 U63 ( .IN1(rnd_out_r[0]), .IN2(n11), .IN3(n9), .Q(pos_out_r[0]) );
  AO21X1 U64 ( .IN1(rnd_out_r[1]), .IN2(n11), .IN3(n9), .Q(pos_out_r[1]) );
  AO21X1 U65 ( .IN1(rnd_out_r[2]), .IN2(n11), .IN3(n9), .Q(pos_out_r[2]) );
  AO21X1 U66 ( .IN1(rnd_out_r[3]), .IN2(n11), .IN3(n9), .Q(pos_out_r[3]) );
  AO21X1 U67 ( .IN1(rnd_out_r[4]), .IN2(n11), .IN3(n9), .Q(pos_out_r[4]) );
  AO21X1 U68 ( .IN1(rnd_out_r[5]), .IN2(n11), .IN3(n9), .Q(pos_out_r[5]) );
  AO21X1 U69 ( .IN1(rnd_out_r[6]), .IN2(n11), .IN3(n9), .Q(pos_out_r[6]) );
  AO21X1 U70 ( .IN1(rnd_out_r[7]), .IN2(n11), .IN3(n9), .Q(pos_out_r[7]) );
  AO21X1 U71 ( .IN1(rnd_out_r[8]), .IN2(n11), .IN3(n9), .Q(pos_out_r[8]) );
  AO21X1 U72 ( .IN1(rnd_out_r[9]), .IN2(n11), .IN3(n9), .Q(pos_out_r[9]) );
  AO21X1 U73 ( .IN1(rnd_out_r[10]), .IN2(n11), .IN3(n9), .Q(pos_out_r[10]) );
  MUX21X1 U74 ( .IN1(pre_out_r[23]), .IN2(rnd_out_r[11]), .S(n45), .Q(n49) );
  AO21X1 U75 ( .IN1(n49), .IN2(n48), .IN3(n47), .Q(pos_out_r[11]) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_3_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561;

  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U21 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n23), .B(n151), .CI(n134), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n460), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n462), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n464), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n466), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n120), .CI(n122), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  FADDX1 U311 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  AND3X1 U312 ( .IN1(n414), .IN2(n415), .IN3(n416), .Q(product[23]) );
  DELLN1X2 U313 ( .INP(b[1]), .Z(n409) );
  XOR3X2 U314 ( .IN1(n27), .IN2(n458), .IN3(n5), .Q(product[21]) );
  NAND2X0 U315 ( .IN1(n27), .IN2(n458), .QN(n410) );
  NAND2X0 U316 ( .IN1(n27), .IN2(n5), .QN(n411) );
  NAND2X0 U317 ( .IN1(n458), .IN2(n5), .QN(n412) );
  NAND3X0 U318 ( .IN1(n410), .IN2(n411), .IN3(n412), .QN(n4) );
  XOR2X2 U319 ( .IN1(n25), .IN2(n153), .Q(n413) );
  XOR2X1 U320 ( .IN1(n413), .IN2(n4), .Q(product[22]) );
  NAND2X0 U321 ( .IN1(n25), .IN2(n153), .QN(n414) );
  NAND2X0 U322 ( .IN1(n25), .IN2(n4), .QN(n415) );
  NAND2X0 U323 ( .IN1(n153), .IN2(n4), .QN(n416) );
  XOR3X2 U324 ( .IN1(n118), .IN2(n123), .IN3(n19), .Q(product[7]) );
  NAND2X0 U325 ( .IN1(n118), .IN2(n123), .QN(n417) );
  NAND2X0 U326 ( .IN1(n118), .IN2(n19), .QN(n418) );
  NAND2X0 U327 ( .IN1(n123), .IN2(n19), .QN(n419) );
  NAND3X0 U328 ( .IN1(n417), .IN2(n418), .IN3(n419), .QN(n18) );
  XOR2X2 U329 ( .IN1(n112), .IN2(n117), .Q(n420) );
  XOR2X1 U330 ( .IN1(n420), .IN2(n18), .Q(product[8]) );
  NAND2X0 U331 ( .IN1(n112), .IN2(n117), .QN(n421) );
  NAND2X0 U332 ( .IN1(n112), .IN2(n18), .QN(n422) );
  NAND2X0 U333 ( .IN1(n117), .IN2(n18), .QN(n423) );
  NAND3X0 U334 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n17) );
  XOR2X2 U335 ( .IN1(n127), .IN2(n124), .Q(n424) );
  XOR2X1 U336 ( .IN1(n424), .IN2(n20), .Q(product[6]) );
  NAND2X0 U337 ( .IN1(n124), .IN2(n20), .QN(n425) );
  NAND2X0 U338 ( .IN1(n127), .IN2(n20), .QN(n426) );
  NAND2X0 U339 ( .IN1(n127), .IN2(n124), .QN(n427) );
  NAND3X0 U340 ( .IN1(n425), .IN2(n427), .IN3(n426), .QN(n19) );
  XOR2X2 U341 ( .IN1(b[9]), .IN2(n457), .Q(n551) );
  XOR2X2 U342 ( .IN1(b[9]), .IN2(n455), .Q(n540) );
  XOR2X2 U343 ( .IN1(b[9]), .IN2(n453), .Q(n529) );
  XOR2X2 U344 ( .IN1(b[9]), .IN2(n451), .Q(n518) );
  XOR2X2 U345 ( .IN1(b[9]), .IN2(n449), .Q(n472) );
  XOR2X2 U346 ( .IN1(b[9]), .IN2(n443), .Q(n496) );
  XOR2X2 U347 ( .IN1(b[6]), .IN2(n457), .Q(n548) );
  XOR2X2 U348 ( .IN1(b[6]), .IN2(n455), .Q(n537) );
  XOR2X2 U349 ( .IN1(b[6]), .IN2(n453), .Q(n526) );
  XOR2X2 U350 ( .IN1(b[6]), .IN2(n451), .Q(n515) );
  XOR2X2 U351 ( .IN1(b[6]), .IN2(n449), .Q(n505) );
  XOR2X2 U352 ( .IN1(b[6]), .IN2(n443), .Q(n493) );
  XNOR2X2 U353 ( .IN1(n10), .IN2(n428), .Q(product[16]) );
  XNOR2X2 U354 ( .IN1(n6), .IN2(n429), .Q(product[20]) );
  XOR2X2 U355 ( .IN1(b[8]), .IN2(n457), .Q(n550) );
  XOR2X2 U356 ( .IN1(b[8]), .IN2(n455), .Q(n539) );
  XOR2X2 U357 ( .IN1(b[8]), .IN2(n453), .Q(n528) );
  XOR2X2 U358 ( .IN1(b[8]), .IN2(n451), .Q(n517) );
  XOR2X2 U359 ( .IN1(b[8]), .IN2(n449), .Q(n507) );
  XOR2X2 U360 ( .IN1(b[8]), .IN2(n443), .Q(n495) );
  XOR2X2 U361 ( .IN1(b[4]), .IN2(n457), .Q(n546) );
  XOR2X2 U362 ( .IN1(b[4]), .IN2(n455), .Q(n535) );
  XOR2X2 U363 ( .IN1(b[4]), .IN2(n453), .Q(n524) );
  XOR2X2 U364 ( .IN1(b[4]), .IN2(n451), .Q(n513) );
  XOR2X2 U365 ( .IN1(b[4]), .IN2(n449), .Q(n503) );
  XOR2X2 U366 ( .IN1(b[4]), .IN2(n443), .Q(n491) );
  XOR2X2 U367 ( .IN1(b[3]), .IN2(n457), .Q(n545) );
  XOR2X2 U368 ( .IN1(b[3]), .IN2(n455), .Q(n534) );
  XOR2X2 U369 ( .IN1(b[3]), .IN2(n453), .Q(n523) );
  XOR2X2 U370 ( .IN1(b[3]), .IN2(n451), .Q(n512) );
  XOR2X2 U371 ( .IN1(b[3]), .IN2(n449), .Q(n502) );
  XOR2X2 U372 ( .IN1(b[3]), .IN2(n443), .Q(n490) );
  XOR3X1 U373 ( .IN1(n57), .IN2(n50), .IN3(n11), .Q(product[15]) );
  XNOR2X1 U374 ( .IN1(n49), .IN2(n44), .Q(n428) );
  INVX0 U375 ( .INP(n25), .ZN(n458) );
  INVX0 U376 ( .INP(n55), .ZN(n464) );
  XOR3X1 U377 ( .IN1(n33), .IN2(n30), .IN3(n7), .Q(product[19]) );
  XNOR2X1 U378 ( .IN1(n29), .IN2(n28), .Q(n429) );
  XOR2X1 U379 ( .IN1(b[2]), .IN2(n443), .Q(n489) );
  XOR2X1 U380 ( .IN1(n409), .IN2(n443), .Q(n488) );
  XOR2X1 U381 ( .IN1(n409), .IN2(n449), .Q(n499) );
  XOR2X1 U382 ( .IN1(n409), .IN2(n451), .Q(n509) );
  XOR2X1 U383 ( .IN1(n409), .IN2(n453), .Q(n520) );
  INVX0 U384 ( .INP(n73), .ZN(n466) );
  XOR2X1 U385 ( .IN1(n409), .IN2(n455), .Q(n531) );
  XOR2X1 U386 ( .IN1(n409), .IN2(n457), .Q(n542) );
  INVX0 U387 ( .INP(n41), .ZN(n462) );
  NBUFFX2 U388 ( .INP(a[1]), .Z(n443) );
  AND2X1 U389 ( .IN1(n443), .IN2(n448), .Q(n473) );
  INVX0 U390 ( .INP(n31), .ZN(n460) );
  INVX0 U391 ( .INP(n498), .ZN(n467) );
  INVX0 U392 ( .INP(n508), .ZN(n465) );
  INVX0 U393 ( .INP(n519), .ZN(n463) );
  INVX0 U394 ( .INP(n530), .ZN(n461) );
  INVX0 U395 ( .INP(n541), .ZN(n459) );
  NBUFFX2 U396 ( .INP(a[3]), .Z(n450) );
  NBUFFX2 U397 ( .INP(a[5]), .Z(n452) );
  NBUFFX2 U398 ( .INP(b[5]), .Z(n430) );
  AND2X1 U399 ( .IN1(n498), .IN2(n553), .Q(n471) );
  AND2X1 U400 ( .IN1(n519), .IN2(n557), .Q(n480) );
  AND2X1 U401 ( .IN1(n508), .IN2(n555), .Q(n477) );
  AND2X1 U402 ( .IN1(n530), .IN2(n559), .Q(n483) );
  AND2X1 U403 ( .IN1(n541), .IN2(n561), .Q(n486) );
  NBUFFX2 U404 ( .INP(a[7]), .Z(n454) );
  NBUFFX2 U405 ( .INP(a[9]), .Z(n456) );
  NAND2X0 U406 ( .IN1(n33), .IN2(n30), .QN(n431) );
  NAND2X0 U407 ( .IN1(n33), .IN2(n7), .QN(n432) );
  NAND2X0 U408 ( .IN1(n30), .IN2(n7), .QN(n433) );
  NAND3X0 U409 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(n6) );
  NAND2X0 U410 ( .IN1(n29), .IN2(n28), .QN(n434) );
  NAND2X0 U411 ( .IN1(n29), .IN2(n6), .QN(n435) );
  NAND2X0 U412 ( .IN1(n28), .IN2(n6), .QN(n436) );
  NAND3X0 U413 ( .IN1(n436), .IN2(n435), .IN3(n434), .QN(n5) );
  NAND2X0 U414 ( .IN1(n57), .IN2(n50), .QN(n437) );
  NAND2X0 U415 ( .IN1(n57), .IN2(n11), .QN(n438) );
  NAND2X0 U416 ( .IN1(n50), .IN2(n11), .QN(n439) );
  NAND3X0 U417 ( .IN1(n437), .IN2(n438), .IN3(n439), .QN(n10) );
  NAND2X0 U418 ( .IN1(n49), .IN2(n44), .QN(n440) );
  NAND2X0 U419 ( .IN1(n49), .IN2(n10), .QN(n441) );
  NAND2X0 U420 ( .IN1(n44), .IN2(n10), .QN(n442) );
  NAND3X0 U421 ( .IN1(n442), .IN2(n441), .IN3(n440), .QN(n9) );
  DELLN1X2 U422 ( .INP(a[11]), .Z(n457) );
  INVX0 U423 ( .INP(n446), .ZN(n444) );
  INVX0 U424 ( .INP(b[0]), .ZN(n445) );
  INVX0 U425 ( .INP(b[0]), .ZN(n446) );
  INVX0 U426 ( .INP(n448), .ZN(n447) );
  INVX0 U427 ( .INP(a[0]), .ZN(n448) );
  DELLN1X2 U428 ( .INP(a[3]), .Z(n449) );
  DELLN1X2 U429 ( .INP(a[5]), .Z(n451) );
  DELLN1X2 U430 ( .INP(a[7]), .Z(n453) );
  DELLN1X2 U431 ( .INP(a[9]), .Z(n455) );
  NOR2X0 U432 ( .IN1(n448), .IN2(n446), .QN(product[0]) );
  XNOR2X1 U433 ( .IN1(n468), .IN2(n469), .Q(n84) );
  NAND2X0 U434 ( .IN1(n469), .IN2(n468), .QN(n83) );
  AOI22X1 U435 ( .IN1(n470), .IN2(n467), .IN3(n471), .IN4(n472), .QN(n468) );
  OA21X1 U436 ( .IN1(n473), .IN2(n447), .IN3(n474), .Q(n469) );
  AO22X1 U437 ( .IN1(n475), .IN2(n467), .IN3(n471), .IN4(n470), .Q(n73) );
  XOR2X1 U438 ( .IN1(b[10]), .IN2(n449), .Q(n470) );
  AO22X1 U439 ( .IN1(n476), .IN2(n465), .IN3(n477), .IN4(n478), .Q(n55) );
  AO22X1 U440 ( .IN1(n479), .IN2(n463), .IN3(n480), .IN4(n481), .Q(n41) );
  AO22X1 U441 ( .IN1(n482), .IN2(n461), .IN3(n483), .IN4(n484), .Q(n31) );
  AO22X1 U442 ( .IN1(n485), .IN2(n459), .IN3(n486), .IN4(n487), .Q(n25) );
  AO22X1 U443 ( .IN1(n447), .IN2(n488), .IN3(n473), .IN4(n445), .Q(n224) );
  AO22X1 U444 ( .IN1(n447), .IN2(n489), .IN3(n473), .IN4(n488), .Q(n223) );
  AO22X1 U445 ( .IN1(n447), .IN2(n490), .IN3(n473), .IN4(n489), .Q(n222) );
  AO22X1 U446 ( .IN1(n447), .IN2(n491), .IN3(n473), .IN4(n490), .Q(n221) );
  AO22X1 U447 ( .IN1(n447), .IN2(n492), .IN3(n473), .IN4(n491), .Q(n220) );
  AO22X1 U448 ( .IN1(n447), .IN2(n493), .IN3(n473), .IN4(n492), .Q(n219) );
  XOR2X1 U449 ( .IN1(n430), .IN2(n443), .Q(n492) );
  AO22X1 U450 ( .IN1(n447), .IN2(n494), .IN3(n473), .IN4(n493), .Q(n218) );
  AO22X1 U451 ( .IN1(n447), .IN2(n495), .IN3(n473), .IN4(n494), .Q(n217) );
  XOR2X1 U452 ( .IN1(b[7]), .IN2(n443), .Q(n494) );
  AO22X1 U453 ( .IN1(n447), .IN2(n496), .IN3(n473), .IN4(n495), .Q(n216) );
  AO22X1 U454 ( .IN1(n447), .IN2(n497), .IN3(n473), .IN4(n496), .Q(n215) );
  AO22X1 U455 ( .IN1(n447), .IN2(n474), .IN3(n473), .IN4(n497), .Q(n214) );
  XOR2X1 U456 ( .IN1(b[10]), .IN2(n443), .Q(n497) );
  XOR2X1 U457 ( .IN1(b[11]), .IN2(n443), .Q(n474) );
  NOR2X0 U458 ( .IN1(n498), .IN2(n446), .QN(n212) );
  AO22X1 U459 ( .IN1(n499), .IN2(n467), .IN3(n471), .IN4(n500), .Q(n211) );
  XOR2X1 U460 ( .IN1(n444), .IN2(n449), .Q(n500) );
  AO22X1 U461 ( .IN1(n501), .IN2(n467), .IN3(n471), .IN4(n499), .Q(n210) );
  AO22X1 U462 ( .IN1(n502), .IN2(n467), .IN3(n471), .IN4(n501), .Q(n209) );
  XOR2X1 U463 ( .IN1(b[2]), .IN2(n449), .Q(n501) );
  AO22X1 U464 ( .IN1(n503), .IN2(n467), .IN3(n471), .IN4(n502), .Q(n208) );
  AO22X1 U465 ( .IN1(n504), .IN2(n467), .IN3(n471), .IN4(n503), .Q(n207) );
  AO22X1 U466 ( .IN1(n505), .IN2(n467), .IN3(n471), .IN4(n504), .Q(n206) );
  XOR2X1 U467 ( .IN1(n430), .IN2(n449), .Q(n504) );
  AO22X1 U468 ( .IN1(n506), .IN2(n467), .IN3(n471), .IN4(n505), .Q(n205) );
  AO22X1 U469 ( .IN1(n507), .IN2(n467), .IN3(n471), .IN4(n506), .Q(n204) );
  XOR2X1 U470 ( .IN1(b[7]), .IN2(n449), .Q(n506) );
  AO22X1 U471 ( .IN1(n472), .IN2(n467), .IN3(n471), .IN4(n507), .Q(n203) );
  OAI21X1 U472 ( .IN1(n467), .IN2(n471), .IN3(n475), .QN(n201) );
  XOR2X1 U473 ( .IN1(b[11]), .IN2(n449), .Q(n475) );
  NOR2X0 U474 ( .IN1(n508), .IN2(n446), .QN(n200) );
  AO22X1 U475 ( .IN1(n509), .IN2(n465), .IN3(n477), .IN4(n510), .Q(n199) );
  XOR2X1 U476 ( .IN1(n444), .IN2(n451), .Q(n510) );
  AO22X1 U477 ( .IN1(n511), .IN2(n465), .IN3(n477), .IN4(n509), .Q(n198) );
  AO22X1 U478 ( .IN1(n512), .IN2(n465), .IN3(n477), .IN4(n511), .Q(n197) );
  XOR2X1 U479 ( .IN1(b[2]), .IN2(n451), .Q(n511) );
  AO22X1 U480 ( .IN1(n513), .IN2(n465), .IN3(n477), .IN4(n512), .Q(n196) );
  AO22X1 U481 ( .IN1(n514), .IN2(n465), .IN3(n477), .IN4(n513), .Q(n195) );
  AO22X1 U482 ( .IN1(n515), .IN2(n465), .IN3(n477), .IN4(n514), .Q(n194) );
  XOR2X1 U483 ( .IN1(n430), .IN2(n451), .Q(n514) );
  AO22X1 U484 ( .IN1(n516), .IN2(n465), .IN3(n477), .IN4(n515), .Q(n193) );
  AO22X1 U485 ( .IN1(n517), .IN2(n465), .IN3(n477), .IN4(n516), .Q(n192) );
  XOR2X1 U486 ( .IN1(b[7]), .IN2(n451), .Q(n516) );
  AO22X1 U487 ( .IN1(n518), .IN2(n465), .IN3(n477), .IN4(n517), .Q(n191) );
  AO22X1 U488 ( .IN1(n478), .IN2(n465), .IN3(n477), .IN4(n518), .Q(n190) );
  XOR2X1 U489 ( .IN1(b[10]), .IN2(n451), .Q(n478) );
  OAI21X1 U490 ( .IN1(n465), .IN2(n477), .IN3(n476), .QN(n189) );
  XOR2X1 U491 ( .IN1(b[11]), .IN2(n451), .Q(n476) );
  NOR2X0 U492 ( .IN1(n519), .IN2(n445), .QN(n188) );
  AO22X1 U493 ( .IN1(n520), .IN2(n463), .IN3(n480), .IN4(n521), .Q(n187) );
  XOR2X1 U494 ( .IN1(n444), .IN2(n453), .Q(n521) );
  AO22X1 U495 ( .IN1(n522), .IN2(n463), .IN3(n480), .IN4(n520), .Q(n186) );
  AO22X1 U496 ( .IN1(n523), .IN2(n463), .IN3(n480), .IN4(n522), .Q(n185) );
  XOR2X1 U497 ( .IN1(b[2]), .IN2(n453), .Q(n522) );
  AO22X1 U498 ( .IN1(n524), .IN2(n463), .IN3(n480), .IN4(n523), .Q(n184) );
  AO22X1 U499 ( .IN1(n525), .IN2(n463), .IN3(n480), .IN4(n524), .Q(n183) );
  AO22X1 U500 ( .IN1(n526), .IN2(n463), .IN3(n480), .IN4(n525), .Q(n182) );
  XOR2X1 U501 ( .IN1(n430), .IN2(n453), .Q(n525) );
  AO22X1 U502 ( .IN1(n527), .IN2(n463), .IN3(n480), .IN4(n526), .Q(n181) );
  AO22X1 U503 ( .IN1(n528), .IN2(n463), .IN3(n480), .IN4(n527), .Q(n180) );
  XOR2X1 U504 ( .IN1(b[7]), .IN2(n453), .Q(n527) );
  AO22X1 U505 ( .IN1(n529), .IN2(n463), .IN3(n480), .IN4(n528), .Q(n179) );
  AO22X1 U506 ( .IN1(n481), .IN2(n463), .IN3(n480), .IN4(n529), .Q(n178) );
  XOR2X1 U507 ( .IN1(b[10]), .IN2(n453), .Q(n481) );
  OAI21X1 U508 ( .IN1(n463), .IN2(n480), .IN3(n479), .QN(n177) );
  XOR2X1 U509 ( .IN1(b[11]), .IN2(n453), .Q(n479) );
  NOR2X0 U510 ( .IN1(n530), .IN2(n445), .QN(n176) );
  AO22X1 U511 ( .IN1(n531), .IN2(n461), .IN3(n483), .IN4(n532), .Q(n175) );
  XOR2X1 U512 ( .IN1(n444), .IN2(n455), .Q(n532) );
  AO22X1 U513 ( .IN1(n533), .IN2(n461), .IN3(n483), .IN4(n531), .Q(n174) );
  AO22X1 U514 ( .IN1(n534), .IN2(n461), .IN3(n483), .IN4(n533), .Q(n173) );
  XOR2X1 U515 ( .IN1(b[2]), .IN2(n455), .Q(n533) );
  AO22X1 U516 ( .IN1(n535), .IN2(n461), .IN3(n483), .IN4(n534), .Q(n172) );
  AO22X1 U517 ( .IN1(n536), .IN2(n461), .IN3(n483), .IN4(n535), .Q(n171) );
  AO22X1 U518 ( .IN1(n537), .IN2(n461), .IN3(n483), .IN4(n536), .Q(n170) );
  XOR2X1 U519 ( .IN1(n430), .IN2(n455), .Q(n536) );
  AO22X1 U520 ( .IN1(n538), .IN2(n461), .IN3(n483), .IN4(n537), .Q(n169) );
  AO22X1 U521 ( .IN1(n539), .IN2(n461), .IN3(n483), .IN4(n538), .Q(n168) );
  XOR2X1 U522 ( .IN1(b[7]), .IN2(n455), .Q(n538) );
  AO22X1 U523 ( .IN1(n540), .IN2(n461), .IN3(n483), .IN4(n539), .Q(n167) );
  AO22X1 U524 ( .IN1(n484), .IN2(n461), .IN3(n483), .IN4(n540), .Q(n166) );
  XOR2X1 U525 ( .IN1(b[10]), .IN2(n455), .Q(n484) );
  OAI21X1 U526 ( .IN1(n461), .IN2(n483), .IN3(n482), .QN(n165) );
  XOR2X1 U527 ( .IN1(b[11]), .IN2(n455), .Q(n482) );
  NOR2X0 U528 ( .IN1(n541), .IN2(n445), .QN(n164) );
  AO22X1 U529 ( .IN1(n542), .IN2(n459), .IN3(n486), .IN4(n543), .Q(n163) );
  XOR2X1 U530 ( .IN1(n444), .IN2(n457), .Q(n543) );
  AO22X1 U531 ( .IN1(n544), .IN2(n459), .IN3(n486), .IN4(n542), .Q(n162) );
  AO22X1 U532 ( .IN1(n545), .IN2(n459), .IN3(n486), .IN4(n544), .Q(n161) );
  XOR2X1 U533 ( .IN1(b[2]), .IN2(n457), .Q(n544) );
  AO22X1 U534 ( .IN1(n546), .IN2(n459), .IN3(n486), .IN4(n545), .Q(n160) );
  AO22X1 U535 ( .IN1(n547), .IN2(n459), .IN3(n486), .IN4(n546), .Q(n159) );
  AO22X1 U536 ( .IN1(n548), .IN2(n459), .IN3(n486), .IN4(n547), .Q(n158) );
  XOR2X1 U537 ( .IN1(n430), .IN2(n457), .Q(n547) );
  AO22X1 U538 ( .IN1(n549), .IN2(n459), .IN3(n486), .IN4(n548), .Q(n157) );
  AO22X1 U539 ( .IN1(n550), .IN2(n459), .IN3(n486), .IN4(n549), .Q(n156) );
  XOR2X1 U540 ( .IN1(b[7]), .IN2(n457), .Q(n549) );
  AO22X1 U541 ( .IN1(n551), .IN2(n459), .IN3(n486), .IN4(n550), .Q(n155) );
  AO22X1 U542 ( .IN1(n487), .IN2(n459), .IN3(n486), .IN4(n551), .Q(n154) );
  XOR2X1 U543 ( .IN1(b[10]), .IN2(n457), .Q(n487) );
  OAI21X1 U544 ( .IN1(n459), .IN2(n486), .IN3(n485), .QN(n153) );
  XOR2X1 U545 ( .IN1(b[11]), .IN2(n457), .Q(n485) );
  AO21X1 U546 ( .IN1(n443), .IN2(n445), .IN3(n473), .Q(n152) );
  AO22X1 U547 ( .IN1(n552), .IN2(n450), .IN3(n471), .IN4(n450), .Q(n151) );
  XOR2X1 U548 ( .IN1(n449), .IN2(a[2]), .Q(n553) );
  NOR2X0 U549 ( .IN1(n444), .IN2(n498), .QN(n552) );
  XNOR2X1 U550 ( .IN1(a[2]), .IN2(n443), .Q(n498) );
  AO22X1 U551 ( .IN1(n554), .IN2(n452), .IN3(n477), .IN4(n452), .Q(n150) );
  XOR2X1 U552 ( .IN1(n451), .IN2(a[4]), .Q(n555) );
  NOR2X0 U553 ( .IN1(n444), .IN2(n508), .QN(n554) );
  XNOR2X1 U554 ( .IN1(a[4]), .IN2(n449), .Q(n508) );
  AO22X1 U555 ( .IN1(n556), .IN2(n454), .IN3(n480), .IN4(n454), .Q(n149) );
  XOR2X1 U556 ( .IN1(n453), .IN2(a[6]), .Q(n557) );
  NOR2X0 U557 ( .IN1(n444), .IN2(n519), .QN(n556) );
  XNOR2X1 U558 ( .IN1(a[6]), .IN2(n451), .Q(n519) );
  AO22X1 U559 ( .IN1(n558), .IN2(n456), .IN3(n483), .IN4(n456), .Q(n148) );
  XOR2X1 U560 ( .IN1(n455), .IN2(a[8]), .Q(n559) );
  NOR2X0 U561 ( .IN1(n444), .IN2(n530), .QN(n558) );
  XNOR2X1 U562 ( .IN1(a[8]), .IN2(n453), .Q(n530) );
  AO22X1 U563 ( .IN1(n560), .IN2(n457), .IN3(n486), .IN4(n457), .Q(n147) );
  XOR2X1 U564 ( .IN1(n457), .IN2(a[10]), .Q(n561) );
  NOR2X0 U565 ( .IN1(n444), .IN2(n541), .QN(n560) );
  XNOR2X1 U566 ( .IN1(a[10]), .IN2(n455), .Q(n541) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_3 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_3_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_2_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n450), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U19 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n452), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n454), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n456), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n458), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n200), .B(n221), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  INVX0 U311 ( .INP(b[11]), .ZN(n408) );
  INVX0 U312 ( .INP(n408), .ZN(n409) );
  XOR2X1 U313 ( .IN1(n435), .IN2(n440), .Q(n492) );
  INVX0 U314 ( .INP(b[4]), .ZN(n410) );
  INVX0 U315 ( .INP(n410), .ZN(n411) );
  DELLN2X2 U316 ( .INP(n7), .Z(n412) );
  INVX0 U317 ( .INP(n437), .ZN(n413) );
  INVX0 U318 ( .INP(n437), .ZN(n414) );
  DELLN2X2 U319 ( .INP(n13), .Z(n415) );
  XOR2X2 U320 ( .IN1(n413), .IN2(n448), .Q(n535) );
  XOR2X2 U321 ( .IN1(n413), .IN2(n446), .Q(n524) );
  XOR2X2 U322 ( .IN1(n414), .IN2(n444), .Q(n513) );
  XOR2X2 U323 ( .IN1(n413), .IN2(n442), .Q(n502) );
  INVX0 U324 ( .INP(b[3]), .ZN(n416) );
  INVX0 U325 ( .INP(n416), .ZN(n417) );
  INVX0 U326 ( .INP(b[1]), .ZN(n418) );
  INVX0 U327 ( .INP(n418), .ZN(n419) );
  XOR2X2 U328 ( .IN1(n409), .IN2(n448), .Q(n477) );
  XOR2X2 U329 ( .IN1(n409), .IN2(n446), .Q(n474) );
  XOR2X2 U330 ( .IN1(n409), .IN2(n444), .Q(n471) );
  XOR2X2 U331 ( .IN1(n409), .IN2(n442), .Q(n468) );
  XOR2X2 U332 ( .IN1(n409), .IN2(n440), .Q(n467) );
  XOR2X2 U333 ( .IN1(n409), .IN2(n434), .Q(n466) );
  XOR2X2 U334 ( .IN1(n411), .IN2(n448), .Q(n538) );
  XOR2X2 U335 ( .IN1(n411), .IN2(n446), .Q(n527) );
  XOR2X2 U336 ( .IN1(n411), .IN2(n444), .Q(n516) );
  XOR2X2 U337 ( .IN1(n411), .IN2(n442), .Q(n505) );
  XOR2X2 U338 ( .IN1(n411), .IN2(n440), .Q(n495) );
  XOR2X2 U339 ( .IN1(n411), .IN2(n434), .Q(n483) );
  XOR3X1 U340 ( .IN1(n37), .IN2(n34), .IN3(n8), .Q(product[18]) );
  XOR3X1 U341 ( .IN1(n76), .IN2(n85), .IN3(n14), .Q(product[12]) );
  XNOR2X1 U342 ( .IN1(n420), .IN2(n415), .Q(product[13]) );
  XNOR2X1 U343 ( .IN1(n66), .IN2(n75), .Q(n420) );
  FADDX1 U344 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  INVX0 U345 ( .INP(n25), .ZN(n450) );
  INVX0 U346 ( .INP(n3), .ZN(product[23]) );
  INVX0 U347 ( .INP(n55), .ZN(n456) );
  XNOR2X1 U348 ( .IN1(n421), .IN2(n412), .Q(product[19]) );
  XNOR2X1 U349 ( .IN1(n33), .IN2(n30), .Q(n421) );
  XOR2X1 U350 ( .IN1(n419), .IN2(n434), .Q(n480) );
  XOR2X1 U351 ( .IN1(n417), .IN2(n434), .Q(n482) );
  XOR2X1 U352 ( .IN1(n419), .IN2(n440), .Q(n491) );
  XOR2X1 U353 ( .IN1(n419), .IN2(n442), .Q(n501) );
  XOR2X1 U354 ( .IN1(n419), .IN2(n444), .Q(n512) );
  XOR2X1 U355 ( .IN1(n417), .IN2(n440), .Q(n494) );
  XOR2X1 U356 ( .IN1(n417), .IN2(n442), .Q(n504) );
  INVX0 U357 ( .INP(n73), .ZN(n458) );
  FADDX1 U358 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U359 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X1 U360 ( .IN1(n419), .IN2(n446), .Q(n523) );
  XOR2X1 U361 ( .IN1(n419), .IN2(n448), .Q(n534) );
  XOR2X1 U362 ( .IN1(n417), .IN2(n444), .Q(n515) );
  XOR2X1 U363 ( .IN1(n417), .IN2(n446), .Q(n526) );
  INVX0 U364 ( .INP(n41), .ZN(n454) );
  INVX0 U365 ( .INP(n31), .ZN(n452) );
  XOR2X1 U366 ( .IN1(n417), .IN2(n448), .Q(n537) );
  XOR2X1 U367 ( .IN1(b[2]), .IN2(n434), .Q(n481) );
  NBUFFX2 U368 ( .INP(a[1]), .Z(n434) );
  INVX0 U369 ( .INP(n490), .ZN(n459) );
  AND2X1 U370 ( .IN1(n434), .IN2(n439), .Q(n465) );
  INVX0 U371 ( .INP(n500), .ZN(n457) );
  INVX0 U372 ( .INP(n511), .ZN(n455) );
  INVX0 U373 ( .INP(n522), .ZN(n453) );
  INVX0 U374 ( .INP(n533), .ZN(n451) );
  NBUFFX2 U375 ( .INP(a[5]), .Z(n443) );
  FADDX1 U376 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  NBUFFX2 U377 ( .INP(a[3]), .Z(n441) );
  AND2X1 U378 ( .IN1(n490), .IN2(n545), .Q(n463) );
  AND2X1 U379 ( .IN1(n511), .IN2(n549), .Q(n472) );
  AND2X1 U380 ( .IN1(n500), .IN2(n547), .Q(n469) );
  AND2X1 U381 ( .IN1(n522), .IN2(n551), .Q(n475) );
  AND2X1 U382 ( .IN1(n533), .IN2(n553), .Q(n478) );
  NBUFFX2 U383 ( .INP(a[7]), .Z(n445) );
  NBUFFX2 U384 ( .INP(a[9]), .Z(n447) );
  NAND2X0 U385 ( .IN1(n37), .IN2(n34), .QN(n422) );
  NAND2X0 U386 ( .IN1(n37), .IN2(n8), .QN(n423) );
  NAND2X0 U387 ( .IN1(n34), .IN2(n8), .QN(n424) );
  NAND3X0 U388 ( .IN1(n422), .IN2(n423), .IN3(n424), .QN(n7) );
  NAND2X0 U389 ( .IN1(n33), .IN2(n30), .QN(n425) );
  NAND2X0 U390 ( .IN1(n33), .IN2(n7), .QN(n426) );
  NAND2X0 U391 ( .IN1(n30), .IN2(n7), .QN(n427) );
  NAND3X0 U392 ( .IN1(n425), .IN2(n426), .IN3(n427), .QN(n6) );
  NAND2X0 U393 ( .IN1(n76), .IN2(n85), .QN(n428) );
  NAND2X0 U394 ( .IN1(n76), .IN2(n14), .QN(n429) );
  NAND2X0 U395 ( .IN1(n85), .IN2(n14), .QN(n430) );
  NAND3X0 U396 ( .IN1(n428), .IN2(n429), .IN3(n430), .QN(n13) );
  NAND2X0 U397 ( .IN1(n66), .IN2(n75), .QN(n431) );
  NAND2X0 U398 ( .IN1(n66), .IN2(n13), .QN(n432) );
  NAND2X0 U399 ( .IN1(n75), .IN2(n13), .QN(n433) );
  NAND3X0 U400 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(n12) );
  DELLN1X2 U401 ( .INP(a[11]), .Z(n448) );
  INVX0 U402 ( .INP(n437), .ZN(n435) );
  INVX0 U403 ( .INP(b[0]), .ZN(n436) );
  INVX0 U404 ( .INP(b[0]), .ZN(n437) );
  INVX0 U405 ( .INP(n439), .ZN(n438) );
  INVX0 U406 ( .INP(a[0]), .ZN(n439) );
  DELLN1X2 U407 ( .INP(a[3]), .Z(n440) );
  DELLN1X2 U408 ( .INP(a[5]), .Z(n442) );
  DELLN1X2 U409 ( .INP(a[7]), .Z(n444) );
  DELLN1X2 U410 ( .INP(a[9]), .Z(n446) );
  NOR2X0 U411 ( .IN1(n439), .IN2(n436), .QN(product[0]) );
  XNOR2X1 U412 ( .IN1(n460), .IN2(n461), .Q(n84) );
  NAND2X0 U413 ( .IN1(n461), .IN2(n460), .QN(n83) );
  AOI22X1 U414 ( .IN1(n462), .IN2(n459), .IN3(n463), .IN4(n464), .QN(n460) );
  OA21X1 U415 ( .IN1(n465), .IN2(n438), .IN3(n466), .Q(n461) );
  AO22X1 U416 ( .IN1(n467), .IN2(n459), .IN3(n463), .IN4(n462), .Q(n73) );
  XOR2X1 U417 ( .IN1(b[10]), .IN2(n440), .Q(n462) );
  AO22X1 U418 ( .IN1(n468), .IN2(n457), .IN3(n469), .IN4(n470), .Q(n55) );
  AO22X1 U419 ( .IN1(n471), .IN2(n455), .IN3(n472), .IN4(n473), .Q(n41) );
  AO22X1 U420 ( .IN1(n474), .IN2(n453), .IN3(n475), .IN4(n476), .Q(n31) );
  AO22X1 U421 ( .IN1(n477), .IN2(n451), .IN3(n478), .IN4(n479), .Q(n25) );
  AO22X1 U422 ( .IN1(n438), .IN2(n480), .IN3(n465), .IN4(n437), .Q(n224) );
  AO22X1 U423 ( .IN1(n438), .IN2(n481), .IN3(n465), .IN4(n480), .Q(n223) );
  AO22X1 U424 ( .IN1(n438), .IN2(n482), .IN3(n465), .IN4(n481), .Q(n222) );
  AO22X1 U425 ( .IN1(n438), .IN2(n483), .IN3(n465), .IN4(n482), .Q(n221) );
  AO22X1 U426 ( .IN1(n438), .IN2(n484), .IN3(n465), .IN4(n483), .Q(n220) );
  AO22X1 U427 ( .IN1(n438), .IN2(n485), .IN3(n465), .IN4(n484), .Q(n219) );
  XOR2X1 U428 ( .IN1(b[5]), .IN2(n434), .Q(n484) );
  AO22X1 U429 ( .IN1(n438), .IN2(n486), .IN3(n465), .IN4(n485), .Q(n218) );
  XOR2X1 U430 ( .IN1(b[6]), .IN2(n434), .Q(n485) );
  AO22X1 U431 ( .IN1(n438), .IN2(n487), .IN3(n465), .IN4(n486), .Q(n217) );
  XOR2X1 U432 ( .IN1(b[7]), .IN2(n434), .Q(n486) );
  AO22X1 U433 ( .IN1(n438), .IN2(n488), .IN3(n465), .IN4(n487), .Q(n216) );
  XOR2X1 U434 ( .IN1(b[8]), .IN2(n434), .Q(n487) );
  AO22X1 U435 ( .IN1(n438), .IN2(n489), .IN3(n465), .IN4(n488), .Q(n215) );
  XOR2X1 U436 ( .IN1(b[9]), .IN2(n434), .Q(n488) );
  AO22X1 U437 ( .IN1(n438), .IN2(n466), .IN3(n465), .IN4(n489), .Q(n214) );
  XOR2X1 U438 ( .IN1(b[10]), .IN2(n434), .Q(n489) );
  NOR2X0 U439 ( .IN1(n490), .IN2(n436), .QN(n212) );
  AO22X1 U440 ( .IN1(n491), .IN2(n459), .IN3(n463), .IN4(n492), .Q(n211) );
  AO22X1 U441 ( .IN1(n493), .IN2(n459), .IN3(n463), .IN4(n491), .Q(n210) );
  AO22X1 U442 ( .IN1(n494), .IN2(n459), .IN3(n463), .IN4(n493), .Q(n209) );
  XOR2X1 U443 ( .IN1(b[2]), .IN2(n440), .Q(n493) );
  AO22X1 U444 ( .IN1(n495), .IN2(n459), .IN3(n463), .IN4(n494), .Q(n208) );
  AO22X1 U445 ( .IN1(n496), .IN2(n459), .IN3(n463), .IN4(n495), .Q(n207) );
  AO22X1 U446 ( .IN1(n497), .IN2(n459), .IN3(n463), .IN4(n496), .Q(n206) );
  XOR2X1 U447 ( .IN1(b[5]), .IN2(n440), .Q(n496) );
  AO22X1 U448 ( .IN1(n498), .IN2(n459), .IN3(n463), .IN4(n497), .Q(n205) );
  XOR2X1 U449 ( .IN1(b[6]), .IN2(n440), .Q(n497) );
  AO22X1 U450 ( .IN1(n499), .IN2(n459), .IN3(n463), .IN4(n498), .Q(n204) );
  XOR2X1 U451 ( .IN1(b[7]), .IN2(n440), .Q(n498) );
  AO22X1 U452 ( .IN1(n464), .IN2(n459), .IN3(n463), .IN4(n499), .Q(n203) );
  XOR2X1 U453 ( .IN1(b[8]), .IN2(n440), .Q(n499) );
  XOR2X1 U454 ( .IN1(b[9]), .IN2(n440), .Q(n464) );
  OAI21X1 U455 ( .IN1(n459), .IN2(n463), .IN3(n467), .QN(n201) );
  NOR2X0 U456 ( .IN1(n500), .IN2(n436), .QN(n200) );
  AO22X1 U457 ( .IN1(n501), .IN2(n457), .IN3(n469), .IN4(n502), .Q(n199) );
  AO22X1 U458 ( .IN1(n503), .IN2(n457), .IN3(n469), .IN4(n501), .Q(n198) );
  AO22X1 U459 ( .IN1(n504), .IN2(n457), .IN3(n469), .IN4(n503), .Q(n197) );
  XOR2X1 U460 ( .IN1(b[2]), .IN2(n442), .Q(n503) );
  AO22X1 U461 ( .IN1(n505), .IN2(n457), .IN3(n469), .IN4(n504), .Q(n196) );
  AO22X1 U462 ( .IN1(n506), .IN2(n457), .IN3(n469), .IN4(n505), .Q(n195) );
  AO22X1 U463 ( .IN1(n507), .IN2(n457), .IN3(n469), .IN4(n506), .Q(n194) );
  XOR2X1 U464 ( .IN1(b[5]), .IN2(n442), .Q(n506) );
  AO22X1 U465 ( .IN1(n508), .IN2(n457), .IN3(n469), .IN4(n507), .Q(n193) );
  XOR2X1 U466 ( .IN1(b[6]), .IN2(n442), .Q(n507) );
  AO22X1 U467 ( .IN1(n509), .IN2(n457), .IN3(n469), .IN4(n508), .Q(n192) );
  XOR2X1 U468 ( .IN1(b[7]), .IN2(n442), .Q(n508) );
  AO22X1 U469 ( .IN1(n510), .IN2(n457), .IN3(n469), .IN4(n509), .Q(n191) );
  XOR2X1 U470 ( .IN1(b[8]), .IN2(n442), .Q(n509) );
  AO22X1 U471 ( .IN1(n470), .IN2(n457), .IN3(n469), .IN4(n510), .Q(n190) );
  XOR2X1 U472 ( .IN1(b[9]), .IN2(n442), .Q(n510) );
  XOR2X1 U473 ( .IN1(b[10]), .IN2(n442), .Q(n470) );
  OAI21X1 U474 ( .IN1(n457), .IN2(n469), .IN3(n468), .QN(n189) );
  NOR2X0 U475 ( .IN1(n511), .IN2(n436), .QN(n188) );
  AO22X1 U476 ( .IN1(n512), .IN2(n455), .IN3(n472), .IN4(n513), .Q(n187) );
  AO22X1 U477 ( .IN1(n514), .IN2(n455), .IN3(n472), .IN4(n512), .Q(n186) );
  AO22X1 U478 ( .IN1(n515), .IN2(n455), .IN3(n472), .IN4(n514), .Q(n185) );
  XOR2X1 U479 ( .IN1(b[2]), .IN2(n444), .Q(n514) );
  AO22X1 U480 ( .IN1(n516), .IN2(n455), .IN3(n472), .IN4(n515), .Q(n184) );
  AO22X1 U481 ( .IN1(n517), .IN2(n455), .IN3(n472), .IN4(n516), .Q(n183) );
  AO22X1 U482 ( .IN1(n518), .IN2(n455), .IN3(n472), .IN4(n517), .Q(n182) );
  XOR2X1 U483 ( .IN1(b[5]), .IN2(n444), .Q(n517) );
  AO22X1 U484 ( .IN1(n519), .IN2(n455), .IN3(n472), .IN4(n518), .Q(n181) );
  XOR2X1 U485 ( .IN1(b[6]), .IN2(n444), .Q(n518) );
  AO22X1 U486 ( .IN1(n520), .IN2(n455), .IN3(n472), .IN4(n519), .Q(n180) );
  XOR2X1 U487 ( .IN1(b[7]), .IN2(n444), .Q(n519) );
  AO22X1 U488 ( .IN1(n521), .IN2(n455), .IN3(n472), .IN4(n520), .Q(n179) );
  XOR2X1 U489 ( .IN1(b[8]), .IN2(n444), .Q(n520) );
  AO22X1 U490 ( .IN1(n473), .IN2(n455), .IN3(n472), .IN4(n521), .Q(n178) );
  XOR2X1 U491 ( .IN1(b[9]), .IN2(n444), .Q(n521) );
  XOR2X1 U492 ( .IN1(b[10]), .IN2(n444), .Q(n473) );
  OAI21X1 U493 ( .IN1(n455), .IN2(n472), .IN3(n471), .QN(n177) );
  NOR2X0 U494 ( .IN1(n522), .IN2(n436), .QN(n176) );
  AO22X1 U495 ( .IN1(n523), .IN2(n453), .IN3(n475), .IN4(n524), .Q(n175) );
  AO22X1 U496 ( .IN1(n525), .IN2(n453), .IN3(n475), .IN4(n523), .Q(n174) );
  AO22X1 U497 ( .IN1(n526), .IN2(n453), .IN3(n475), .IN4(n525), .Q(n173) );
  XOR2X1 U498 ( .IN1(b[2]), .IN2(n446), .Q(n525) );
  AO22X1 U499 ( .IN1(n527), .IN2(n453), .IN3(n475), .IN4(n526), .Q(n172) );
  AO22X1 U500 ( .IN1(n528), .IN2(n453), .IN3(n475), .IN4(n527), .Q(n171) );
  AO22X1 U501 ( .IN1(n529), .IN2(n453), .IN3(n475), .IN4(n528), .Q(n170) );
  XOR2X1 U502 ( .IN1(b[5]), .IN2(n446), .Q(n528) );
  AO22X1 U503 ( .IN1(n530), .IN2(n453), .IN3(n475), .IN4(n529), .Q(n169) );
  XOR2X1 U504 ( .IN1(b[6]), .IN2(n446), .Q(n529) );
  AO22X1 U505 ( .IN1(n531), .IN2(n453), .IN3(n475), .IN4(n530), .Q(n168) );
  XOR2X1 U506 ( .IN1(b[7]), .IN2(n446), .Q(n530) );
  AO22X1 U507 ( .IN1(n532), .IN2(n453), .IN3(n475), .IN4(n531), .Q(n167) );
  XOR2X1 U508 ( .IN1(b[8]), .IN2(n446), .Q(n531) );
  AO22X1 U509 ( .IN1(n476), .IN2(n453), .IN3(n475), .IN4(n532), .Q(n166) );
  XOR2X1 U510 ( .IN1(b[9]), .IN2(n446), .Q(n532) );
  XOR2X1 U511 ( .IN1(b[10]), .IN2(n446), .Q(n476) );
  OAI21X1 U512 ( .IN1(n453), .IN2(n475), .IN3(n474), .QN(n165) );
  NOR2X0 U513 ( .IN1(n533), .IN2(n436), .QN(n164) );
  AO22X1 U514 ( .IN1(n534), .IN2(n451), .IN3(n478), .IN4(n535), .Q(n163) );
  AO22X1 U515 ( .IN1(n536), .IN2(n451), .IN3(n478), .IN4(n534), .Q(n162) );
  AO22X1 U516 ( .IN1(n537), .IN2(n451), .IN3(n478), .IN4(n536), .Q(n161) );
  XOR2X1 U517 ( .IN1(b[2]), .IN2(n448), .Q(n536) );
  AO22X1 U518 ( .IN1(n538), .IN2(n451), .IN3(n478), .IN4(n537), .Q(n160) );
  AO22X1 U519 ( .IN1(n539), .IN2(n451), .IN3(n478), .IN4(n538), .Q(n159) );
  AO22X1 U520 ( .IN1(n540), .IN2(n451), .IN3(n478), .IN4(n539), .Q(n158) );
  XOR2X1 U521 ( .IN1(b[5]), .IN2(n448), .Q(n539) );
  AO22X1 U522 ( .IN1(n541), .IN2(n451), .IN3(n478), .IN4(n540), .Q(n157) );
  XOR2X1 U523 ( .IN1(b[6]), .IN2(n448), .Q(n540) );
  AO22X1 U524 ( .IN1(n542), .IN2(n451), .IN3(n478), .IN4(n541), .Q(n156) );
  XOR2X1 U525 ( .IN1(b[7]), .IN2(n448), .Q(n541) );
  AO22X1 U526 ( .IN1(n543), .IN2(n451), .IN3(n478), .IN4(n542), .Q(n155) );
  XOR2X1 U527 ( .IN1(b[8]), .IN2(n448), .Q(n542) );
  AO22X1 U528 ( .IN1(n479), .IN2(n451), .IN3(n478), .IN4(n543), .Q(n154) );
  XOR2X1 U529 ( .IN1(b[9]), .IN2(n448), .Q(n543) );
  XOR2X1 U530 ( .IN1(b[10]), .IN2(n448), .Q(n479) );
  OAI21X1 U531 ( .IN1(n451), .IN2(n478), .IN3(n477), .QN(n153) );
  AO21X1 U532 ( .IN1(n434), .IN2(n437), .IN3(n465), .Q(n152) );
  AO22X1 U533 ( .IN1(n544), .IN2(n441), .IN3(n463), .IN4(n441), .Q(n151) );
  XOR2X1 U534 ( .IN1(n440), .IN2(a[2]), .Q(n545) );
  NOR2X0 U535 ( .IN1(n414), .IN2(n490), .QN(n544) );
  XNOR2X1 U536 ( .IN1(a[2]), .IN2(n434), .Q(n490) );
  AO22X1 U537 ( .IN1(n546), .IN2(n443), .IN3(n469), .IN4(n443), .Q(n150) );
  XOR2X1 U538 ( .IN1(n442), .IN2(a[4]), .Q(n547) );
  NOR2X0 U539 ( .IN1(n414), .IN2(n500), .QN(n546) );
  XNOR2X1 U540 ( .IN1(a[4]), .IN2(n440), .Q(n500) );
  AO22X1 U541 ( .IN1(n548), .IN2(n445), .IN3(n472), .IN4(n445), .Q(n149) );
  XOR2X1 U542 ( .IN1(n444), .IN2(a[6]), .Q(n549) );
  NOR2X0 U543 ( .IN1(n413), .IN2(n511), .QN(n548) );
  XNOR2X1 U544 ( .IN1(a[6]), .IN2(n442), .Q(n511) );
  AO22X1 U545 ( .IN1(n550), .IN2(n447), .IN3(n475), .IN4(n447), .Q(n148) );
  XOR2X1 U546 ( .IN1(n446), .IN2(a[8]), .Q(n551) );
  NOR2X0 U547 ( .IN1(n414), .IN2(n522), .QN(n550) );
  XNOR2X1 U548 ( .IN1(a[8]), .IN2(n444), .Q(n522) );
  AO22X1 U549 ( .IN1(n552), .IN2(n448), .IN3(n478), .IN4(n448), .Q(n147) );
  XOR2X1 U550 ( .IN1(n448), .IN2(a[10]), .Q(n553) );
  NOR2X0 U551 ( .IN1(n414), .IN2(n533), .QN(n552) );
  XNOR2X1 U552 ( .IN1(a[10]), .IN2(n446), .Q(n533) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_2 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_2_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_1_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n449), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U16 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  FADDX1 U18 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n451), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n453), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n455), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n457), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n221), .B(n200), .CI(n210), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  DELLN1X2 U311 ( .INP(b[1]), .Z(n408) );
  INVX0 U312 ( .INP(b[5]), .ZN(n409) );
  INVX0 U313 ( .INP(n409), .ZN(n410) );
  INVX0 U314 ( .INP(b[11]), .ZN(n411) );
  INVX0 U315 ( .INP(n411), .ZN(n412) );
  XOR2X2 U316 ( .IN1(n412), .IN2(n447), .Q(n476) );
  XOR2X2 U317 ( .IN1(n412), .IN2(n445), .Q(n473) );
  XOR2X2 U318 ( .IN1(n412), .IN2(n443), .Q(n470) );
  XOR2X2 U319 ( .IN1(n412), .IN2(n441), .Q(n467) );
  XOR2X2 U320 ( .IN1(n412), .IN2(n439), .Q(n466) );
  XOR2X2 U321 ( .IN1(n412), .IN2(a[1]), .Q(n465) );
  XOR2X2 U322 ( .IN1(b[4]), .IN2(n447), .Q(n537) );
  XOR2X2 U323 ( .IN1(b[4]), .IN2(n445), .Q(n526) );
  XOR2X2 U324 ( .IN1(b[4]), .IN2(n443), .Q(n515) );
  XOR2X2 U325 ( .IN1(b[4]), .IN2(n441), .Q(n504) );
  XOR3X1 U326 ( .IN1(n66), .IN2(n75), .IN3(n13), .Q(product[13]) );
  NAND2X0 U327 ( .IN1(n66), .IN2(n75), .QN(n413) );
  NAND2X0 U328 ( .IN1(n65), .IN2(n58), .QN(n417) );
  XOR2X1 U329 ( .IN1(n132), .IN2(n133), .Q(n430) );
  NAND2X0 U330 ( .IN1(n151), .IN2(n23), .QN(n429) );
  NAND2X0 U331 ( .IN1(n66), .IN2(n13), .QN(n414) );
  NAND2X0 U332 ( .IN1(n75), .IN2(n13), .QN(n415) );
  NAND3X0 U333 ( .IN1(n413), .IN2(n414), .IN3(n415), .QN(n12) );
  XOR2X1 U334 ( .IN1(n65), .IN2(n58), .Q(n416) );
  XOR2X1 U335 ( .IN1(n416), .IN2(n12), .Q(product[14]) );
  NAND2X0 U336 ( .IN1(n65), .IN2(n12), .QN(n418) );
  NAND2X0 U337 ( .IN1(n58), .IN2(n12), .QN(n419) );
  NAND3X0 U338 ( .IN1(n417), .IN2(n418), .IN3(n419), .QN(n11) );
  XOR3X1 U339 ( .IN1(n124), .IN2(n127), .IN3(n20), .Q(product[6]) );
  NAND2X0 U340 ( .IN1(n124), .IN2(n127), .QN(n420) );
  NAND2X0 U341 ( .IN1(n124), .IN2(n20), .QN(n421) );
  NAND2X0 U342 ( .IN1(n127), .IN2(n20), .QN(n422) );
  NAND3X0 U343 ( .IN1(n420), .IN2(n421), .IN3(n422), .QN(n19) );
  XOR2X1 U344 ( .IN1(n118), .IN2(n123), .Q(n423) );
  XOR2X1 U345 ( .IN1(n423), .IN2(n19), .Q(product[7]) );
  NAND2X0 U346 ( .IN1(n118), .IN2(n123), .QN(n424) );
  NAND2X0 U347 ( .IN1(n118), .IN2(n19), .QN(n425) );
  NAND2X0 U348 ( .IN1(n123), .IN2(n19), .QN(n426) );
  NAND3X0 U349 ( .IN1(n424), .IN2(n425), .IN3(n426), .QN(n18) );
  XOR3X1 U350 ( .IN1(n134), .IN2(n151), .IN3(n23), .Q(product[3]) );
  NAND2X0 U351 ( .IN1(n134), .IN2(n151), .QN(n427) );
  NAND2X0 U352 ( .IN1(n134), .IN2(n23), .QN(n428) );
  NAND3X0 U353 ( .IN1(n427), .IN2(n428), .IN3(n429), .QN(n22) );
  XOR2X1 U354 ( .IN1(n430), .IN2(n22), .Q(product[4]) );
  NAND2X0 U355 ( .IN1(n132), .IN2(n133), .QN(n431) );
  NAND2X0 U356 ( .IN1(n132), .IN2(n22), .QN(n432) );
  NAND2X0 U357 ( .IN1(n133), .IN2(n22), .QN(n433) );
  NAND3X0 U358 ( .IN1(n431), .IN2(n432), .IN3(n433), .QN(n21) );
  FADDX1 U359 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U360 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  INVX0 U361 ( .INP(n25), .ZN(n449) );
  FADDX1 U362 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  INVX0 U363 ( .INP(n3), .ZN(product[23]) );
  INVX0 U364 ( .INP(n55), .ZN(n455) );
  XOR2X1 U365 ( .IN1(n408), .IN2(n439), .Q(n490) );
  INVX0 U366 ( .INP(n73), .ZN(n457) );
  XOR2X1 U367 ( .IN1(n408), .IN2(n445), .Q(n522) );
  XOR2X1 U368 ( .IN1(n408), .IN2(n443), .Q(n511) );
  XOR2X1 U369 ( .IN1(n408), .IN2(n441), .Q(n500) );
  XOR2X1 U370 ( .IN1(b[3]), .IN2(n443), .Q(n514) );
  XOR2X1 U371 ( .IN1(b[3]), .IN2(n441), .Q(n503) );
  XOR2X1 U372 ( .IN1(b[3]), .IN2(n439), .Q(n493) );
  XOR2X1 U373 ( .IN1(n408), .IN2(n447), .Q(n533) );
  XOR2X1 U374 ( .IN1(b[3]), .IN2(n447), .Q(n536) );
  INVX0 U375 ( .INP(n31), .ZN(n451) );
  INVX0 U376 ( .INP(n41), .ZN(n453) );
  XOR2X1 U377 ( .IN1(b[2]), .IN2(a[1]), .Q(n480) );
  XOR2X1 U378 ( .IN1(b[2]), .IN2(n439), .Q(n492) );
  INVX0 U379 ( .INP(n499), .ZN(n456) );
  INVX0 U380 ( .INP(n489), .ZN(n458) );
  AND2X1 U381 ( .IN1(a[1]), .IN2(n438), .Q(n464) );
  INVX0 U382 ( .INP(n521), .ZN(n452) );
  INVX0 U383 ( .INP(n510), .ZN(n454) );
  INVX0 U384 ( .INP(n532), .ZN(n450) );
  NBUFFX2 U385 ( .INP(a[3]), .Z(n440) );
  NBUFFX2 U386 ( .INP(a[5]), .Z(n442) );
  XOR2X1 U387 ( .IN1(n410), .IN2(a[1]), .Q(n483) );
  NBUFFX2 U388 ( .INP(a[7]), .Z(n444) );
  NBUFFX2 U389 ( .INP(a[9]), .Z(n446) );
  XOR2X2 U390 ( .IN1(b[4]), .IN2(n439), .Q(n494) );
  XOR2X2 U391 ( .IN1(b[4]), .IN2(a[1]), .Q(n482) );
  XOR2X2 U392 ( .IN1(b[3]), .IN2(n445), .Q(n525) );
  XOR2X2 U393 ( .IN1(b[3]), .IN2(a[1]), .Q(n481) );
  XOR2X2 U394 ( .IN1(n408), .IN2(a[1]), .Q(n479) );
  XOR2X2 U395 ( .IN1(b[10]), .IN2(a[1]), .Q(n488) );
  XOR2X2 U396 ( .IN1(b[8]), .IN2(a[1]), .Q(n486) );
  XOR2X2 U397 ( .IN1(b[7]), .IN2(a[1]), .Q(n485) );
  FADDX1 U398 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  FADDX1 U399 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  DELLN1X2 U400 ( .INP(a[11]), .Z(n447) );
  AND2X2 U401 ( .IN1(n489), .IN2(n544), .Q(n462) );
  AND2X2 U402 ( .IN1(n499), .IN2(n546), .Q(n468) );
  AND2X2 U403 ( .IN1(n510), .IN2(n548), .Q(n471) );
  AND2X2 U404 ( .IN1(n521), .IN2(n550), .Q(n474) );
  AND2X2 U405 ( .IN1(n532), .IN2(n552), .Q(n477) );
  INVX0 U406 ( .INP(n436), .ZN(n434) );
  INVX0 U407 ( .INP(b[0]), .ZN(n435) );
  INVX0 U408 ( .INP(b[0]), .ZN(n436) );
  INVX0 U409 ( .INP(n438), .ZN(n437) );
  INVX0 U410 ( .INP(a[0]), .ZN(n438) );
  DELLN1X2 U411 ( .INP(a[3]), .Z(n439) );
  DELLN1X2 U412 ( .INP(a[5]), .Z(n441) );
  DELLN1X2 U413 ( .INP(a[7]), .Z(n443) );
  DELLN1X2 U414 ( .INP(a[9]), .Z(n445) );
  NOR2X0 U415 ( .IN1(n438), .IN2(n435), .QN(product[0]) );
  XNOR2X1 U416 ( .IN1(n459), .IN2(n460), .Q(n84) );
  NAND2X0 U417 ( .IN1(n460), .IN2(n459), .QN(n83) );
  AOI22X1 U418 ( .IN1(n461), .IN2(n458), .IN3(n462), .IN4(n463), .QN(n459) );
  OA21X1 U419 ( .IN1(n464), .IN2(n437), .IN3(n465), .Q(n460) );
  AO22X1 U420 ( .IN1(n466), .IN2(n458), .IN3(n462), .IN4(n461), .Q(n73) );
  XOR2X1 U421 ( .IN1(b[10]), .IN2(n439), .Q(n461) );
  AO22X1 U422 ( .IN1(n467), .IN2(n456), .IN3(n468), .IN4(n469), .Q(n55) );
  AO22X1 U423 ( .IN1(n470), .IN2(n454), .IN3(n471), .IN4(n472), .Q(n41) );
  AO22X1 U424 ( .IN1(n473), .IN2(n452), .IN3(n474), .IN4(n475), .Q(n31) );
  AO22X1 U425 ( .IN1(n476), .IN2(n450), .IN3(n477), .IN4(n478), .Q(n25) );
  AO22X1 U426 ( .IN1(n437), .IN2(n479), .IN3(n464), .IN4(n436), .Q(n224) );
  AO22X1 U427 ( .IN1(n437), .IN2(n480), .IN3(n464), .IN4(n479), .Q(n223) );
  AO22X1 U428 ( .IN1(n437), .IN2(n481), .IN3(n464), .IN4(n480), .Q(n222) );
  AO22X1 U429 ( .IN1(n437), .IN2(n482), .IN3(n464), .IN4(n481), .Q(n221) );
  AO22X1 U430 ( .IN1(n437), .IN2(n483), .IN3(n464), .IN4(n482), .Q(n220) );
  AO22X1 U431 ( .IN1(n437), .IN2(n484), .IN3(n464), .IN4(n483), .Q(n219) );
  AO22X1 U432 ( .IN1(n437), .IN2(n485), .IN3(n464), .IN4(n484), .Q(n218) );
  XOR2X1 U433 ( .IN1(b[6]), .IN2(a[1]), .Q(n484) );
  AO22X1 U434 ( .IN1(n437), .IN2(n486), .IN3(n464), .IN4(n485), .Q(n217) );
  AO22X1 U435 ( .IN1(n437), .IN2(n487), .IN3(n464), .IN4(n486), .Q(n216) );
  AO22X1 U436 ( .IN1(n437), .IN2(n488), .IN3(n464), .IN4(n487), .Q(n215) );
  XOR2X1 U437 ( .IN1(b[9]), .IN2(a[1]), .Q(n487) );
  AO22X1 U438 ( .IN1(n437), .IN2(n465), .IN3(n464), .IN4(n488), .Q(n214) );
  NOR2X0 U439 ( .IN1(n489), .IN2(n435), .QN(n212) );
  AO22X1 U440 ( .IN1(n490), .IN2(n458), .IN3(n462), .IN4(n491), .Q(n211) );
  XOR2X1 U441 ( .IN1(n434), .IN2(n439), .Q(n491) );
  AO22X1 U442 ( .IN1(n492), .IN2(n458), .IN3(n462), .IN4(n490), .Q(n210) );
  AO22X1 U443 ( .IN1(n493), .IN2(n458), .IN3(n462), .IN4(n492), .Q(n209) );
  AO22X1 U444 ( .IN1(n494), .IN2(n458), .IN3(n462), .IN4(n493), .Q(n208) );
  AO22X1 U445 ( .IN1(n495), .IN2(n458), .IN3(n462), .IN4(n494), .Q(n207) );
  AO22X1 U446 ( .IN1(n496), .IN2(n458), .IN3(n462), .IN4(n495), .Q(n206) );
  XOR2X1 U447 ( .IN1(n410), .IN2(n439), .Q(n495) );
  AO22X1 U448 ( .IN1(n497), .IN2(n458), .IN3(n462), .IN4(n496), .Q(n205) );
  XOR2X1 U449 ( .IN1(b[6]), .IN2(n439), .Q(n496) );
  AO22X1 U450 ( .IN1(n498), .IN2(n458), .IN3(n462), .IN4(n497), .Q(n204) );
  XOR2X1 U451 ( .IN1(b[7]), .IN2(n439), .Q(n497) );
  AO22X1 U452 ( .IN1(n463), .IN2(n458), .IN3(n462), .IN4(n498), .Q(n203) );
  XOR2X1 U453 ( .IN1(b[8]), .IN2(n439), .Q(n498) );
  XOR2X1 U454 ( .IN1(b[9]), .IN2(n439), .Q(n463) );
  OAI21X1 U455 ( .IN1(n458), .IN2(n462), .IN3(n466), .QN(n201) );
  NOR2X0 U456 ( .IN1(n499), .IN2(n435), .QN(n200) );
  AO22X1 U457 ( .IN1(n500), .IN2(n456), .IN3(n468), .IN4(n501), .Q(n199) );
  XOR2X1 U458 ( .IN1(n434), .IN2(n441), .Q(n501) );
  AO22X1 U459 ( .IN1(n502), .IN2(n456), .IN3(n468), .IN4(n500), .Q(n198) );
  AO22X1 U460 ( .IN1(n503), .IN2(n456), .IN3(n468), .IN4(n502), .Q(n197) );
  XOR2X1 U461 ( .IN1(b[2]), .IN2(n441), .Q(n502) );
  AO22X1 U462 ( .IN1(n504), .IN2(n456), .IN3(n468), .IN4(n503), .Q(n196) );
  AO22X1 U463 ( .IN1(n505), .IN2(n456), .IN3(n468), .IN4(n504), .Q(n195) );
  AO22X1 U464 ( .IN1(n506), .IN2(n456), .IN3(n468), .IN4(n505), .Q(n194) );
  XOR2X1 U465 ( .IN1(n410), .IN2(n441), .Q(n505) );
  AO22X1 U466 ( .IN1(n507), .IN2(n456), .IN3(n468), .IN4(n506), .Q(n193) );
  XOR2X1 U467 ( .IN1(b[6]), .IN2(n441), .Q(n506) );
  AO22X1 U468 ( .IN1(n508), .IN2(n456), .IN3(n468), .IN4(n507), .Q(n192) );
  XOR2X1 U469 ( .IN1(b[7]), .IN2(n441), .Q(n507) );
  AO22X1 U470 ( .IN1(n509), .IN2(n456), .IN3(n468), .IN4(n508), .Q(n191) );
  XOR2X1 U471 ( .IN1(b[8]), .IN2(n441), .Q(n508) );
  AO22X1 U472 ( .IN1(n469), .IN2(n456), .IN3(n468), .IN4(n509), .Q(n190) );
  XOR2X1 U473 ( .IN1(b[9]), .IN2(n441), .Q(n509) );
  XOR2X1 U474 ( .IN1(b[10]), .IN2(n441), .Q(n469) );
  OAI21X1 U475 ( .IN1(n456), .IN2(n468), .IN3(n467), .QN(n189) );
  NOR2X0 U476 ( .IN1(n510), .IN2(n435), .QN(n188) );
  AO22X1 U477 ( .IN1(n511), .IN2(n454), .IN3(n471), .IN4(n512), .Q(n187) );
  XOR2X1 U478 ( .IN1(n434), .IN2(n443), .Q(n512) );
  AO22X1 U479 ( .IN1(n513), .IN2(n454), .IN3(n471), .IN4(n511), .Q(n186) );
  AO22X1 U480 ( .IN1(n514), .IN2(n454), .IN3(n471), .IN4(n513), .Q(n185) );
  XOR2X1 U481 ( .IN1(b[2]), .IN2(n443), .Q(n513) );
  AO22X1 U482 ( .IN1(n515), .IN2(n454), .IN3(n471), .IN4(n514), .Q(n184) );
  AO22X1 U483 ( .IN1(n516), .IN2(n454), .IN3(n471), .IN4(n515), .Q(n183) );
  AO22X1 U484 ( .IN1(n517), .IN2(n454), .IN3(n471), .IN4(n516), .Q(n182) );
  XOR2X1 U485 ( .IN1(n410), .IN2(n443), .Q(n516) );
  AO22X1 U486 ( .IN1(n518), .IN2(n454), .IN3(n471), .IN4(n517), .Q(n181) );
  XOR2X1 U487 ( .IN1(b[6]), .IN2(n443), .Q(n517) );
  AO22X1 U488 ( .IN1(n519), .IN2(n454), .IN3(n471), .IN4(n518), .Q(n180) );
  XOR2X1 U489 ( .IN1(b[7]), .IN2(n443), .Q(n518) );
  AO22X1 U490 ( .IN1(n520), .IN2(n454), .IN3(n471), .IN4(n519), .Q(n179) );
  XOR2X1 U491 ( .IN1(b[8]), .IN2(n443), .Q(n519) );
  AO22X1 U492 ( .IN1(n472), .IN2(n454), .IN3(n471), .IN4(n520), .Q(n178) );
  XOR2X1 U493 ( .IN1(b[9]), .IN2(n443), .Q(n520) );
  XOR2X1 U494 ( .IN1(b[10]), .IN2(n443), .Q(n472) );
  OAI21X1 U495 ( .IN1(n454), .IN2(n471), .IN3(n470), .QN(n177) );
  NOR2X0 U496 ( .IN1(n521), .IN2(n435), .QN(n176) );
  AO22X1 U497 ( .IN1(n522), .IN2(n452), .IN3(n474), .IN4(n523), .Q(n175) );
  XOR2X1 U498 ( .IN1(n434), .IN2(n445), .Q(n523) );
  AO22X1 U499 ( .IN1(n524), .IN2(n452), .IN3(n474), .IN4(n522), .Q(n174) );
  AO22X1 U500 ( .IN1(n525), .IN2(n452), .IN3(n474), .IN4(n524), .Q(n173) );
  XOR2X1 U501 ( .IN1(b[2]), .IN2(n445), .Q(n524) );
  AO22X1 U502 ( .IN1(n526), .IN2(n452), .IN3(n474), .IN4(n525), .Q(n172) );
  AO22X1 U503 ( .IN1(n527), .IN2(n452), .IN3(n474), .IN4(n526), .Q(n171) );
  AO22X1 U504 ( .IN1(n528), .IN2(n452), .IN3(n474), .IN4(n527), .Q(n170) );
  XOR2X1 U505 ( .IN1(n410), .IN2(n445), .Q(n527) );
  AO22X1 U506 ( .IN1(n529), .IN2(n452), .IN3(n474), .IN4(n528), .Q(n169) );
  XOR2X1 U507 ( .IN1(b[6]), .IN2(n445), .Q(n528) );
  AO22X1 U508 ( .IN1(n530), .IN2(n452), .IN3(n474), .IN4(n529), .Q(n168) );
  XOR2X1 U509 ( .IN1(b[7]), .IN2(n445), .Q(n529) );
  AO22X1 U510 ( .IN1(n531), .IN2(n452), .IN3(n474), .IN4(n530), .Q(n167) );
  XOR2X1 U511 ( .IN1(b[8]), .IN2(n445), .Q(n530) );
  AO22X1 U512 ( .IN1(n475), .IN2(n452), .IN3(n474), .IN4(n531), .Q(n166) );
  XOR2X1 U513 ( .IN1(b[9]), .IN2(n445), .Q(n531) );
  XOR2X1 U514 ( .IN1(b[10]), .IN2(n445), .Q(n475) );
  OAI21X1 U515 ( .IN1(n452), .IN2(n474), .IN3(n473), .QN(n165) );
  NOR2X0 U516 ( .IN1(n532), .IN2(n435), .QN(n164) );
  AO22X1 U517 ( .IN1(n533), .IN2(n450), .IN3(n477), .IN4(n534), .Q(n163) );
  XOR2X1 U518 ( .IN1(n434), .IN2(n447), .Q(n534) );
  AO22X1 U519 ( .IN1(n535), .IN2(n450), .IN3(n477), .IN4(n533), .Q(n162) );
  AO22X1 U520 ( .IN1(n536), .IN2(n450), .IN3(n477), .IN4(n535), .Q(n161) );
  XOR2X1 U521 ( .IN1(b[2]), .IN2(n447), .Q(n535) );
  AO22X1 U522 ( .IN1(n537), .IN2(n450), .IN3(n477), .IN4(n536), .Q(n160) );
  AO22X1 U523 ( .IN1(n538), .IN2(n450), .IN3(n477), .IN4(n537), .Q(n159) );
  AO22X1 U524 ( .IN1(n539), .IN2(n450), .IN3(n477), .IN4(n538), .Q(n158) );
  XOR2X1 U525 ( .IN1(n410), .IN2(n447), .Q(n538) );
  AO22X1 U526 ( .IN1(n540), .IN2(n450), .IN3(n477), .IN4(n539), .Q(n157) );
  XOR2X1 U527 ( .IN1(b[6]), .IN2(n447), .Q(n539) );
  AO22X1 U528 ( .IN1(n541), .IN2(n450), .IN3(n477), .IN4(n540), .Q(n156) );
  XOR2X1 U529 ( .IN1(b[7]), .IN2(n447), .Q(n540) );
  AO22X1 U530 ( .IN1(n542), .IN2(n450), .IN3(n477), .IN4(n541), .Q(n155) );
  XOR2X1 U531 ( .IN1(b[8]), .IN2(n447), .Q(n541) );
  AO22X1 U532 ( .IN1(n478), .IN2(n450), .IN3(n477), .IN4(n542), .Q(n154) );
  XOR2X1 U533 ( .IN1(b[9]), .IN2(n447), .Q(n542) );
  XOR2X1 U534 ( .IN1(b[10]), .IN2(n447), .Q(n478) );
  OAI21X1 U535 ( .IN1(n450), .IN2(n477), .IN3(n476), .QN(n153) );
  AO21X1 U536 ( .IN1(a[1]), .IN2(n436), .IN3(n464), .Q(n152) );
  AO22X1 U537 ( .IN1(n543), .IN2(n440), .IN3(n462), .IN4(n440), .Q(n151) );
  XOR2X1 U538 ( .IN1(n439), .IN2(a[2]), .Q(n544) );
  NOR2X0 U539 ( .IN1(n434), .IN2(n489), .QN(n543) );
  XNOR2X1 U540 ( .IN1(a[2]), .IN2(a[1]), .Q(n489) );
  AO22X1 U541 ( .IN1(n545), .IN2(n442), .IN3(n468), .IN4(n442), .Q(n150) );
  XOR2X1 U542 ( .IN1(n441), .IN2(a[4]), .Q(n546) );
  NOR2X0 U543 ( .IN1(n434), .IN2(n499), .QN(n545) );
  XNOR2X1 U544 ( .IN1(a[4]), .IN2(n439), .Q(n499) );
  AO22X1 U545 ( .IN1(n547), .IN2(n444), .IN3(n471), .IN4(n444), .Q(n149) );
  XOR2X1 U546 ( .IN1(n443), .IN2(a[6]), .Q(n548) );
  NOR2X0 U547 ( .IN1(n434), .IN2(n510), .QN(n547) );
  XNOR2X1 U548 ( .IN1(a[6]), .IN2(n441), .Q(n510) );
  AO22X1 U549 ( .IN1(n549), .IN2(n446), .IN3(n474), .IN4(n446), .Q(n148) );
  XOR2X1 U550 ( .IN1(n445), .IN2(a[8]), .Q(n550) );
  NOR2X0 U551 ( .IN1(n434), .IN2(n521), .QN(n549) );
  XNOR2X1 U552 ( .IN1(a[8]), .IN2(n443), .Q(n521) );
  AO22X1 U553 ( .IN1(n551), .IN2(n447), .IN3(n477), .IN4(n447), .Q(n147) );
  XOR2X1 U554 ( .IN1(n447), .IN2(a[10]), .Q(n552) );
  NOR2X0 U555 ( .IN1(n434), .IN2(n532), .QN(n551) );
  XNOR2X1 U556 ( .IN1(a[10]), .IN2(n445), .Q(n532) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_1 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;

  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_1_DW_mult_tc_0 mult_30 ( .a(in_a), .b(in_b), 
        .product(pre_out) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_0_DW_mult_tc_0 ( a, b, product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556;

  FADDX1 U4 ( .A(n25), .B(n153), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n453), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U22 ( .A(n132), .B(n133), .CI(n22), .CO(n21), .S(product[4]) );
  FADDX1 U23 ( .A(n134), .B(n151), .CI(n23), .CO(n22), .S(product[3]) );
  FADDX1 U24 ( .A(n223), .B(n212), .CI(n24), .CO(n23), .S(product[2]) );
  HADDX1 U25 ( .A0(n152), .B0(n224), .C1(n24), .SO(product[1]) );
  FADDX1 U27 ( .A(n154), .B(n165), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n455), .B(n155), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n166), .B(n177), .CI(n156), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n157), .B(n167), .CI(n457), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n168), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n158), .B(n189), .CI(n178), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n459), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n159), .B(n169), .CI(n179), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n170), .B(n73), .CI(n180), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n160), .B(n201), .CI(n190), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n461), .B(n181), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n191), .B(n171), .CI(n161), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n182), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n162), .B(n192), .CI(n172), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n173), .B(n193), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n147), .B(n183), .CI(n203), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n214), .B0(n163), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n184), .B(n174), .CI(n194), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n215), .B(n164), .CI(n204), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n205), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n148), .B(n185), .CI(n195), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n216), .B0(n175), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n119), .B(n116), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n186), .B(n196), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n217), .B(n176), .CI(n206), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n149), .B(n207), .CI(n197), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n218), .B0(n187), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n198), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n219), .B(n188), .CI(n208), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n150), .B(n199), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n220), .B0(n209), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n210), .B(n200), .CI(n221), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n222), .B0(n211), .C1(n133), .SO(n134) );
  FADDX1 U311 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  XOR3X1 U312 ( .IN1(n33), .IN2(n30), .IN3(n414), .Q(product[19]) );
  XOR2X2 U313 ( .IN1(n438), .IN2(n451), .Q(n538) );
  XOR2X2 U314 ( .IN1(n438), .IN2(n449), .Q(n527) );
  XOR2X2 U315 ( .IN1(n438), .IN2(n447), .Q(n516) );
  XOR2X2 U316 ( .IN1(n438), .IN2(n445), .Q(n505) );
  INVX0 U317 ( .INP(b[3]), .ZN(n408) );
  INVX0 U318 ( .INP(n408), .ZN(n409) );
  DELLN2X2 U319 ( .INP(n8), .Z(n410) );
  INVX0 U320 ( .INP(b[6]), .ZN(n411) );
  INVX0 U321 ( .INP(n411), .ZN(n412) );
  DELLN2X2 U322 ( .INP(n16), .Z(n413) );
  DELLN2X2 U323 ( .INP(n7), .Z(n414) );
  INVX0 U324 ( .INP(b[1]), .ZN(n415) );
  INVX0 U325 ( .INP(n415), .ZN(n416) );
  XOR2X2 U326 ( .IN1(b[9]), .IN2(n451), .Q(n546) );
  XOR2X2 U327 ( .IN1(b[9]), .IN2(n449), .Q(n535) );
  XOR2X2 U328 ( .IN1(b[9]), .IN2(n447), .Q(n524) );
  XOR2X2 U329 ( .IN1(b[9]), .IN2(n445), .Q(n513) );
  XOR2X2 U330 ( .IN1(b[9]), .IN2(n443), .Q(n467) );
  XOR2X2 U331 ( .IN1(b[9]), .IN2(a[1]), .Q(n491) );
  XOR2X2 U332 ( .IN1(n412), .IN2(n451), .Q(n543) );
  XOR2X2 U333 ( .IN1(n412), .IN2(n449), .Q(n532) );
  XOR2X2 U334 ( .IN1(n412), .IN2(n447), .Q(n521) );
  XOR2X2 U335 ( .IN1(n412), .IN2(n445), .Q(n510) );
  XOR2X2 U336 ( .IN1(n412), .IN2(n443), .Q(n500) );
  XOR2X2 U337 ( .IN1(n412), .IN2(a[1]), .Q(n488) );
  XOR2X2 U338 ( .IN1(b[8]), .IN2(n451), .Q(n545) );
  XOR2X2 U339 ( .IN1(b[8]), .IN2(n449), .Q(n534) );
  XOR2X2 U340 ( .IN1(b[8]), .IN2(n447), .Q(n523) );
  XOR2X2 U341 ( .IN1(b[8]), .IN2(n445), .Q(n512) );
  XOR2X2 U342 ( .IN1(b[8]), .IN2(n443), .Q(n502) );
  XOR2X2 U343 ( .IN1(b[8]), .IN2(a[1]), .Q(n490) );
  XOR2X2 U344 ( .IN1(b[4]), .IN2(n451), .Q(n541) );
  XOR2X2 U345 ( .IN1(b[4]), .IN2(n449), .Q(n530) );
  XOR2X2 U346 ( .IN1(b[4]), .IN2(n447), .Q(n519) );
  XOR2X2 U347 ( .IN1(b[4]), .IN2(n445), .Q(n508) );
  XOR2X2 U348 ( .IN1(b[4]), .IN2(n443), .Q(n498) );
  XOR2X2 U349 ( .IN1(b[4]), .IN2(a[1]), .Q(n486) );
  XOR2X2 U350 ( .IN1(n409), .IN2(n451), .Q(n540) );
  XOR2X2 U351 ( .IN1(n409), .IN2(n449), .Q(n529) );
  XOR2X2 U352 ( .IN1(n409), .IN2(n447), .Q(n518) );
  XOR2X2 U353 ( .IN1(n409), .IN2(n445), .Q(n507) );
  XOR2X2 U354 ( .IN1(n409), .IN2(n443), .Q(n497) );
  XOR2X2 U355 ( .IN1(n409), .IN2(a[1]), .Q(n485) );
  NAND2X1 U356 ( .IN1(n33), .IN2(n30), .QN(n417) );
  NAND2X0 U357 ( .IN1(n33), .IN2(n7), .QN(n418) );
  NAND2X0 U358 ( .IN1(n30), .IN2(n7), .QN(n419) );
  NAND3X0 U359 ( .IN1(n419), .IN2(n418), .IN3(n417), .QN(n6) );
  XOR2X1 U360 ( .IN1(n29), .IN2(n28), .Q(n420) );
  XOR2X1 U361 ( .IN1(n420), .IN2(n6), .Q(product[20]) );
  NAND2X1 U362 ( .IN1(n29), .IN2(n28), .QN(n421) );
  NAND2X0 U363 ( .IN1(n29), .IN2(n6), .QN(n422) );
  NAND2X0 U364 ( .IN1(n28), .IN2(n6), .QN(n423) );
  NAND3X0 U365 ( .IN1(n421), .IN2(n422), .IN3(n423), .QN(n5) );
  FADDX1 U366 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U367 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U368 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  XNOR2X1 U369 ( .IN1(n424), .IN2(n410), .Q(product[18]) );
  XNOR2X1 U370 ( .IN1(n37), .IN2(n34), .Q(n424) );
  XOR3X1 U371 ( .IN1(n43), .IN2(n38), .IN3(n9), .Q(product[17]) );
  XOR3X1 U372 ( .IN1(n104), .IN2(n111), .IN3(n17), .Q(product[9]) );
  XNOR2X1 U373 ( .IN1(n425), .IN2(n413), .Q(product[10]) );
  XNOR2X1 U374 ( .IN1(n96), .IN2(n103), .Q(n425) );
  INVX0 U375 ( .INP(n25), .ZN(n453) );
  FADDX1 U376 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  INVX0 U377 ( .INP(n3), .ZN(product[23]) );
  INVX0 U378 ( .INP(n55), .ZN(n459) );
  FADDX1 U379 ( .A(n124), .B(n127), .CI(n20), .CO(n19), .S(product[6]) );
  FADDX1 U380 ( .A(n128), .B(n131), .CI(n21), .CO(n20), .S(product[5]) );
  XOR2X1 U381 ( .IN1(b[2]), .IN2(a[1]), .Q(n484) );
  XOR2X1 U382 ( .IN1(n416), .IN2(a[1]), .Q(n483) );
  XOR2X1 U383 ( .IN1(n416), .IN2(n443), .Q(n494) );
  XOR2X1 U384 ( .IN1(n416), .IN2(n445), .Q(n504) );
  XOR2X1 U385 ( .IN1(n416), .IN2(n447), .Q(n515) );
  INVX0 U386 ( .INP(n73), .ZN(n461) );
  XOR2X1 U387 ( .IN1(n416), .IN2(n449), .Q(n526) );
  XOR2X1 U388 ( .IN1(n416), .IN2(n451), .Q(n537) );
  INVX0 U389 ( .INP(n31), .ZN(n455) );
  INVX0 U390 ( .INP(n41), .ZN(n457) );
  INVX0 U391 ( .INP(n493), .ZN(n462) );
  INVX0 U392 ( .INP(n503), .ZN(n460) );
  INVX0 U393 ( .INP(n514), .ZN(n458) );
  AND2X1 U394 ( .IN1(a[1]), .IN2(n442), .Q(n468) );
  INVX0 U395 ( .INP(n525), .ZN(n456) );
  INVX0 U396 ( .INP(n536), .ZN(n454) );
  NBUFFX2 U397 ( .INP(a[5]), .Z(n446) );
  NBUFFX2 U398 ( .INP(a[3]), .Z(n444) );
  AND2X1 U399 ( .IN1(n493), .IN2(n548), .Q(n466) );
  AND2X1 U400 ( .IN1(n514), .IN2(n552), .Q(n475) );
  AND2X1 U401 ( .IN1(n503), .IN2(n550), .Q(n472) );
  AND2X1 U402 ( .IN1(n525), .IN2(n554), .Q(n478) );
  AND2X1 U403 ( .IN1(n536), .IN2(n556), .Q(n481) );
  NBUFFX2 U404 ( .INP(a[7]), .Z(n448) );
  NBUFFX2 U405 ( .INP(a[9]), .Z(n450) );
  NAND2X0 U406 ( .IN1(n43), .IN2(n38), .QN(n426) );
  NAND2X0 U407 ( .IN1(n43), .IN2(n9), .QN(n427) );
  NAND2X0 U408 ( .IN1(n38), .IN2(n9), .QN(n428) );
  NAND3X0 U409 ( .IN1(n428), .IN2(n427), .IN3(n426), .QN(n8) );
  NAND2X0 U410 ( .IN1(n37), .IN2(n34), .QN(n429) );
  NAND2X0 U411 ( .IN1(n37), .IN2(n8), .QN(n430) );
  NAND2X0 U412 ( .IN1(n34), .IN2(n8), .QN(n431) );
  NAND3X0 U413 ( .IN1(n431), .IN2(n430), .IN3(n429), .QN(n7) );
  NAND2X0 U414 ( .IN1(n104), .IN2(n111), .QN(n432) );
  NAND2X0 U415 ( .IN1(n104), .IN2(n17), .QN(n433) );
  NAND2X0 U416 ( .IN1(n111), .IN2(n17), .QN(n434) );
  NAND3X0 U417 ( .IN1(n432), .IN2(n433), .IN3(n434), .QN(n16) );
  NAND2X0 U418 ( .IN1(n96), .IN2(n103), .QN(n435) );
  NAND2X0 U419 ( .IN1(n96), .IN2(n16), .QN(n436) );
  NAND2X0 U420 ( .IN1(n103), .IN2(n16), .QN(n437) );
  NAND3X0 U421 ( .IN1(n435), .IN2(n436), .IN3(n437), .QN(n15) );
  DELLN1X2 U422 ( .INP(a[11]), .Z(n451) );
  INVX0 U423 ( .INP(n440), .ZN(n438) );
  INVX0 U424 ( .INP(b[0]), .ZN(n439) );
  INVX0 U425 ( .INP(b[0]), .ZN(n440) );
  INVX0 U426 ( .INP(n442), .ZN(n441) );
  INVX0 U427 ( .INP(a[0]), .ZN(n442) );
  DELLN1X2 U428 ( .INP(a[3]), .Z(n443) );
  DELLN1X2 U429 ( .INP(a[5]), .Z(n445) );
  DELLN1X2 U430 ( .INP(a[7]), .Z(n447) );
  DELLN1X2 U431 ( .INP(a[9]), .Z(n449) );
  NOR2X0 U432 ( .IN1(n442), .IN2(n439), .QN(product[0]) );
  XNOR2X1 U433 ( .IN1(n463), .IN2(n464), .Q(n84) );
  NAND2X0 U434 ( .IN1(n464), .IN2(n463), .QN(n83) );
  AOI22X1 U435 ( .IN1(n465), .IN2(n462), .IN3(n466), .IN4(n467), .QN(n463) );
  OA21X1 U436 ( .IN1(n468), .IN2(n441), .IN3(n469), .Q(n464) );
  AO22X1 U437 ( .IN1(n470), .IN2(n462), .IN3(n466), .IN4(n465), .Q(n73) );
  XOR2X1 U438 ( .IN1(b[10]), .IN2(n443), .Q(n465) );
  AO22X1 U439 ( .IN1(n471), .IN2(n460), .IN3(n472), .IN4(n473), .Q(n55) );
  AO22X1 U440 ( .IN1(n474), .IN2(n458), .IN3(n475), .IN4(n476), .Q(n41) );
  AO22X1 U441 ( .IN1(n477), .IN2(n456), .IN3(n478), .IN4(n479), .Q(n31) );
  AO22X1 U442 ( .IN1(n480), .IN2(n454), .IN3(n481), .IN4(n482), .Q(n25) );
  AO22X1 U443 ( .IN1(n441), .IN2(n483), .IN3(n468), .IN4(n440), .Q(n224) );
  AO22X1 U444 ( .IN1(n441), .IN2(n484), .IN3(n468), .IN4(n483), .Q(n223) );
  AO22X1 U445 ( .IN1(n441), .IN2(n485), .IN3(n468), .IN4(n484), .Q(n222) );
  AO22X1 U446 ( .IN1(n441), .IN2(n486), .IN3(n468), .IN4(n485), .Q(n221) );
  AO22X1 U447 ( .IN1(n441), .IN2(n487), .IN3(n468), .IN4(n486), .Q(n220) );
  AO22X1 U448 ( .IN1(n441), .IN2(n488), .IN3(n468), .IN4(n487), .Q(n219) );
  XOR2X1 U449 ( .IN1(b[5]), .IN2(a[1]), .Q(n487) );
  AO22X1 U450 ( .IN1(n441), .IN2(n489), .IN3(n468), .IN4(n488), .Q(n218) );
  AO22X1 U451 ( .IN1(n441), .IN2(n490), .IN3(n468), .IN4(n489), .Q(n217) );
  XOR2X1 U452 ( .IN1(b[7]), .IN2(a[1]), .Q(n489) );
  AO22X1 U453 ( .IN1(n441), .IN2(n491), .IN3(n468), .IN4(n490), .Q(n216) );
  AO22X1 U454 ( .IN1(n441), .IN2(n492), .IN3(n468), .IN4(n491), .Q(n215) );
  AO22X1 U455 ( .IN1(n441), .IN2(n469), .IN3(n468), .IN4(n492), .Q(n214) );
  XOR2X1 U456 ( .IN1(b[10]), .IN2(a[1]), .Q(n492) );
  XOR2X1 U457 ( .IN1(b[11]), .IN2(a[1]), .Q(n469) );
  NOR2X0 U458 ( .IN1(n493), .IN2(n439), .QN(n212) );
  AO22X1 U459 ( .IN1(n494), .IN2(n462), .IN3(n466), .IN4(n495), .Q(n211) );
  XOR2X1 U460 ( .IN1(n438), .IN2(n443), .Q(n495) );
  AO22X1 U461 ( .IN1(n496), .IN2(n462), .IN3(n466), .IN4(n494), .Q(n210) );
  AO22X1 U462 ( .IN1(n497), .IN2(n462), .IN3(n466), .IN4(n496), .Q(n209) );
  XOR2X1 U463 ( .IN1(b[2]), .IN2(n443), .Q(n496) );
  AO22X1 U464 ( .IN1(n498), .IN2(n462), .IN3(n466), .IN4(n497), .Q(n208) );
  AO22X1 U465 ( .IN1(n499), .IN2(n462), .IN3(n466), .IN4(n498), .Q(n207) );
  AO22X1 U466 ( .IN1(n500), .IN2(n462), .IN3(n466), .IN4(n499), .Q(n206) );
  XOR2X1 U467 ( .IN1(b[5]), .IN2(n443), .Q(n499) );
  AO22X1 U468 ( .IN1(n501), .IN2(n462), .IN3(n466), .IN4(n500), .Q(n205) );
  AO22X1 U469 ( .IN1(n502), .IN2(n462), .IN3(n466), .IN4(n501), .Q(n204) );
  XOR2X1 U470 ( .IN1(b[7]), .IN2(n443), .Q(n501) );
  AO22X1 U471 ( .IN1(n467), .IN2(n462), .IN3(n466), .IN4(n502), .Q(n203) );
  OAI21X1 U472 ( .IN1(n462), .IN2(n466), .IN3(n470), .QN(n201) );
  XOR2X1 U473 ( .IN1(b[11]), .IN2(n443), .Q(n470) );
  NOR2X0 U474 ( .IN1(n503), .IN2(n439), .QN(n200) );
  AO22X1 U475 ( .IN1(n504), .IN2(n460), .IN3(n472), .IN4(n505), .Q(n199) );
  AO22X1 U476 ( .IN1(n506), .IN2(n460), .IN3(n472), .IN4(n504), .Q(n198) );
  AO22X1 U477 ( .IN1(n507), .IN2(n460), .IN3(n472), .IN4(n506), .Q(n197) );
  XOR2X1 U478 ( .IN1(b[2]), .IN2(n445), .Q(n506) );
  AO22X1 U479 ( .IN1(n508), .IN2(n460), .IN3(n472), .IN4(n507), .Q(n196) );
  AO22X1 U480 ( .IN1(n509), .IN2(n460), .IN3(n472), .IN4(n508), .Q(n195) );
  AO22X1 U481 ( .IN1(n510), .IN2(n460), .IN3(n472), .IN4(n509), .Q(n194) );
  XOR2X1 U482 ( .IN1(b[5]), .IN2(n445), .Q(n509) );
  AO22X1 U483 ( .IN1(n511), .IN2(n460), .IN3(n472), .IN4(n510), .Q(n193) );
  AO22X1 U484 ( .IN1(n512), .IN2(n460), .IN3(n472), .IN4(n511), .Q(n192) );
  XOR2X1 U485 ( .IN1(b[7]), .IN2(n445), .Q(n511) );
  AO22X1 U486 ( .IN1(n513), .IN2(n460), .IN3(n472), .IN4(n512), .Q(n191) );
  AO22X1 U487 ( .IN1(n473), .IN2(n460), .IN3(n472), .IN4(n513), .Q(n190) );
  XOR2X1 U488 ( .IN1(b[10]), .IN2(n445), .Q(n473) );
  OAI21X1 U489 ( .IN1(n460), .IN2(n472), .IN3(n471), .QN(n189) );
  XOR2X1 U490 ( .IN1(b[11]), .IN2(n445), .Q(n471) );
  NOR2X0 U491 ( .IN1(n514), .IN2(n439), .QN(n188) );
  AO22X1 U492 ( .IN1(n515), .IN2(n458), .IN3(n475), .IN4(n516), .Q(n187) );
  AO22X1 U493 ( .IN1(n517), .IN2(n458), .IN3(n475), .IN4(n515), .Q(n186) );
  AO22X1 U494 ( .IN1(n518), .IN2(n458), .IN3(n475), .IN4(n517), .Q(n185) );
  XOR2X1 U495 ( .IN1(b[2]), .IN2(n447), .Q(n517) );
  AO22X1 U496 ( .IN1(n519), .IN2(n458), .IN3(n475), .IN4(n518), .Q(n184) );
  AO22X1 U497 ( .IN1(n520), .IN2(n458), .IN3(n475), .IN4(n519), .Q(n183) );
  AO22X1 U498 ( .IN1(n521), .IN2(n458), .IN3(n475), .IN4(n520), .Q(n182) );
  XOR2X1 U499 ( .IN1(b[5]), .IN2(n447), .Q(n520) );
  AO22X1 U500 ( .IN1(n522), .IN2(n458), .IN3(n475), .IN4(n521), .Q(n181) );
  AO22X1 U501 ( .IN1(n523), .IN2(n458), .IN3(n475), .IN4(n522), .Q(n180) );
  XOR2X1 U502 ( .IN1(b[7]), .IN2(n447), .Q(n522) );
  AO22X1 U503 ( .IN1(n524), .IN2(n458), .IN3(n475), .IN4(n523), .Q(n179) );
  AO22X1 U504 ( .IN1(n476), .IN2(n458), .IN3(n475), .IN4(n524), .Q(n178) );
  XOR2X1 U505 ( .IN1(b[10]), .IN2(n447), .Q(n476) );
  OAI21X1 U506 ( .IN1(n458), .IN2(n475), .IN3(n474), .QN(n177) );
  XOR2X1 U507 ( .IN1(b[11]), .IN2(n447), .Q(n474) );
  NOR2X0 U508 ( .IN1(n525), .IN2(n439), .QN(n176) );
  AO22X1 U509 ( .IN1(n526), .IN2(n456), .IN3(n478), .IN4(n527), .Q(n175) );
  AO22X1 U510 ( .IN1(n528), .IN2(n456), .IN3(n478), .IN4(n526), .Q(n174) );
  AO22X1 U511 ( .IN1(n529), .IN2(n456), .IN3(n478), .IN4(n528), .Q(n173) );
  XOR2X1 U512 ( .IN1(b[2]), .IN2(n449), .Q(n528) );
  AO22X1 U513 ( .IN1(n530), .IN2(n456), .IN3(n478), .IN4(n529), .Q(n172) );
  AO22X1 U514 ( .IN1(n531), .IN2(n456), .IN3(n478), .IN4(n530), .Q(n171) );
  AO22X1 U515 ( .IN1(n532), .IN2(n456), .IN3(n478), .IN4(n531), .Q(n170) );
  XOR2X1 U516 ( .IN1(b[5]), .IN2(n449), .Q(n531) );
  AO22X1 U517 ( .IN1(n533), .IN2(n456), .IN3(n478), .IN4(n532), .Q(n169) );
  AO22X1 U518 ( .IN1(n534), .IN2(n456), .IN3(n478), .IN4(n533), .Q(n168) );
  XOR2X1 U519 ( .IN1(b[7]), .IN2(n449), .Q(n533) );
  AO22X1 U520 ( .IN1(n535), .IN2(n456), .IN3(n478), .IN4(n534), .Q(n167) );
  AO22X1 U521 ( .IN1(n479), .IN2(n456), .IN3(n478), .IN4(n535), .Q(n166) );
  XOR2X1 U522 ( .IN1(b[10]), .IN2(n449), .Q(n479) );
  OAI21X1 U523 ( .IN1(n456), .IN2(n478), .IN3(n477), .QN(n165) );
  XOR2X1 U524 ( .IN1(b[11]), .IN2(n449), .Q(n477) );
  NOR2X0 U525 ( .IN1(n536), .IN2(n439), .QN(n164) );
  AO22X1 U526 ( .IN1(n537), .IN2(n454), .IN3(n481), .IN4(n538), .Q(n163) );
  AO22X1 U527 ( .IN1(n539), .IN2(n454), .IN3(n481), .IN4(n537), .Q(n162) );
  AO22X1 U528 ( .IN1(n540), .IN2(n454), .IN3(n481), .IN4(n539), .Q(n161) );
  XOR2X1 U529 ( .IN1(b[2]), .IN2(n451), .Q(n539) );
  AO22X1 U530 ( .IN1(n541), .IN2(n454), .IN3(n481), .IN4(n540), .Q(n160) );
  AO22X1 U531 ( .IN1(n542), .IN2(n454), .IN3(n481), .IN4(n541), .Q(n159) );
  AO22X1 U532 ( .IN1(n543), .IN2(n454), .IN3(n481), .IN4(n542), .Q(n158) );
  XOR2X1 U533 ( .IN1(b[5]), .IN2(n451), .Q(n542) );
  AO22X1 U534 ( .IN1(n544), .IN2(n454), .IN3(n481), .IN4(n543), .Q(n157) );
  AO22X1 U535 ( .IN1(n545), .IN2(n454), .IN3(n481), .IN4(n544), .Q(n156) );
  XOR2X1 U536 ( .IN1(b[7]), .IN2(n451), .Q(n544) );
  AO22X1 U537 ( .IN1(n546), .IN2(n454), .IN3(n481), .IN4(n545), .Q(n155) );
  AO22X1 U538 ( .IN1(n482), .IN2(n454), .IN3(n481), .IN4(n546), .Q(n154) );
  XOR2X1 U539 ( .IN1(b[10]), .IN2(n451), .Q(n482) );
  OAI21X1 U540 ( .IN1(n454), .IN2(n481), .IN3(n480), .QN(n153) );
  XOR2X1 U541 ( .IN1(b[11]), .IN2(n451), .Q(n480) );
  AO21X1 U542 ( .IN1(a[1]), .IN2(n440), .IN3(n468), .Q(n152) );
  AO22X1 U543 ( .IN1(n547), .IN2(n444), .IN3(n466), .IN4(n444), .Q(n151) );
  XOR2X1 U544 ( .IN1(n443), .IN2(a[2]), .Q(n548) );
  NOR2X0 U545 ( .IN1(n438), .IN2(n493), .QN(n547) );
  XNOR2X1 U546 ( .IN1(a[2]), .IN2(a[1]), .Q(n493) );
  AO22X1 U547 ( .IN1(n549), .IN2(n446), .IN3(n472), .IN4(n446), .Q(n150) );
  XOR2X1 U548 ( .IN1(n445), .IN2(a[4]), .Q(n550) );
  NOR2X0 U549 ( .IN1(n438), .IN2(n503), .QN(n549) );
  XNOR2X1 U550 ( .IN1(a[4]), .IN2(n443), .Q(n503) );
  AO22X1 U551 ( .IN1(n551), .IN2(n448), .IN3(n475), .IN4(n448), .Q(n149) );
  XOR2X1 U552 ( .IN1(n447), .IN2(a[6]), .Q(n552) );
  NOR2X0 U553 ( .IN1(n438), .IN2(n514), .QN(n551) );
  XNOR2X1 U554 ( .IN1(a[6]), .IN2(n445), .Q(n514) );
  AO22X1 U555 ( .IN1(n553), .IN2(n450), .IN3(n478), .IN4(n450), .Q(n148) );
  XOR2X1 U556 ( .IN1(n449), .IN2(a[8]), .Q(n554) );
  NOR2X0 U557 ( .IN1(n438), .IN2(n525), .QN(n553) );
  XNOR2X1 U558 ( .IN1(a[8]), .IN2(n447), .Q(n525) );
  AO22X1 U559 ( .IN1(n555), .IN2(n451), .IN3(n481), .IN4(n451), .Q(n147) );
  XOR2X1 U560 ( .IN1(n451), .IN2(a[10]), .Q(n556) );
  NOR2X0 U561 ( .IN1(n438), .IN2(n536), .QN(n555) );
  XNOR2X1 U562 ( .IN1(a[10]), .IN2(n449), .Q(n536) );
endmodule


module mult_pipe_WORD_WIDTH12_INT_BITS4_0 ( in_a, in_b, clk, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [23:0] \output ;
  input clk;
  wire   n1, n2, n3;
  wire   [23:0] pre_out;

  DFFX1 \out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(\output [23]) );
  DFFX1 \out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(\output [22]) );
  DFFX1 \out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(\output [21]) );
  DFFX1 \out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(\output [20]) );
  DFFX1 \out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(\output [19]) );
  DFFX1 \out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(\output [18]) );
  DFFX1 \out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(\output [17]) );
  DFFX1 \out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(\output [16]) );
  DFFX1 \out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(\output [15]) );
  DFFX1 \out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(\output [14]) );
  DFFX1 \out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(\output [13]) );
  DFFX1 \out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(\output [12]) );
  DFFX1 \out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(\output [11]) );
  DFFX1 \out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(\output [10]) );
  DFFX1 \out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(\output [9]) );
  DFFX1 \out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(\output [8]) );
  DFFX1 \out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(\output [7]) );
  DFFX1 \out_reg_reg[6]  ( .D(pre_out[6]), .CLK(clk), .Q(\output [6]) );
  DFFX1 \out_reg_reg[5]  ( .D(pre_out[5]), .CLK(clk), .Q(\output [5]) );
  DFFX1 \out_reg_reg[4]  ( .D(pre_out[4]), .CLK(clk), .Q(\output [4]) );
  DFFX1 \out_reg_reg[3]  ( .D(pre_out[3]), .CLK(clk), .Q(\output [3]) );
  DFFX1 \out_reg_reg[2]  ( .D(pre_out[2]), .CLK(clk), .Q(\output [2]) );
  DFFX1 \out_reg_reg[1]  ( .D(pre_out[1]), .CLK(clk), .Q(\output [1]) );
  DFFX1 \out_reg_reg[0]  ( .D(pre_out[0]), .CLK(clk), .Q(\output [0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_0_DW_mult_tc_0 mult_30 ( .a(in_a), .b({
        in_b[11:6], n3, in_b[4:3], n2, in_b[1:0]}), .product(pre_out) );
  INVX0 U3 ( .INP(in_b[2]), .ZN(n1) );
  INVX0 U4 ( .INP(n1), .ZN(n2) );
  NBUFFX2 U5 ( .INP(in_b[5]), .Z(n3) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_0_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  wire   [24:0] carry;

  FADDX1 U2_22 ( .A(A[22]), .B(n7), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n8), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n9), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n10), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n11), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n12), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n13), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n14), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n16), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n17), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n18), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n19), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n20), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n21), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8])
         );
  FADDX1 U2_7 ( .A(A[7]), .B(n22), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  XNOR3X1 U1 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(DIFF[23]) );
  INVX0 U2 ( .INP(B[21]), .ZN(n8) );
  INVX0 U3 ( .INP(B[20]), .ZN(n9) );
  INVX0 U4 ( .INP(B[22]), .ZN(n7) );
  INVX0 U5 ( .INP(B[19]), .ZN(n10) );
  INVX0 U6 ( .INP(B[18]), .ZN(n11) );
  INVX0 U7 ( .INP(B[17]), .ZN(n12) );
  INVX0 U8 ( .INP(B[16]), .ZN(n13) );
  INVX0 U9 ( .INP(B[15]), .ZN(n14) );
  INVX0 U10 ( .INP(B[14]), .ZN(n15) );
  INVX0 U11 ( .INP(B[13]), .ZN(n16) );
  INVX0 U12 ( .INP(B[12]), .ZN(n17) );
  INVX0 U13 ( .INP(B[11]), .ZN(n18) );
  INVX0 U14 ( .INP(B[10]), .ZN(n19) );
  INVX0 U15 ( .INP(B[9]), .ZN(n20) );
  INVX0 U16 ( .INP(B[8]), .ZN(n21) );
  INVX0 U17 ( .INP(B[7]), .ZN(n22) );
  INVX0 U18 ( .INP(A[3]), .ZN(n4) );
  INVX0 U19 ( .INP(A[1]), .ZN(n6) );
  INVX0 U20 ( .INP(A[5]), .ZN(n2) );
  INVX0 U21 ( .INP(A[2]), .ZN(n5) );
  INVX0 U22 ( .INP(B[0]), .ZN(n23) );
  INVX0 U23 ( .INP(A[4]), .ZN(n3) );
  INVX0 U24 ( .INP(A[6]), .ZN(n1) );
  OAI22X1 U25 ( .IN1(n24), .IN2(n1), .IN3(B[6]), .IN4(n25), .QN(carry[7]) );
  AND2X1 U26 ( .IN1(n1), .IN2(n24), .Q(n25) );
  OA22X1 U27 ( .IN1(n26), .IN2(n2), .IN3(B[5]), .IN4(n27), .Q(n24) );
  AND2X1 U28 ( .IN1(n2), .IN2(n26), .Q(n27) );
  OA22X1 U29 ( .IN1(n28), .IN2(n3), .IN3(B[4]), .IN4(n29), .Q(n26) );
  AND2X1 U30 ( .IN1(n3), .IN2(n28), .Q(n29) );
  OA22X1 U31 ( .IN1(n30), .IN2(n4), .IN3(B[3]), .IN4(n31), .Q(n28) );
  AND2X1 U32 ( .IN1(n4), .IN2(n30), .Q(n31) );
  OA22X1 U33 ( .IN1(n32), .IN2(n5), .IN3(B[2]), .IN4(n33), .Q(n30) );
  AND2X1 U34 ( .IN1(n5), .IN2(n32), .Q(n33) );
  OA22X1 U35 ( .IN1(n34), .IN2(n6), .IN3(B[1]), .IN4(n35), .Q(n32) );
  AND2X1 U36 ( .IN1(n6), .IN2(n34), .Q(n35) );
  NOR2X0 U37 ( .IN1(n23), .IN2(A[0]), .QN(n34) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_0 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_0_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(\output ) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_0_DW01_add_0 ( A, B, CI, SUM, 
        CO );
  input [23:0] A;
  input [23:0] B;
  output [23:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [23:1] carry;

  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  XOR3X1 U1_23 ( .IN1(A[23]), .IN2(B[23]), .IN3(carry[23]), .Q(SUM[23]) );
  AO22X1 U1 ( .IN1(A[6]), .IN2(n1), .IN3(B[6]), .IN4(n2), .Q(carry[7]) );
  OR2X1 U2 ( .IN1(n1), .IN2(A[6]), .Q(n2) );
  AO22X1 U3 ( .IN1(A[5]), .IN2(n3), .IN3(B[5]), .IN4(n4), .Q(n1) );
  OR2X1 U4 ( .IN1(n3), .IN2(A[5]), .Q(n4) );
  AO22X1 U5 ( .IN1(A[4]), .IN2(n5), .IN3(B[4]), .IN4(n6), .Q(n3) );
  OR2X1 U6 ( .IN1(n5), .IN2(A[4]), .Q(n6) );
  AO22X1 U7 ( .IN1(A[3]), .IN2(n7), .IN3(B[3]), .IN4(n8), .Q(n5) );
  OR2X1 U8 ( .IN1(n7), .IN2(A[3]), .Q(n8) );
  AO22X1 U9 ( .IN1(A[2]), .IN2(n9), .IN3(B[2]), .IN4(n10), .Q(n7) );
  OR2X1 U10 ( .IN1(n9), .IN2(A[2]), .Q(n10) );
  AO22X1 U11 ( .IN1(B[1]), .IN2(A[1]), .IN3(n11), .IN4(B[0]), .Q(n9) );
  OA21X1 U12 ( .IN1(A[1]), .IN2(B[1]), .IN3(A[0]), .Q(n11) );
endmodule


module add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_0 ( a, b, \output  );
  input [23:0] a;
  input [23:0] b;
  output [23:0] \output ;


  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_0_DW01_add_0 add_37 ( .A(a), .B(b), 
        .CI(1'b0), .SUM(\output ) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_DW01_inc_1 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0 ( a_r, a_i, b_r, b_i, out_r, 
        out_i, clk );
  input [11:0] a_r;
  input [11:0] a_i;
  input [11:0] b_r;
  input [11:0] b_i;
  output [11:0] out_r;
  output [11:0] out_i;
  input clk;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47;
  wire   [23:0] mult1_out;
  wire   [23:0] mult2_out;
  wire   [23:0] mult3_out;
  wire   [23:0] mult4_out;
  wire   [23:7] pre_out_r;
  wire   [23:7] pre_out_i;
  wire   [11:0] rnd_out_r;
  wire   [11:0] rnd_out_i;
  wire   [11:0] pos_out_r;
  wire   [11:0] pos_out_i;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFFX1 \out_r_reg_reg[11]  ( .D(pos_out_r[11]), .CLK(clk), .Q(out_r[11]) );
  DFFX1 \out_r_reg_reg[10]  ( .D(pos_out_r[10]), .CLK(clk), .Q(out_r[10]) );
  DFFX1 \out_r_reg_reg[9]  ( .D(pos_out_r[9]), .CLK(clk), .Q(out_r[9]) );
  DFFX1 \out_r_reg_reg[8]  ( .D(pos_out_r[8]), .CLK(clk), .Q(out_r[8]) );
  DFFX1 \out_r_reg_reg[7]  ( .D(pos_out_r[7]), .CLK(clk), .Q(out_r[7]) );
  DFFX1 \out_r_reg_reg[6]  ( .D(pos_out_r[6]), .CLK(clk), .Q(out_r[6]) );
  DFFX1 \out_r_reg_reg[5]  ( .D(pos_out_r[5]), .CLK(clk), .Q(out_r[5]) );
  DFFX1 \out_r_reg_reg[4]  ( .D(pos_out_r[4]), .CLK(clk), .Q(out_r[4]) );
  DFFX1 \out_r_reg_reg[3]  ( .D(pos_out_r[3]), .CLK(clk), .Q(out_r[3]) );
  DFFX1 \out_r_reg_reg[2]  ( .D(pos_out_r[2]), .CLK(clk), .Q(out_r[2]) );
  DFFX1 \out_r_reg_reg[1]  ( .D(pos_out_r[1]), .CLK(clk), .Q(out_r[1]) );
  DFFX1 \out_r_reg_reg[0]  ( .D(pos_out_r[0]), .CLK(clk), .Q(out_r[0]) );
  DFFX1 \out_i_reg_reg[11]  ( .D(pos_out_i[11]), .CLK(clk), .Q(out_i[11]) );
  DFFX1 \out_i_reg_reg[10]  ( .D(pos_out_i[10]), .CLK(clk), .Q(out_i[10]) );
  DFFX1 \out_i_reg_reg[9]  ( .D(pos_out_i[9]), .CLK(clk), .Q(out_i[9]) );
  DFFX1 \out_i_reg_reg[8]  ( .D(pos_out_i[8]), .CLK(clk), .Q(out_i[8]) );
  DFFX1 \out_i_reg_reg[7]  ( .D(pos_out_i[7]), .CLK(clk), .Q(out_i[7]) );
  DFFX1 \out_i_reg_reg[6]  ( .D(pos_out_i[6]), .CLK(clk), .Q(out_i[6]) );
  DFFX1 \out_i_reg_reg[5]  ( .D(pos_out_i[5]), .CLK(clk), .Q(out_i[5]) );
  DFFX1 \out_i_reg_reg[4]  ( .D(pos_out_i[4]), .CLK(clk), .Q(out_i[4]) );
  DFFX1 \out_i_reg_reg[3]  ( .D(pos_out_i[3]), .CLK(clk), .Q(out_i[3]) );
  DFFX1 \out_i_reg_reg[2]  ( .D(pos_out_i[2]), .CLK(clk), .Q(out_i[2]) );
  DFFX1 \out_i_reg_reg[1]  ( .D(pos_out_i[1]), .CLK(clk), .Q(out_i[1]) );
  DFFX1 \out_i_reg_reg[0]  ( .D(pos_out_i[0]), .CLK(clk), .Q(out_i[0]) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_3 mult1 ( .in_a({a_r[11:2], n17, a_r[0]}), 
        .in_b({b_r[11], n8, b_r[9:8], n6, b_r[6:5], n5, b_r[3:0]}), .clk(clk), 
        .\output (mult1_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_2 mult2 ( .in_a({a_i[11:2], n16, a_i[0]}), 
        .in_b({b_i[11:10], n14, b_i[8:7], n15, b_i[5:3], n13, b_i[1], n3}), 
        .clk(clk), .\output (mult2_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_1 mult3 ( .in_a({a_r[11:2], n17, a_r[0]}), 
        .in_b({b_i[11:10], n14, b_i[8:7], n15, b_i[5:3], n13, b_i[1], n2}), 
        .clk(clk), .\output (mult3_out) );
  mult_pipe_WORD_WIDTH12_INT_BITS4_0 mult4 ( .in_a({a_i[11:2], n16, a_i[0]}), 
        .in_b({b_r[11], n8, b_r[9:8], n6, b_r[6:5], n5, b_r[3:0]}), .clk(clk), 
        .\output (mult4_out) );
  add_sub_WORD_WIDTH24_OPERATION0_USE_SAT0_0 sub ( .a(mult1_out), .b(mult2_out), .\output ({pre_out_r, SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6}) );
  add_sub_WORD_WIDTH24_OPERATION1_USE_SAT0_0 add ( .a(mult3_out), .b(mult4_out), .\output ({pre_out_i, SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_DW01_inc_0 add_154_round ( .A(
        pre_out_i[19:7]), .SUM({rnd_out_i, SYNOPSYS_UNCONNECTED__14}) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0_DW01_inc_1 add_140_round ( .A(
        pre_out_r[19:7]), .SUM({rnd_out_r, SYNOPSYS_UNCONNECTED__15}) );
  DELLN2X2 U3 ( .INP(b_i[2]), .Z(n13) );
  DELLN2X2 U4 ( .INP(b_i[6]), .Z(n15) );
  INVX0 U5 ( .INP(n3), .ZN(n1) );
  INVX0 U6 ( .INP(n1), .ZN(n2) );
  DELLN2X2 U7 ( .INP(b_i[0]), .Z(n3) );
  INVX0 U8 ( .INP(b_r[4]), .ZN(n4) );
  INVX1 U9 ( .INP(n4), .ZN(n5) );
  DELLN2X2 U10 ( .INP(b_r[7]), .Z(n6) );
  INVX0 U11 ( .INP(b_r[10]), .ZN(n7) );
  INVX0 U12 ( .INP(n7), .ZN(n8) );
  INVX0 U13 ( .INP(pre_out_r[23]), .ZN(n40) );
  INVX0 U14 ( .INP(pre_out_i[23]), .ZN(n25) );
  INVX0 U15 ( .INP(n41), .ZN(n43) );
  INVX0 U16 ( .INP(n26), .ZN(n28) );
  AND2X1 U17 ( .IN1(n27), .IN2(n29), .Q(n9) );
  AND2X1 U18 ( .IN1(n42), .IN2(n44), .Q(n10) );
  AND2X1 U19 ( .IN1(n28), .IN2(n29), .Q(n11) );
  AND2X1 U20 ( .IN1(n43), .IN2(n44), .Q(n12) );
  NOR2X0 U21 ( .IN1(pre_out_r[21]), .IN2(pre_out_r[22]), .QN(n33) );
  NOR2X0 U22 ( .IN1(pre_out_i[21]), .IN2(pre_out_i[22]), .QN(n18) );
  NAND2X0 U23 ( .IN1(n34), .IN2(n33), .QN(n36) );
  NOR2X0 U24 ( .IN1(pre_out_r[19]), .IN2(pre_out_r[20]), .QN(n34) );
  NAND2X0 U25 ( .IN1(n19), .IN2(n18), .QN(n21) );
  NOR2X0 U26 ( .IN1(pre_out_i[19]), .IN2(pre_out_i[20]), .QN(n19) );
  INVX0 U27 ( .INP(n31), .ZN(n24) );
  INVX0 U28 ( .INP(n29), .ZN(n30) );
  INVX0 U29 ( .INP(n44), .ZN(n45) );
  INVX0 U30 ( .INP(n46), .ZN(n39) );
  DELLN1X2 U31 ( .INP(b_i[9]), .Z(n14) );
  XNOR2X1 U32 ( .IN1(mult3_out[23]), .IN2(mult4_out[23]), .Q(n23) );
  NAND2X0 U33 ( .IN1(n38), .IN2(n37), .QN(n46) );
  DELLN1X2 U34 ( .INP(a_i[1]), .Z(n16) );
  DELLN1X2 U35 ( .INP(a_r[1]), .Z(n17) );
  NAND4X0 U36 ( .IN1(pre_out_i[22]), .IN2(pre_out_i[21]), .IN3(pre_out_i[20]), 
        .IN4(pre_out_i[19]), .QN(n20) );
  MUX21X1 U37 ( .IN1(n21), .IN2(n20), .S(pre_out_i[23]), .Q(n26) );
  XOR2X1 U38 ( .IN1(pre_out_i[23]), .IN2(mult3_out[23]), .Q(n22) );
  NAND2X1 U39 ( .IN1(n23), .IN2(n22), .QN(n31) );
  NAND2X1 U40 ( .IN1(mult3_out[23]), .IN2(n24), .QN(n29) );
  AO21X1 U41 ( .IN1(n26), .IN2(n25), .IN3(n24), .Q(n27) );
  AO21X1 U42 ( .IN1(rnd_out_i[0]), .IN2(n11), .IN3(n9), .Q(pos_out_i[0]) );
  AO21X1 U43 ( .IN1(rnd_out_i[1]), .IN2(n11), .IN3(n9), .Q(pos_out_i[1]) );
  AO21X1 U44 ( .IN1(rnd_out_i[2]), .IN2(n11), .IN3(n9), .Q(pos_out_i[2]) );
  AO21X1 U45 ( .IN1(rnd_out_i[3]), .IN2(n11), .IN3(n9), .Q(pos_out_i[3]) );
  AO21X1 U46 ( .IN1(rnd_out_i[4]), .IN2(n11), .IN3(n9), .Q(pos_out_i[4]) );
  AO21X1 U47 ( .IN1(rnd_out_i[5]), .IN2(n11), .IN3(n9), .Q(pos_out_i[5]) );
  AO21X1 U48 ( .IN1(rnd_out_i[6]), .IN2(n11), .IN3(n9), .Q(pos_out_i[6]) );
  AO21X1 U49 ( .IN1(rnd_out_i[7]), .IN2(n11), .IN3(n9), .Q(pos_out_i[7]) );
  AO21X1 U50 ( .IN1(rnd_out_i[8]), .IN2(n11), .IN3(n9), .Q(pos_out_i[8]) );
  AO21X1 U51 ( .IN1(rnd_out_i[9]), .IN2(n11), .IN3(n9), .Q(pos_out_i[9]) );
  AO21X1 U52 ( .IN1(rnd_out_i[10]), .IN2(n11), .IN3(n9), .Q(pos_out_i[10]) );
  MUX21X1 U53 ( .IN1(pre_out_i[23]), .IN2(rnd_out_i[11]), .S(n28), .Q(n32) );
  AO21X1 U54 ( .IN1(n32), .IN2(n31), .IN3(n30), .Q(pos_out_i[11]) );
  NAND4X0 U55 ( .IN1(pre_out_r[22]), .IN2(pre_out_r[21]), .IN3(pre_out_r[20]), 
        .IN4(pre_out_r[19]), .QN(n35) );
  MUX21X1 U56 ( .IN1(n36), .IN2(n35), .S(pre_out_r[23]), .Q(n41) );
  XOR2X1 U57 ( .IN1(mult2_out[23]), .IN2(mult1_out[23]), .Q(n38) );
  XOR2X1 U58 ( .IN1(pre_out_r[23]), .IN2(mult1_out[23]), .Q(n37) );
  NAND2X1 U59 ( .IN1(mult1_out[23]), .IN2(n39), .QN(n44) );
  AO21X1 U60 ( .IN1(n41), .IN2(n40), .IN3(n39), .Q(n42) );
  AO21X1 U61 ( .IN1(rnd_out_r[0]), .IN2(n12), .IN3(n10), .Q(pos_out_r[0]) );
  AO21X1 U62 ( .IN1(rnd_out_r[1]), .IN2(n12), .IN3(n10), .Q(pos_out_r[1]) );
  AO21X1 U63 ( .IN1(rnd_out_r[2]), .IN2(n12), .IN3(n10), .Q(pos_out_r[2]) );
  AO21X1 U64 ( .IN1(rnd_out_r[3]), .IN2(n12), .IN3(n10), .Q(pos_out_r[3]) );
  AO21X1 U65 ( .IN1(rnd_out_r[4]), .IN2(n12), .IN3(n10), .Q(pos_out_r[4]) );
  AO21X1 U66 ( .IN1(rnd_out_r[5]), .IN2(n12), .IN3(n10), .Q(pos_out_r[5]) );
  AO21X1 U67 ( .IN1(rnd_out_r[6]), .IN2(n12), .IN3(n10), .Q(pos_out_r[6]) );
  AO21X1 U68 ( .IN1(rnd_out_r[7]), .IN2(n12), .IN3(n10), .Q(pos_out_r[7]) );
  AO21X1 U69 ( .IN1(rnd_out_r[8]), .IN2(n12), .IN3(n10), .Q(pos_out_r[8]) );
  AO21X1 U70 ( .IN1(rnd_out_r[9]), .IN2(n12), .IN3(n10), .Q(pos_out_r[9]) );
  AO21X1 U71 ( .IN1(rnd_out_r[10]), .IN2(n12), .IN3(n10), .Q(pos_out_r[10]) );
  MUX21X1 U72 ( .IN1(pre_out_r[23]), .IN2(rnd_out_r[11]), .S(n43), .Q(n47) );
  AO21X1 U73 ( .IN1(n47), .IN2(n46), .IN3(n45), .Q(pos_out_r[11]) );
endmodule


module vec_mult_N4_WORD_WIDTH12_INT_BITS4 ( .in_a_r({\in_a_r[0][11] , 
        \in_a_r[0][10] , \in_a_r[0][9] , \in_a_r[0][8] , \in_a_r[0][7] , 
        \in_a_r[0][6] , \in_a_r[0][5] , \in_a_r[0][4] , \in_a_r[0][3] , 
        \in_a_r[0][2] , \in_a_r[0][1] , \in_a_r[0][0] , \in_a_r[1][11] , 
        \in_a_r[1][10] , \in_a_r[1][9] , \in_a_r[1][8] , \in_a_r[1][7] , 
        \in_a_r[1][6] , \in_a_r[1][5] , \in_a_r[1][4] , \in_a_r[1][3] , 
        \in_a_r[1][2] , \in_a_r[1][1] , \in_a_r[1][0] , \in_a_r[2][11] , 
        \in_a_r[2][10] , \in_a_r[2][9] , \in_a_r[2][8] , \in_a_r[2][7] , 
        \in_a_r[2][6] , \in_a_r[2][5] , \in_a_r[2][4] , \in_a_r[2][3] , 
        \in_a_r[2][2] , \in_a_r[2][1] , \in_a_r[2][0] , \in_a_r[3][11] , 
        \in_a_r[3][10] , \in_a_r[3][9] , \in_a_r[3][8] , \in_a_r[3][7] , 
        \in_a_r[3][6] , \in_a_r[3][5] , \in_a_r[3][4] , \in_a_r[3][3] , 
        \in_a_r[3][2] , \in_a_r[3][1] , \in_a_r[3][0] }), .in_a_i({
        \in_a_i[0][11] , \in_a_i[0][10] , \in_a_i[0][9] , \in_a_i[0][8] , 
        \in_a_i[0][7] , \in_a_i[0][6] , \in_a_i[0][5] , \in_a_i[0][4] , 
        \in_a_i[0][3] , \in_a_i[0][2] , \in_a_i[0][1] , \in_a_i[0][0] , 
        \in_a_i[1][11] , \in_a_i[1][10] , \in_a_i[1][9] , \in_a_i[1][8] , 
        \in_a_i[1][7] , \in_a_i[1][6] , \in_a_i[1][5] , \in_a_i[1][4] , 
        \in_a_i[1][3] , \in_a_i[1][2] , \in_a_i[1][1] , \in_a_i[1][0] , 
        \in_a_i[2][11] , \in_a_i[2][10] , \in_a_i[2][9] , \in_a_i[2][8] , 
        \in_a_i[2][7] , \in_a_i[2][6] , \in_a_i[2][5] , \in_a_i[2][4] , 
        \in_a_i[2][3] , \in_a_i[2][2] , \in_a_i[2][1] , \in_a_i[2][0] , 
        \in_a_i[3][11] , \in_a_i[3][10] , \in_a_i[3][9] , \in_a_i[3][8] , 
        \in_a_i[3][7] , \in_a_i[3][6] , \in_a_i[3][5] , \in_a_i[3][4] , 
        \in_a_i[3][3] , \in_a_i[3][2] , \in_a_i[3][1] , \in_a_i[3][0] }), 
        in_b_r, in_b_i, .out_r({\out_r[0][11] , \out_r[0][10] , \out_r[0][9] , 
        \out_r[0][8] , \out_r[0][7] , \out_r[0][6] , \out_r[0][5] , 
        \out_r[0][4] , \out_r[0][3] , \out_r[0][2] , \out_r[0][1] , 
        \out_r[0][0] , \out_r[1][11] , \out_r[1][10] , \out_r[1][9] , 
        \out_r[1][8] , \out_r[1][7] , \out_r[1][6] , \out_r[1][5] , 
        \out_r[1][4] , \out_r[1][3] , \out_r[1][2] , \out_r[1][1] , 
        \out_r[1][0] , \out_r[2][11] , \out_r[2][10] , \out_r[2][9] , 
        \out_r[2][8] , \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , 
        \out_r[2][4] , \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , 
        \out_r[2][0] , \out_r[3][11] , \out_r[3][10] , \out_r[3][9] , 
        \out_r[3][8] , \out_r[3][7] , \out_r[3][6] , \out_r[3][5] , 
        \out_r[3][4] , \out_r[3][3] , \out_r[3][2] , \out_r[3][1] , 
        \out_r[3][0] }), .out_i({\out_i[0][11] , \out_i[0][10] , \out_i[0][9] , 
        \out_i[0][8] , \out_i[0][7] , \out_i[0][6] , \out_i[0][5] , 
        \out_i[0][4] , \out_i[0][3] , \out_i[0][2] , \out_i[0][1] , 
        \out_i[0][0] , \out_i[1][11] , \out_i[1][10] , \out_i[1][9] , 
        \out_i[1][8] , \out_i[1][7] , \out_i[1][6] , \out_i[1][5] , 
        \out_i[1][4] , \out_i[1][3] , \out_i[1][2] , \out_i[1][1] , 
        \out_i[1][0] , \out_i[2][11] , \out_i[2][10] , \out_i[2][9] , 
        \out_i[2][8] , \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , 
        \out_i[2][4] , \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , 
        \out_i[2][0] , \out_i[3][11] , \out_i[3][10] , \out_i[3][9] , 
        \out_i[3][8] , \out_i[3][7] , \out_i[3][6] , \out_i[3][5] , 
        \out_i[3][4] , \out_i[3][3] , \out_i[3][2] , \out_i[3][1] , 
        \out_i[3][0] }), clk );
  input [11:0] in_b_r;
  input [11:0] in_b_i;
  input \in_a_r[0][11] , \in_a_r[0][10] , \in_a_r[0][9] , \in_a_r[0][8] ,
         \in_a_r[0][7] , \in_a_r[0][6] , \in_a_r[0][5] , \in_a_r[0][4] ,
         \in_a_r[0][3] , \in_a_r[0][2] , \in_a_r[0][1] , \in_a_r[0][0] ,
         \in_a_r[1][11] , \in_a_r[1][10] , \in_a_r[1][9] , \in_a_r[1][8] ,
         \in_a_r[1][7] , \in_a_r[1][6] , \in_a_r[1][5] , \in_a_r[1][4] ,
         \in_a_r[1][3] , \in_a_r[1][2] , \in_a_r[1][1] , \in_a_r[1][0] ,
         \in_a_r[2][11] , \in_a_r[2][10] , \in_a_r[2][9] , \in_a_r[2][8] ,
         \in_a_r[2][7] , \in_a_r[2][6] , \in_a_r[2][5] , \in_a_r[2][4] ,
         \in_a_r[2][3] , \in_a_r[2][2] , \in_a_r[2][1] , \in_a_r[2][0] ,
         \in_a_r[3][11] , \in_a_r[3][10] , \in_a_r[3][9] , \in_a_r[3][8] ,
         \in_a_r[3][7] , \in_a_r[3][6] , \in_a_r[3][5] , \in_a_r[3][4] ,
         \in_a_r[3][3] , \in_a_r[3][2] , \in_a_r[3][1] , \in_a_r[3][0] ,
         \in_a_i[0][11] , \in_a_i[0][10] , \in_a_i[0][9] , \in_a_i[0][8] ,
         \in_a_i[0][7] , \in_a_i[0][6] , \in_a_i[0][5] , \in_a_i[0][4] ,
         \in_a_i[0][3] , \in_a_i[0][2] , \in_a_i[0][1] , \in_a_i[0][0] ,
         \in_a_i[1][11] , \in_a_i[1][10] , \in_a_i[1][9] , \in_a_i[1][8] ,
         \in_a_i[1][7] , \in_a_i[1][6] , \in_a_i[1][5] , \in_a_i[1][4] ,
         \in_a_i[1][3] , \in_a_i[1][2] , \in_a_i[1][1] , \in_a_i[1][0] ,
         \in_a_i[2][11] , \in_a_i[2][10] , \in_a_i[2][9] , \in_a_i[2][8] ,
         \in_a_i[2][7] , \in_a_i[2][6] , \in_a_i[2][5] , \in_a_i[2][4] ,
         \in_a_i[2][3] , \in_a_i[2][2] , \in_a_i[2][1] , \in_a_i[2][0] ,
         \in_a_i[3][11] , \in_a_i[3][10] , \in_a_i[3][9] , \in_a_i[3][8] ,
         \in_a_i[3][7] , \in_a_i[3][6] , \in_a_i[3][5] , \in_a_i[3][4] ,
         \in_a_i[3][3] , \in_a_i[3][2] , \in_a_i[3][1] , \in_a_i[3][0] , clk;
  output \out_r[0][11] , \out_r[0][10] , \out_r[0][9] , \out_r[0][8] ,
         \out_r[0][7] , \out_r[0][6] , \out_r[0][5] , \out_r[0][4] ,
         \out_r[0][3] , \out_r[0][2] , \out_r[0][1] , \out_r[0][0] ,
         \out_r[1][11] , \out_r[1][10] , \out_r[1][9] , \out_r[1][8] ,
         \out_r[1][7] , \out_r[1][6] , \out_r[1][5] , \out_r[1][4] ,
         \out_r[1][3] , \out_r[1][2] , \out_r[1][1] , \out_r[1][0] ,
         \out_r[2][11] , \out_r[2][10] , \out_r[2][9] , \out_r[2][8] ,
         \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , \out_r[2][4] ,
         \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , \out_r[2][0] ,
         \out_r[3][11] , \out_r[3][10] , \out_r[3][9] , \out_r[3][8] ,
         \out_r[3][7] , \out_r[3][6] , \out_r[3][5] , \out_r[3][4] ,
         \out_r[3][3] , \out_r[3][2] , \out_r[3][1] , \out_r[3][0] ,
         \out_i[0][11] , \out_i[0][10] , \out_i[0][9] , \out_i[0][8] ,
         \out_i[0][7] , \out_i[0][6] , \out_i[0][5] , \out_i[0][4] ,
         \out_i[0][3] , \out_i[0][2] , \out_i[0][1] , \out_i[0][0] ,
         \out_i[1][11] , \out_i[1][10] , \out_i[1][9] , \out_i[1][8] ,
         \out_i[1][7] , \out_i[1][6] , \out_i[1][5] , \out_i[1][4] ,
         \out_i[1][3] , \out_i[1][2] , \out_i[1][1] , \out_i[1][0] ,
         \out_i[2][11] , \out_i[2][10] , \out_i[2][9] , \out_i[2][8] ,
         \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , \out_i[2][4] ,
         \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , \out_i[2][0] ,
         \out_i[3][11] , \out_i[3][10] , \out_i[3][9] , \out_i[3][8] ,
         \out_i[3][7] , \out_i[3][6] , \out_i[3][5] , \out_i[3][4] ,
         \out_i[3][3] , \out_i[3][2] , \out_i[3][1] , \out_i[3][0] ;
  wire   \in_a_r_reg[0][11] , \in_a_r_reg[0][10] , \in_a_r_reg[0][9] ,
         \in_a_r_reg[0][8] , \in_a_r_reg[0][7] , \in_a_r_reg[0][6] ,
         \in_a_r_reg[0][5] , \in_a_r_reg[0][4] , \in_a_r_reg[0][3] ,
         \in_a_r_reg[0][2] , \in_a_r_reg[0][1] , \in_a_r_reg[0][0] ,
         \in_a_r_reg[1][11] , \in_a_r_reg[1][10] , \in_a_r_reg[1][9] ,
         \in_a_r_reg[1][8] , \in_a_r_reg[1][7] , \in_a_r_reg[1][6] ,
         \in_a_r_reg[1][5] , \in_a_r_reg[1][4] , \in_a_r_reg[1][3] ,
         \in_a_r_reg[1][2] , \in_a_r_reg[1][1] , \in_a_r_reg[1][0] ,
         \in_a_r_reg[2][11] , \in_a_r_reg[2][10] , \in_a_r_reg[2][9] ,
         \in_a_r_reg[2][8] , \in_a_r_reg[2][7] , \in_a_r_reg[2][6] ,
         \in_a_r_reg[2][5] , \in_a_r_reg[2][4] , \in_a_r_reg[2][3] ,
         \in_a_r_reg[2][2] , \in_a_r_reg[2][1] , \in_a_r_reg[2][0] ,
         \in_a_r_reg[3][11] , \in_a_r_reg[3][10] , \in_a_r_reg[3][9] ,
         \in_a_r_reg[3][8] , \in_a_r_reg[3][7] , \in_a_r_reg[3][6] ,
         \in_a_r_reg[3][5] , \in_a_r_reg[3][4] , \in_a_r_reg[3][3] ,
         \in_a_r_reg[3][2] , \in_a_r_reg[3][1] , \in_a_r_reg[3][0] ,
         \in_a_i_reg[0][11] , \in_a_i_reg[0][10] , \in_a_i_reg[0][9] ,
         \in_a_i_reg[0][8] , \in_a_i_reg[0][7] , \in_a_i_reg[0][6] ,
         \in_a_i_reg[0][5] , \in_a_i_reg[0][4] , \in_a_i_reg[0][3] ,
         \in_a_i_reg[0][2] , \in_a_i_reg[0][1] , \in_a_i_reg[0][0] ,
         \in_a_i_reg[1][11] , \in_a_i_reg[1][10] , \in_a_i_reg[1][9] ,
         \in_a_i_reg[1][8] , \in_a_i_reg[1][7] , \in_a_i_reg[1][6] ,
         \in_a_i_reg[1][5] , \in_a_i_reg[1][4] , \in_a_i_reg[1][3] ,
         \in_a_i_reg[1][2] , \in_a_i_reg[1][1] , \in_a_i_reg[1][0] ,
         \in_a_i_reg[2][11] , \in_a_i_reg[2][10] , \in_a_i_reg[2][9] ,
         \in_a_i_reg[2][8] , \in_a_i_reg[2][7] , \in_a_i_reg[2][6] ,
         \in_a_i_reg[2][5] , \in_a_i_reg[2][4] , \in_a_i_reg[2][3] ,
         \in_a_i_reg[2][2] , \in_a_i_reg[2][1] , \in_a_i_reg[2][0] ,
         \in_a_i_reg[3][11] , \in_a_i_reg[3][10] , \in_a_i_reg[3][9] ,
         \in_a_i_reg[3][8] , \in_a_i_reg[3][7] , \in_a_i_reg[3][6] ,
         \in_a_i_reg[3][5] , \in_a_i_reg[3][4] , \in_a_i_reg[3][3] ,
         \in_a_i_reg[3][2] , \in_a_i_reg[3][1] , \in_a_i_reg[3][0] , n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65;
  wire   [11:0] in_b_r_reg;
  wire   [11:0] in_b_i_reg;

  DFFX1 \in_a_r_reg_reg[0][11]  ( .D(\in_a_r[0][11] ), .CLK(clk), .Q(
        \in_a_r_reg[0][11] ) );
  DFFX1 \in_a_r_reg_reg[0][10]  ( .D(\in_a_r[0][10] ), .CLK(clk), .Q(
        \in_a_r_reg[0][10] ) );
  DFFX1 \in_a_r_reg_reg[0][9]  ( .D(\in_a_r[0][9] ), .CLK(clk), .Q(
        \in_a_r_reg[0][9] ) );
  DFFX1 \in_a_r_reg_reg[0][8]  ( .D(\in_a_r[0][8] ), .CLK(clk), .Q(
        \in_a_r_reg[0][8] ) );
  DFFX1 \in_a_r_reg_reg[0][7]  ( .D(\in_a_r[0][7] ), .CLK(clk), .Q(
        \in_a_r_reg[0][7] ) );
  DFFX1 \in_a_r_reg_reg[0][6]  ( .D(\in_a_r[0][6] ), .CLK(clk), .Q(
        \in_a_r_reg[0][6] ) );
  DFFX1 \in_a_r_reg_reg[0][5]  ( .D(\in_a_r[0][5] ), .CLK(clk), .Q(
        \in_a_r_reg[0][5] ) );
  DFFX1 \in_a_r_reg_reg[0][4]  ( .D(\in_a_r[0][4] ), .CLK(clk), .Q(
        \in_a_r_reg[0][4] ) );
  DFFX1 \in_a_r_reg_reg[0][3]  ( .D(\in_a_r[0][3] ), .CLK(clk), .Q(
        \in_a_r_reg[0][3] ) );
  DFFX1 \in_a_r_reg_reg[0][2]  ( .D(\in_a_r[0][2] ), .CLK(clk), .Q(
        \in_a_r_reg[0][2] ) );
  DFFX1 \in_a_r_reg_reg[0][1]  ( .D(\in_a_r[0][1] ), .CLK(clk), .Q(
        \in_a_r_reg[0][1] ) );
  DFFX1 \in_a_r_reg_reg[0][0]  ( .D(\in_a_r[0][0] ), .CLK(clk), .Q(
        \in_a_r_reg[0][0] ) );
  DFFX1 \in_a_r_reg_reg[1][11]  ( .D(\in_a_r[1][11] ), .CLK(clk), .Q(
        \in_a_r_reg[1][11] ) );
  DFFX1 \in_a_r_reg_reg[1][10]  ( .D(\in_a_r[1][10] ), .CLK(clk), .Q(
        \in_a_r_reg[1][10] ) );
  DFFX1 \in_a_r_reg_reg[1][9]  ( .D(\in_a_r[1][9] ), .CLK(clk), .Q(
        \in_a_r_reg[1][9] ) );
  DFFX1 \in_a_r_reg_reg[1][8]  ( .D(\in_a_r[1][8] ), .CLK(clk), .Q(
        \in_a_r_reg[1][8] ) );
  DFFX1 \in_a_r_reg_reg[1][7]  ( .D(\in_a_r[1][7] ), .CLK(clk), .Q(
        \in_a_r_reg[1][7] ) );
  DFFX1 \in_a_r_reg_reg[1][6]  ( .D(\in_a_r[1][6] ), .CLK(clk), .Q(
        \in_a_r_reg[1][6] ) );
  DFFX1 \in_a_r_reg_reg[1][5]  ( .D(\in_a_r[1][5] ), .CLK(clk), .Q(
        \in_a_r_reg[1][5] ) );
  DFFX1 \in_a_r_reg_reg[1][4]  ( .D(\in_a_r[1][4] ), .CLK(clk), .Q(
        \in_a_r_reg[1][4] ) );
  DFFX1 \in_a_r_reg_reg[1][3]  ( .D(\in_a_r[1][3] ), .CLK(clk), .Q(
        \in_a_r_reg[1][3] ) );
  DFFX1 \in_a_r_reg_reg[1][2]  ( .D(\in_a_r[1][2] ), .CLK(clk), .Q(
        \in_a_r_reg[1][2] ) );
  DFFX1 \in_a_r_reg_reg[1][1]  ( .D(\in_a_r[1][1] ), .CLK(clk), .Q(
        \in_a_r_reg[1][1] ) );
  DFFX1 \in_a_r_reg_reg[1][0]  ( .D(\in_a_r[1][0] ), .CLK(clk), .Q(
        \in_a_r_reg[1][0] ) );
  DFFX1 \in_a_r_reg_reg[2][11]  ( .D(\in_a_r[2][11] ), .CLK(clk), .Q(
        \in_a_r_reg[2][11] ) );
  DFFX1 \in_a_r_reg_reg[2][10]  ( .D(\in_a_r[2][10] ), .CLK(clk), .Q(
        \in_a_r_reg[2][10] ) );
  DFFX1 \in_a_r_reg_reg[2][9]  ( .D(\in_a_r[2][9] ), .CLK(clk), .Q(
        \in_a_r_reg[2][9] ) );
  DFFX1 \in_a_r_reg_reg[2][8]  ( .D(\in_a_r[2][8] ), .CLK(clk), .Q(
        \in_a_r_reg[2][8] ) );
  DFFX1 \in_a_r_reg_reg[2][7]  ( .D(\in_a_r[2][7] ), .CLK(clk), .Q(
        \in_a_r_reg[2][7] ) );
  DFFX1 \in_a_r_reg_reg[2][6]  ( .D(\in_a_r[2][6] ), .CLK(clk), .Q(
        \in_a_r_reg[2][6] ) );
  DFFX1 \in_a_r_reg_reg[2][5]  ( .D(\in_a_r[2][5] ), .CLK(clk), .Q(
        \in_a_r_reg[2][5] ) );
  DFFX1 \in_a_r_reg_reg[2][4]  ( .D(\in_a_r[2][4] ), .CLK(clk), .Q(
        \in_a_r_reg[2][4] ) );
  DFFX1 \in_a_r_reg_reg[2][3]  ( .D(\in_a_r[2][3] ), .CLK(clk), .Q(
        \in_a_r_reg[2][3] ) );
  DFFX1 \in_a_r_reg_reg[2][2]  ( .D(\in_a_r[2][2] ), .CLK(clk), .Q(
        \in_a_r_reg[2][2] ) );
  DFFX1 \in_a_r_reg_reg[2][1]  ( .D(\in_a_r[2][1] ), .CLK(clk), .Q(
        \in_a_r_reg[2][1] ) );
  DFFX1 \in_a_r_reg_reg[2][0]  ( .D(\in_a_r[2][0] ), .CLK(clk), .Q(
        \in_a_r_reg[2][0] ) );
  DFFX1 \in_a_r_reg_reg[3][11]  ( .D(\in_a_r[3][11] ), .CLK(clk), .Q(
        \in_a_r_reg[3][11] ) );
  DFFX1 \in_a_r_reg_reg[3][10]  ( .D(\in_a_r[3][10] ), .CLK(clk), .Q(
        \in_a_r_reg[3][10] ) );
  DFFX1 \in_a_r_reg_reg[3][9]  ( .D(\in_a_r[3][9] ), .CLK(clk), .Q(
        \in_a_r_reg[3][9] ) );
  DFFX1 \in_a_r_reg_reg[3][8]  ( .D(\in_a_r[3][8] ), .CLK(clk), .Q(
        \in_a_r_reg[3][8] ) );
  DFFX1 \in_a_r_reg_reg[3][7]  ( .D(\in_a_r[3][7] ), .CLK(clk), .Q(
        \in_a_r_reg[3][7] ) );
  DFFX1 \in_a_r_reg_reg[3][6]  ( .D(\in_a_r[3][6] ), .CLK(clk), .Q(
        \in_a_r_reg[3][6] ) );
  DFFX1 \in_a_r_reg_reg[3][5]  ( .D(\in_a_r[3][5] ), .CLK(clk), .Q(
        \in_a_r_reg[3][5] ) );
  DFFX1 \in_a_r_reg_reg[3][4]  ( .D(\in_a_r[3][4] ), .CLK(clk), .Q(
        \in_a_r_reg[3][4] ) );
  DFFX1 \in_a_r_reg_reg[3][3]  ( .D(\in_a_r[3][3] ), .CLK(clk), .Q(
        \in_a_r_reg[3][3] ) );
  DFFX1 \in_a_r_reg_reg[3][2]  ( .D(\in_a_r[3][2] ), .CLK(clk), .Q(
        \in_a_r_reg[3][2] ) );
  DFFX1 \in_a_r_reg_reg[3][1]  ( .D(\in_a_r[3][1] ), .CLK(clk), .Q(
        \in_a_r_reg[3][1] ) );
  DFFX1 \in_a_r_reg_reg[3][0]  ( .D(\in_a_r[3][0] ), .CLK(clk), .Q(
        \in_a_r_reg[3][0] ) );
  DFFX1 \in_a_i_reg_reg[0][11]  ( .D(\in_a_i[0][11] ), .CLK(clk), .Q(
        \in_a_i_reg[0][11] ) );
  DFFX1 \in_a_i_reg_reg[0][10]  ( .D(\in_a_i[0][10] ), .CLK(clk), .Q(
        \in_a_i_reg[0][10] ) );
  DFFX1 \in_a_i_reg_reg[0][9]  ( .D(\in_a_i[0][9] ), .CLK(clk), .Q(
        \in_a_i_reg[0][9] ) );
  DFFX1 \in_a_i_reg_reg[0][8]  ( .D(\in_a_i[0][8] ), .CLK(clk), .Q(
        \in_a_i_reg[0][8] ) );
  DFFX1 \in_a_i_reg_reg[0][7]  ( .D(\in_a_i[0][7] ), .CLK(clk), .Q(
        \in_a_i_reg[0][7] ) );
  DFFX1 \in_a_i_reg_reg[0][6]  ( .D(\in_a_i[0][6] ), .CLK(clk), .Q(
        \in_a_i_reg[0][6] ) );
  DFFX1 \in_a_i_reg_reg[0][5]  ( .D(\in_a_i[0][5] ), .CLK(clk), .Q(
        \in_a_i_reg[0][5] ) );
  DFFX1 \in_a_i_reg_reg[0][4]  ( .D(\in_a_i[0][4] ), .CLK(clk), .Q(
        \in_a_i_reg[0][4] ) );
  DFFX1 \in_a_i_reg_reg[0][3]  ( .D(\in_a_i[0][3] ), .CLK(clk), .Q(
        \in_a_i_reg[0][3] ) );
  DFFX1 \in_a_i_reg_reg[0][2]  ( .D(\in_a_i[0][2] ), .CLK(clk), .Q(
        \in_a_i_reg[0][2] ) );
  DFFX1 \in_a_i_reg_reg[0][1]  ( .D(\in_a_i[0][1] ), .CLK(clk), .Q(
        \in_a_i_reg[0][1] ) );
  DFFX1 \in_a_i_reg_reg[0][0]  ( .D(\in_a_i[0][0] ), .CLK(clk), .Q(
        \in_a_i_reg[0][0] ) );
  DFFX1 \in_a_i_reg_reg[1][11]  ( .D(\in_a_i[1][11] ), .CLK(clk), .Q(
        \in_a_i_reg[1][11] ) );
  DFFX1 \in_a_i_reg_reg[1][10]  ( .D(\in_a_i[1][10] ), .CLK(clk), .Q(
        \in_a_i_reg[1][10] ) );
  DFFX1 \in_a_i_reg_reg[1][9]  ( .D(\in_a_i[1][9] ), .CLK(clk), .Q(
        \in_a_i_reg[1][9] ) );
  DFFX1 \in_a_i_reg_reg[1][8]  ( .D(\in_a_i[1][8] ), .CLK(clk), .Q(
        \in_a_i_reg[1][8] ) );
  DFFX1 \in_a_i_reg_reg[1][7]  ( .D(\in_a_i[1][7] ), .CLK(clk), .Q(
        \in_a_i_reg[1][7] ) );
  DFFX1 \in_a_i_reg_reg[1][6]  ( .D(\in_a_i[1][6] ), .CLK(clk), .Q(
        \in_a_i_reg[1][6] ) );
  DFFX1 \in_a_i_reg_reg[1][5]  ( .D(\in_a_i[1][5] ), .CLK(clk), .Q(
        \in_a_i_reg[1][5] ) );
  DFFX1 \in_a_i_reg_reg[1][4]  ( .D(\in_a_i[1][4] ), .CLK(clk), .Q(
        \in_a_i_reg[1][4] ) );
  DFFX1 \in_a_i_reg_reg[1][3]  ( .D(\in_a_i[1][3] ), .CLK(clk), .Q(
        \in_a_i_reg[1][3] ) );
  DFFX1 \in_a_i_reg_reg[1][2]  ( .D(\in_a_i[1][2] ), .CLK(clk), .Q(
        \in_a_i_reg[1][2] ) );
  DFFX1 \in_a_i_reg_reg[1][1]  ( .D(\in_a_i[1][1] ), .CLK(clk), .Q(
        \in_a_i_reg[1][1] ) );
  DFFX1 \in_a_i_reg_reg[1][0]  ( .D(\in_a_i[1][0] ), .CLK(clk), .Q(
        \in_a_i_reg[1][0] ) );
  DFFX1 \in_a_i_reg_reg[2][11]  ( .D(\in_a_i[2][11] ), .CLK(clk), .Q(
        \in_a_i_reg[2][11] ) );
  DFFX1 \in_a_i_reg_reg[2][10]  ( .D(\in_a_i[2][10] ), .CLK(clk), .Q(
        \in_a_i_reg[2][10] ) );
  DFFX1 \in_a_i_reg_reg[2][9]  ( .D(\in_a_i[2][9] ), .CLK(clk), .Q(
        \in_a_i_reg[2][9] ) );
  DFFX1 \in_a_i_reg_reg[2][8]  ( .D(\in_a_i[2][8] ), .CLK(clk), .Q(
        \in_a_i_reg[2][8] ) );
  DFFX1 \in_a_i_reg_reg[2][7]  ( .D(\in_a_i[2][7] ), .CLK(clk), .Q(
        \in_a_i_reg[2][7] ) );
  DFFX1 \in_a_i_reg_reg[2][6]  ( .D(\in_a_i[2][6] ), .CLK(clk), .Q(
        \in_a_i_reg[2][6] ) );
  DFFX1 \in_a_i_reg_reg[2][5]  ( .D(\in_a_i[2][5] ), .CLK(clk), .Q(
        \in_a_i_reg[2][5] ) );
  DFFX1 \in_a_i_reg_reg[2][4]  ( .D(\in_a_i[2][4] ), .CLK(clk), .Q(
        \in_a_i_reg[2][4] ) );
  DFFX1 \in_a_i_reg_reg[2][3]  ( .D(\in_a_i[2][3] ), .CLK(clk), .Q(
        \in_a_i_reg[2][3] ) );
  DFFX1 \in_a_i_reg_reg[2][2]  ( .D(\in_a_i[2][2] ), .CLK(clk), .Q(
        \in_a_i_reg[2][2] ) );
  DFFX1 \in_a_i_reg_reg[2][1]  ( .D(\in_a_i[2][1] ), .CLK(clk), .Q(
        \in_a_i_reg[2][1] ) );
  DFFX1 \in_a_i_reg_reg[2][0]  ( .D(\in_a_i[2][0] ), .CLK(clk), .Q(
        \in_a_i_reg[2][0] ) );
  DFFX1 \in_a_i_reg_reg[3][11]  ( .D(\in_a_i[3][11] ), .CLK(clk), .Q(
        \in_a_i_reg[3][11] ) );
  DFFX1 \in_a_i_reg_reg[3][10]  ( .D(\in_a_i[3][10] ), .CLK(clk), .Q(
        \in_a_i_reg[3][10] ) );
  DFFX1 \in_a_i_reg_reg[3][9]  ( .D(\in_a_i[3][9] ), .CLK(clk), .Q(
        \in_a_i_reg[3][9] ) );
  DFFX1 \in_a_i_reg_reg[3][8]  ( .D(\in_a_i[3][8] ), .CLK(clk), .Q(
        \in_a_i_reg[3][8] ) );
  DFFX1 \in_a_i_reg_reg[3][7]  ( .D(\in_a_i[3][7] ), .CLK(clk), .Q(
        \in_a_i_reg[3][7] ) );
  DFFX1 \in_a_i_reg_reg[3][6]  ( .D(\in_a_i[3][6] ), .CLK(clk), .Q(
        \in_a_i_reg[3][6] ) );
  DFFX1 \in_a_i_reg_reg[3][5]  ( .D(\in_a_i[3][5] ), .CLK(clk), .Q(
        \in_a_i_reg[3][5] ) );
  DFFX1 \in_a_i_reg_reg[3][4]  ( .D(\in_a_i[3][4] ), .CLK(clk), .Q(
        \in_a_i_reg[3][4] ) );
  DFFX1 \in_a_i_reg_reg[3][3]  ( .D(\in_a_i[3][3] ), .CLK(clk), .Q(
        \in_a_i_reg[3][3] ) );
  DFFX1 \in_a_i_reg_reg[3][2]  ( .D(\in_a_i[3][2] ), .CLK(clk), .Q(
        \in_a_i_reg[3][2] ) );
  DFFX1 \in_a_i_reg_reg[3][1]  ( .D(\in_a_i[3][1] ), .CLK(clk), .Q(
        \in_a_i_reg[3][1] ) );
  DFFX1 \in_a_i_reg_reg[3][0]  ( .D(\in_a_i[3][0] ), .CLK(clk), .Q(
        \in_a_i_reg[3][0] ) );
  DFFX1 \in_b_r_reg_reg[0]  ( .D(in_b_r[0]), .CLK(clk), .Q(in_b_r_reg[0]) );
  DFFX1 \in_b_i_reg_reg[0]  ( .D(in_b_i[0]), .CLK(clk), .Q(in_b_i_reg[0]), 
        .QN(n1) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_3 mult_0 ( .a_r({
        \in_a_r_reg[0][11] , \in_a_r_reg[0][10] , \in_a_r_reg[0][9] , 
        \in_a_r_reg[0][8] , \in_a_r_reg[0][7] , \in_a_r_reg[0][6] , 
        \in_a_r_reg[0][5] , \in_a_r_reg[0][4] , \in_a_r_reg[0][3] , 
        \in_a_r_reg[0][2] , \in_a_r_reg[0][1] , \in_a_r_reg[0][0] }), .a_i({
        \in_a_i_reg[0][11] , \in_a_i_reg[0][10] , \in_a_i_reg[0][9] , 
        \in_a_i_reg[0][8] , \in_a_i_reg[0][7] , \in_a_i_reg[0][6] , 
        \in_a_i_reg[0][5] , \in_a_i_reg[0][4] , \in_a_i_reg[0][3] , 
        \in_a_i_reg[0][2] , \in_a_i_reg[0][1] , \in_a_i_reg[0][0] }), .b_r({n5, 
        in_b_r_reg[10:9], n10, n4, n53, n45, n55, n61, n41, n43, in_b_r_reg[0]}), .b_i({in_b_i_reg[11], n9, n14, n18, n36, in_b_i_reg[6], n47, n57, 
        in_b_i_reg[3], n13, in_b_i_reg[1], n2}), .out_r({\out_r[0][11] , 
        \out_r[0][10] , \out_r[0][9] , \out_r[0][8] , \out_r[0][7] , 
        \out_r[0][6] , \out_r[0][5] , \out_r[0][4] , \out_r[0][3] , 
        \out_r[0][2] , \out_r[0][1] , \out_r[0][0] }), .out_i({\out_i[0][11] , 
        \out_i[0][10] , \out_i[0][9] , \out_i[0][8] , \out_i[0][7] , 
        \out_i[0][6] , \out_i[0][5] , \out_i[0][4] , \out_i[0][3] , 
        \out_i[0][2] , \out_i[0][1] , \out_i[0][0] }), .clk(clk) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_2 mult_1 ( .a_r({
        \in_a_r_reg[1][11] , \in_a_r_reg[1][10] , \in_a_r_reg[1][9] , 
        \in_a_r_reg[1][8] , \in_a_r_reg[1][7] , \in_a_r_reg[1][6] , 
        \in_a_r_reg[1][5] , \in_a_r_reg[1][4] , \in_a_r_reg[1][3] , 
        \in_a_r_reg[1][2] , \in_a_r_reg[1][1] , \in_a_r_reg[1][0] }), .a_i({
        \in_a_i_reg[1][11] , \in_a_i_reg[1][10] , \in_a_i_reg[1][9] , 
        \in_a_i_reg[1][8] , \in_a_i_reg[1][7] , \in_a_i_reg[1][6] , 
        \in_a_i_reg[1][5] , \in_a_i_reg[1][4] , \in_a_i_reg[1][3] , 
        \in_a_i_reg[1][2] , \in_a_i_reg[1][1] , \in_a_i_reg[1][0] }), .b_r({
        n17, n8, n16, n19, in_b_r_reg[7], n21, in_b_r_reg[5], n32, n34, 
        in_b_r_reg[2:0]}), .b_i({n11, n25, n27, n29, n36, in_b_i_reg[6], n22, 
        in_b_i_reg[4], n59, in_b_i_reg[2:0]}), .out_r({\out_r[1][11] , 
        \out_r[1][10] , \out_r[1][9] , \out_r[1][8] , \out_r[1][7] , 
        \out_r[1][6] , \out_r[1][5] , \out_r[1][4] , \out_r[1][3] , 
        \out_r[1][2] , \out_r[1][1] , \out_r[1][0] }), .out_i({\out_i[1][11] , 
        \out_i[1][10] , \out_i[1][9] , \out_i[1][8] , \out_i[1][7] , 
        \out_i[1][6] , \out_i[1][5] , \out_i[1][4] , \out_i[1][3] , 
        \out_i[1][2] , \out_i[1][1] , \out_i[1][0] }), .clk(clk) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_1 mult_2 ( .a_r({
        \in_a_r_reg[2][11] , \in_a_r_reg[2][10] , \in_a_r_reg[2][9] , 
        \in_a_r_reg[2][8] , \in_a_r_reg[2][7] , \in_a_r_reg[2][6] , 
        \in_a_r_reg[2][5] , \in_a_r_reg[2][4] , \in_a_r_reg[2][3] , 
        \in_a_r_reg[2][2] , \in_a_r_reg[2][1] , \in_a_r_reg[2][0] }), .a_i({
        \in_a_i_reg[2][11] , \in_a_i_reg[2][10] , \in_a_i_reg[2][9] , 
        \in_a_i_reg[2][8] , \in_a_i_reg[2][7] , \in_a_i_reg[2][6] , 
        \in_a_i_reg[2][5] , \in_a_i_reg[2][4] , \in_a_i_reg[2][3] , 
        \in_a_i_reg[2][2] , \in_a_i_reg[2][1] , \in_a_i_reg[2][0] }), .b_r({
        in_b_r_reg[11:6], n45, in_b_r_reg[4:2], n65, in_b_r_reg[0]}), .b_i({
        n38, in_b_i_reg[10:6], n6, in_b_i_reg[4], n20, in_b_i_reg[2], n63, 
        in_b_i_reg[0]}), .out_r({\out_r[2][11] , \out_r[2][10] , \out_r[2][9] , 
        \out_r[2][8] , \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , 
        \out_r[2][4] , \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , 
        \out_r[2][0] }), .out_i({\out_i[2][11] , \out_i[2][10] , \out_i[2][9] , 
        \out_i[2][8] , \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , 
        \out_i[2][4] , \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , 
        \out_i[2][0] }), .clk(clk) );
  complex_mult_pipe_INT_BITS4_WORD_WIDTH12_0 mult_3 ( .a_r({
        \in_a_r_reg[3][11] , \in_a_r_reg[3][10] , \in_a_r_reg[3][9] , 
        \in_a_r_reg[3][8] , \in_a_r_reg[3][7] , \in_a_r_reg[3][6] , 
        \in_a_r_reg[3][5] , \in_a_r_reg[3][4] , \in_a_r_reg[3][3] , 
        \in_a_r_reg[3][2] , \in_a_r_reg[3][1] , \in_a_r_reg[3][0] }), .a_i({
        \in_a_i_reg[3][11] , \in_a_i_reg[3][10] , \in_a_i_reg[3][9] , 
        \in_a_i_reg[3][8] , \in_a_i_reg[3][7] , \in_a_i_reg[3][6] , 
        \in_a_i_reg[3][5] , \in_a_i_reg[3][4] , \in_a_i_reg[3][3] , 
        \in_a_i_reg[3][2] , \in_a_i_reg[3][1] , \in_a_i_reg[3][0] }), .b_r({
        n40, in_b_r_reg[10], n31, n49, in_b_r_reg[7], n15, in_b_r_reg[5:3], 
        n51, n65, in_b_r_reg[0]}), .b_i({in_b_i_reg[11:5], n23, n33, 
        in_b_i_reg[2], n42, in_b_i_reg[0]}), .out_r({\out_r[3][11] , 
        \out_r[3][10] , \out_r[3][9] , \out_r[3][8] , \out_r[3][7] , 
        \out_r[3][6] , \out_r[3][5] , \out_r[3][4] , \out_r[3][3] , 
        \out_r[3][2] , \out_r[3][1] , \out_r[3][0] }), .out_i({\out_i[3][11] , 
        \out_i[3][10] , \out_i[3][9] , \out_i[3][8] , \out_i[3][7] , 
        \out_i[3][6] , \out_i[3][5] , \out_i[3][4] , \out_i[3][3] , 
        \out_i[3][2] , \out_i[3][1] , \out_i[3][0] }), .clk(clk) );
  DFFX1 \in_b_r_reg_reg[2]  ( .D(in_b_r[2]), .CLK(clk), .Q(in_b_r_reg[2]), 
        .QN(n50) );
  DFFX1 \in_b_i_reg_reg[5]  ( .D(in_b_i[5]), .CLK(clk), .Q(in_b_i_reg[5]), 
        .QN(n46) );
  DFFX1 \in_b_r_reg_reg[5]  ( .D(in_b_r[5]), .CLK(clk), .Q(in_b_r_reg[5]), 
        .QN(n44) );
  DFFX1 \in_b_i_reg_reg[7]  ( .D(in_b_i[7]), .CLK(clk), .Q(in_b_i_reg[7]), 
        .QN(n35) );
  DFFX1 \in_b_r_reg_reg[9]  ( .D(in_b_r[9]), .CLK(clk), .Q(in_b_r_reg[9]), 
        .QN(n30) );
  DFFX1 \in_b_i_reg_reg[8]  ( .D(in_b_i[8]), .CLK(clk), .Q(in_b_i_reg[8]), 
        .QN(n28) );
  DFFX1 \in_b_i_reg_reg[9]  ( .D(in_b_i[9]), .CLK(clk), .Q(in_b_i_reg[9]), 
        .QN(n26) );
  DFFX1 \in_b_i_reg_reg[10]  ( .D(in_b_i[10]), .CLK(clk), .Q(in_b_i_reg[10]), 
        .QN(n24) );
  DFFX2 \in_b_i_reg_reg[11]  ( .D(in_b_i[11]), .CLK(clk), .Q(in_b_i_reg[11]), 
        .QN(n37) );
  DFFX1 \in_b_r_reg_reg[10]  ( .D(in_b_r[10]), .CLK(clk), .Q(in_b_r_reg[10]), 
        .QN(n7) );
  DFFX1 \in_b_r_reg_reg[1]  ( .D(in_b_r[1]), .CLK(clk), .Q(in_b_r_reg[1]), 
        .QN(n64) );
  DFFX1 \in_b_i_reg_reg[1]  ( .D(in_b_i[1]), .CLK(clk), .Q(in_b_i_reg[1]), 
        .QN(n62) );
  DFFX1 \in_b_r_reg_reg[3]  ( .D(in_b_r[3]), .CLK(clk), .Q(in_b_r_reg[3]), 
        .QN(n60) );
  DFFX1 \in_b_r_reg_reg[4]  ( .D(in_b_r[4]), .CLK(clk), .Q(in_b_r_reg[4]), 
        .QN(n54) );
  DFFX1 \in_b_i_reg_reg[6]  ( .D(in_b_i[6]), .CLK(clk), .Q(in_b_i_reg[6]) );
  DFFX1 \in_b_i_reg_reg[2]  ( .D(in_b_i[2]), .CLK(clk), .Q(in_b_i_reg[2]), 
        .QN(n12) );
  DFFX1 \in_b_i_reg_reg[3]  ( .D(in_b_i[3]), .CLK(clk), .Q(in_b_i_reg[3]), 
        .QN(n58) );
  DFFX1 \in_b_r_reg_reg[7]  ( .D(in_b_r[7]), .CLK(clk), .Q(in_b_r_reg[7]), 
        .QN(n3) );
  DFFX1 \in_b_i_reg_reg[4]  ( .D(in_b_i[4]), .CLK(clk), .Q(in_b_i_reg[4]), 
        .QN(n56) );
  DFFX1 \in_b_r_reg_reg[11]  ( .D(in_b_r[11]), .CLK(clk), .Q(in_b_r_reg[11]), 
        .QN(n39) );
  DFFX1 \in_b_r_reg_reg[6]  ( .D(in_b_r[6]), .CLK(clk), .Q(in_b_r_reg[6]), 
        .QN(n52) );
  DFFX1 \in_b_r_reg_reg[8]  ( .D(in_b_r[8]), .CLK(clk), .Q(in_b_r_reg[8]), 
        .QN(n48) );
  INVX0 U3 ( .INP(n1), .ZN(n2) );
  INVX0 U4 ( .INP(n3), .ZN(n4) );
  INVX0 U5 ( .INP(n39), .ZN(n5) );
  INVX0 U6 ( .INP(n46), .ZN(n6) );
  INVX0 U7 ( .INP(n7), .ZN(n8) );
  INVX0 U8 ( .INP(n24), .ZN(n9) );
  INVX0 U9 ( .INP(n48), .ZN(n10) );
  INVX0 U10 ( .INP(n37), .ZN(n11) );
  INVX0 U11 ( .INP(n12), .ZN(n13) );
  INVX0 U12 ( .INP(n26), .ZN(n14) );
  INVX0 U13 ( .INP(n52), .ZN(n15) );
  INVX0 U14 ( .INP(n30), .ZN(n16) );
  INVX0 U15 ( .INP(n39), .ZN(n17) );
  INVX0 U16 ( .INP(n28), .ZN(n18) );
  INVX0 U17 ( .INP(n48), .ZN(n19) );
  INVX0 U18 ( .INP(n58), .ZN(n20) );
  INVX0 U19 ( .INP(n52), .ZN(n21) );
  INVX0 U20 ( .INP(n46), .ZN(n22) );
  INVX0 U21 ( .INP(n56), .ZN(n23) );
  INVX0 U22 ( .INP(n24), .ZN(n25) );
  INVX0 U23 ( .INP(n26), .ZN(n27) );
  INVX0 U24 ( .INP(n28), .ZN(n29) );
  INVX0 U25 ( .INP(n30), .ZN(n31) );
  INVX0 U26 ( .INP(n54), .ZN(n32) );
  INVX0 U27 ( .INP(n58), .ZN(n33) );
  INVX0 U28 ( .INP(n60), .ZN(n34) );
  INVX0 U29 ( .INP(n35), .ZN(n36) );
  INVX0 U30 ( .INP(n37), .ZN(n38) );
  INVX0 U31 ( .INP(n39), .ZN(n40) );
  INVX0 U32 ( .INP(n50), .ZN(n41) );
  INVX0 U33 ( .INP(n62), .ZN(n42) );
  INVX0 U34 ( .INP(n64), .ZN(n43) );
  INVX0 U35 ( .INP(n44), .ZN(n45) );
  INVX0 U36 ( .INP(n46), .ZN(n47) );
  INVX0 U37 ( .INP(n48), .ZN(n49) );
  INVX0 U38 ( .INP(n50), .ZN(n51) );
  INVX0 U39 ( .INP(n52), .ZN(n53) );
  INVX0 U40 ( .INP(n54), .ZN(n55) );
  INVX0 U41 ( .INP(n56), .ZN(n57) );
  INVX0 U42 ( .INP(n58), .ZN(n59) );
  INVX0 U43 ( .INP(n60), .ZN(n61) );
  INVX0 U44 ( .INP(n62), .ZN(n63) );
  INVX0 U45 ( .INP(n64), .ZN(n65) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_7_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_7 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_7_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_6_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_6 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_6_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_5_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_5 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_5_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_4_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_4 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_4_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_3_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_3 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_3_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_2_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_2 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_2_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_1_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_1 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_1_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_0_DW01_sub_0 ( A, B, CI, DIFF, 
        CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;
  wire   [12:0] carry;

  FADDX1 U2_10 ( .A(A[10]), .B(n3), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n4), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n5), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n6), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1 U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1 U2_5 ( .A(A[5]), .B(n8), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1 U2_4 ( .A(A[4]), .B(n9), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1 U2_3 ( .A(A[3]), .B(n10), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n11), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n12), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XNOR3X1 U1 ( .IN1(A[11]), .IN2(B[11]), .IN3(carry[11]), .Q(DIFF[11]) );
  INVX0 U2 ( .INP(B[10]), .ZN(n3) );
  INVX0 U3 ( .INP(B[9]), .ZN(n4) );
  INVX0 U4 ( .INP(B[8]), .ZN(n5) );
  INVX0 U5 ( .INP(B[7]), .ZN(n6) );
  INVX0 U6 ( .INP(B[6]), .ZN(n7) );
  INVX0 U7 ( .INP(B[5]), .ZN(n8) );
  INVX0 U8 ( .INP(B[4]), .ZN(n9) );
  INVX0 U9 ( .INP(B[3]), .ZN(n10) );
  INVX0 U10 ( .INP(B[2]), .ZN(n11) );
  INVX0 U11 ( .INP(B[1]), .ZN(n12) );
  NAND2X0 U12 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U13 ( .INP(A[0]), .ZN(n1) );
  INVX0 U14 ( .INP(n13), .ZN(n2) );
  INVX0 U15 ( .INP(B[0]), .ZN(n13) );
  XOR2X1 U16 ( .IN1(n2), .IN2(A[0]), .Q(DIFF[0]) );
endmodule


module add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_0 ( a, b, \output  );
  input [11:0] a;
  input [11:0] b;
  output [11:0] \output ;
  wire   n1, n2, n4, n5, n6, n7;
  wire   [11:0] pre_out;

  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_0_DW01_sub_0 sub_57 ( .A(a), .B(b), 
        .CI(1'b0), .DIFF(pre_out) );
  NAND2X1 U2 ( .IN1(n1), .IN2(n2), .QN(n5) );
  XOR2X1 U3 ( .IN1(pre_out[11]), .IN2(a[11]), .Q(n1) );
  XOR2X1 U4 ( .IN1(b[11]), .IN2(a[11]), .Q(n2) );
  INVX0 U5 ( .INP(n5), .ZN(n6) );
  AND2X1 U6 ( .IN1(n6), .IN2(b[11]), .Q(n4) );
  INVX0 U7 ( .INP(b[11]), .ZN(n7) );
  AO21X1 U8 ( .IN1(pre_out[0]), .IN2(n5), .IN3(n4), .Q(\output [0]) );
  AO21X1 U9 ( .IN1(pre_out[1]), .IN2(n5), .IN3(n4), .Q(\output [1]) );
  AO21X1 U10 ( .IN1(pre_out[2]), .IN2(n5), .IN3(n4), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(pre_out[3]), .IN2(n5), .IN3(n4), .Q(\output [3]) );
  AO21X1 U12 ( .IN1(pre_out[4]), .IN2(n5), .IN3(n4), .Q(\output [4]) );
  AO21X1 U13 ( .IN1(pre_out[5]), .IN2(n5), .IN3(n4), .Q(\output [5]) );
  AO21X1 U14 ( .IN1(pre_out[6]), .IN2(n5), .IN3(n4), .Q(\output [6]) );
  AO21X1 U15 ( .IN1(pre_out[7]), .IN2(n5), .IN3(n4), .Q(\output [7]) );
  AO21X1 U16 ( .IN1(pre_out[8]), .IN2(n5), .IN3(n4), .Q(\output [8]) );
  AO21X1 U17 ( .IN1(pre_out[9]), .IN2(n5), .IN3(n4), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(pre_out[10]), .IN2(n5), .IN3(n4), .Q(\output [10]) );
  MUX21X1 U19 ( .IN1(pre_out[11]), .IN2(n7), .S(n6), .Q(\output [11]) );
endmodule


module vec_sub_N4_WORD_WIDTH12 ( .in_a_r({\in_a_r[0][11] , \in_a_r[0][10] , 
        \in_a_r[0][9] , \in_a_r[0][8] , \in_a_r[0][7] , \in_a_r[0][6] , 
        \in_a_r[0][5] , \in_a_r[0][4] , \in_a_r[0][3] , \in_a_r[0][2] , 
        \in_a_r[0][1] , \in_a_r[0][0] , \in_a_r[1][11] , \in_a_r[1][10] , 
        \in_a_r[1][9] , \in_a_r[1][8] , \in_a_r[1][7] , \in_a_r[1][6] , 
        \in_a_r[1][5] , \in_a_r[1][4] , \in_a_r[1][3] , \in_a_r[1][2] , 
        \in_a_r[1][1] , \in_a_r[1][0] , \in_a_r[2][11] , \in_a_r[2][10] , 
        \in_a_r[2][9] , \in_a_r[2][8] , \in_a_r[2][7] , \in_a_r[2][6] , 
        \in_a_r[2][5] , \in_a_r[2][4] , \in_a_r[2][3] , \in_a_r[2][2] , 
        \in_a_r[2][1] , \in_a_r[2][0] , \in_a_r[3][11] , \in_a_r[3][10] , 
        \in_a_r[3][9] , \in_a_r[3][8] , \in_a_r[3][7] , \in_a_r[3][6] , 
        \in_a_r[3][5] , \in_a_r[3][4] , \in_a_r[3][3] , \in_a_r[3][2] , 
        \in_a_r[3][1] , \in_a_r[3][0] }), .in_a_i({\in_a_i[0][11] , 
        \in_a_i[0][10] , \in_a_i[0][9] , \in_a_i[0][8] , \in_a_i[0][7] , 
        \in_a_i[0][6] , \in_a_i[0][5] , \in_a_i[0][4] , \in_a_i[0][3] , 
        \in_a_i[0][2] , \in_a_i[0][1] , \in_a_i[0][0] , \in_a_i[1][11] , 
        \in_a_i[1][10] , \in_a_i[1][9] , \in_a_i[1][8] , \in_a_i[1][7] , 
        \in_a_i[1][6] , \in_a_i[1][5] , \in_a_i[1][4] , \in_a_i[1][3] , 
        \in_a_i[1][2] , \in_a_i[1][1] , \in_a_i[1][0] , \in_a_i[2][11] , 
        \in_a_i[2][10] , \in_a_i[2][9] , \in_a_i[2][8] , \in_a_i[2][7] , 
        \in_a_i[2][6] , \in_a_i[2][5] , \in_a_i[2][4] , \in_a_i[2][3] , 
        \in_a_i[2][2] , \in_a_i[2][1] , \in_a_i[2][0] , \in_a_i[3][11] , 
        \in_a_i[3][10] , \in_a_i[3][9] , \in_a_i[3][8] , \in_a_i[3][7] , 
        \in_a_i[3][6] , \in_a_i[3][5] , \in_a_i[3][4] , \in_a_i[3][3] , 
        \in_a_i[3][2] , \in_a_i[3][1] , \in_a_i[3][0] }), .in_b_r({
        \in_b_r[0][11] , \in_b_r[0][10] , \in_b_r[0][9] , \in_b_r[0][8] , 
        \in_b_r[0][7] , \in_b_r[0][6] , \in_b_r[0][5] , \in_b_r[0][4] , 
        \in_b_r[0][3] , \in_b_r[0][2] , \in_b_r[0][1] , \in_b_r[0][0] , 
        \in_b_r[1][11] , \in_b_r[1][10] , \in_b_r[1][9] , \in_b_r[1][8] , 
        \in_b_r[1][7] , \in_b_r[1][6] , \in_b_r[1][5] , \in_b_r[1][4] , 
        \in_b_r[1][3] , \in_b_r[1][2] , \in_b_r[1][1] , \in_b_r[1][0] , 
        \in_b_r[2][11] , \in_b_r[2][10] , \in_b_r[2][9] , \in_b_r[2][8] , 
        \in_b_r[2][7] , \in_b_r[2][6] , \in_b_r[2][5] , \in_b_r[2][4] , 
        \in_b_r[2][3] , \in_b_r[2][2] , \in_b_r[2][1] , \in_b_r[2][0] , 
        \in_b_r[3][11] , \in_b_r[3][10] , \in_b_r[3][9] , \in_b_r[3][8] , 
        \in_b_r[3][7] , \in_b_r[3][6] , \in_b_r[3][5] , \in_b_r[3][4] , 
        \in_b_r[3][3] , \in_b_r[3][2] , \in_b_r[3][1] , \in_b_r[3][0] }), 
    .in_b_i({\in_b_i[0][11] , \in_b_i[0][10] , \in_b_i[0][9] , \in_b_i[0][8] , 
        \in_b_i[0][7] , \in_b_i[0][6] , \in_b_i[0][5] , \in_b_i[0][4] , 
        \in_b_i[0][3] , \in_b_i[0][2] , \in_b_i[0][1] , \in_b_i[0][0] , 
        \in_b_i[1][11] , \in_b_i[1][10] , \in_b_i[1][9] , \in_b_i[1][8] , 
        \in_b_i[1][7] , \in_b_i[1][6] , \in_b_i[1][5] , \in_b_i[1][4] , 
        \in_b_i[1][3] , \in_b_i[1][2] , \in_b_i[1][1] , \in_b_i[1][0] , 
        \in_b_i[2][11] , \in_b_i[2][10] , \in_b_i[2][9] , \in_b_i[2][8] , 
        \in_b_i[2][7] , \in_b_i[2][6] , \in_b_i[2][5] , \in_b_i[2][4] , 
        \in_b_i[2][3] , \in_b_i[2][2] , \in_b_i[2][1] , \in_b_i[2][0] , 
        \in_b_i[3][11] , \in_b_i[3][10] , \in_b_i[3][9] , \in_b_i[3][8] , 
        \in_b_i[3][7] , \in_b_i[3][6] , \in_b_i[3][5] , \in_b_i[3][4] , 
        \in_b_i[3][3] , \in_b_i[3][2] , \in_b_i[3][1] , \in_b_i[3][0] }), 
    .out_r({\out_r[0][11] , \out_r[0][10] , \out_r[0][9] , \out_r[0][8] , 
        \out_r[0][7] , \out_r[0][6] , \out_r[0][5] , \out_r[0][4] , 
        \out_r[0][3] , \out_r[0][2] , \out_r[0][1] , \out_r[0][0] , 
        \out_r[1][11] , \out_r[1][10] , \out_r[1][9] , \out_r[1][8] , 
        \out_r[1][7] , \out_r[1][6] , \out_r[1][5] , \out_r[1][4] , 
        \out_r[1][3] , \out_r[1][2] , \out_r[1][1] , \out_r[1][0] , 
        \out_r[2][11] , \out_r[2][10] , \out_r[2][9] , \out_r[2][8] , 
        \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , \out_r[2][4] , 
        \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , \out_r[2][0] , 
        \out_r[3][11] , \out_r[3][10] , \out_r[3][9] , \out_r[3][8] , 
        \out_r[3][7] , \out_r[3][6] , \out_r[3][5] , \out_r[3][4] , 
        \out_r[3][3] , \out_r[3][2] , \out_r[3][1] , \out_r[3][0] }), .out_i({
        \out_i[0][11] , \out_i[0][10] , \out_i[0][9] , \out_i[0][8] , 
        \out_i[0][7] , \out_i[0][6] , \out_i[0][5] , \out_i[0][4] , 
        \out_i[0][3] , \out_i[0][2] , \out_i[0][1] , \out_i[0][0] , 
        \out_i[1][11] , \out_i[1][10] , \out_i[1][9] , \out_i[1][8] , 
        \out_i[1][7] , \out_i[1][6] , \out_i[1][5] , \out_i[1][4] , 
        \out_i[1][3] , \out_i[1][2] , \out_i[1][1] , \out_i[1][0] , 
        \out_i[2][11] , \out_i[2][10] , \out_i[2][9] , \out_i[2][8] , 
        \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , \out_i[2][4] , 
        \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , \out_i[2][0] , 
        \out_i[3][11] , \out_i[3][10] , \out_i[3][9] , \out_i[3][8] , 
        \out_i[3][7] , \out_i[3][6] , \out_i[3][5] , \out_i[3][4] , 
        \out_i[3][3] , \out_i[3][2] , \out_i[3][1] , \out_i[3][0] }), w_in_a, 
        clk );
  input \in_a_r[0][11] , \in_a_r[0][10] , \in_a_r[0][9] , \in_a_r[0][8] ,
         \in_a_r[0][7] , \in_a_r[0][6] , \in_a_r[0][5] , \in_a_r[0][4] ,
         \in_a_r[0][3] , \in_a_r[0][2] , \in_a_r[0][1] , \in_a_r[0][0] ,
         \in_a_r[1][11] , \in_a_r[1][10] , \in_a_r[1][9] , \in_a_r[1][8] ,
         \in_a_r[1][7] , \in_a_r[1][6] , \in_a_r[1][5] , \in_a_r[1][4] ,
         \in_a_r[1][3] , \in_a_r[1][2] , \in_a_r[1][1] , \in_a_r[1][0] ,
         \in_a_r[2][11] , \in_a_r[2][10] , \in_a_r[2][9] , \in_a_r[2][8] ,
         \in_a_r[2][7] , \in_a_r[2][6] , \in_a_r[2][5] , \in_a_r[2][4] ,
         \in_a_r[2][3] , \in_a_r[2][2] , \in_a_r[2][1] , \in_a_r[2][0] ,
         \in_a_r[3][11] , \in_a_r[3][10] , \in_a_r[3][9] , \in_a_r[3][8] ,
         \in_a_r[3][7] , \in_a_r[3][6] , \in_a_r[3][5] , \in_a_r[3][4] ,
         \in_a_r[3][3] , \in_a_r[3][2] , \in_a_r[3][1] , \in_a_r[3][0] ,
         \in_a_i[0][11] , \in_a_i[0][10] , \in_a_i[0][9] , \in_a_i[0][8] ,
         \in_a_i[0][7] , \in_a_i[0][6] , \in_a_i[0][5] , \in_a_i[0][4] ,
         \in_a_i[0][3] , \in_a_i[0][2] , \in_a_i[0][1] , \in_a_i[0][0] ,
         \in_a_i[1][11] , \in_a_i[1][10] , \in_a_i[1][9] , \in_a_i[1][8] ,
         \in_a_i[1][7] , \in_a_i[1][6] , \in_a_i[1][5] , \in_a_i[1][4] ,
         \in_a_i[1][3] , \in_a_i[1][2] , \in_a_i[1][1] , \in_a_i[1][0] ,
         \in_a_i[2][11] , \in_a_i[2][10] , \in_a_i[2][9] , \in_a_i[2][8] ,
         \in_a_i[2][7] , \in_a_i[2][6] , \in_a_i[2][5] , \in_a_i[2][4] ,
         \in_a_i[2][3] , \in_a_i[2][2] , \in_a_i[2][1] , \in_a_i[2][0] ,
         \in_a_i[3][11] , \in_a_i[3][10] , \in_a_i[3][9] , \in_a_i[3][8] ,
         \in_a_i[3][7] , \in_a_i[3][6] , \in_a_i[3][5] , \in_a_i[3][4] ,
         \in_a_i[3][3] , \in_a_i[3][2] , \in_a_i[3][1] , \in_a_i[3][0] ,
         \in_b_r[0][11] , \in_b_r[0][10] , \in_b_r[0][9] , \in_b_r[0][8] ,
         \in_b_r[0][7] , \in_b_r[0][6] , \in_b_r[0][5] , \in_b_r[0][4] ,
         \in_b_r[0][3] , \in_b_r[0][2] , \in_b_r[0][1] , \in_b_r[0][0] ,
         \in_b_r[1][11] , \in_b_r[1][10] , \in_b_r[1][9] , \in_b_r[1][8] ,
         \in_b_r[1][7] , \in_b_r[1][6] , \in_b_r[1][5] , \in_b_r[1][4] ,
         \in_b_r[1][3] , \in_b_r[1][2] , \in_b_r[1][1] , \in_b_r[1][0] ,
         \in_b_r[2][11] , \in_b_r[2][10] , \in_b_r[2][9] , \in_b_r[2][8] ,
         \in_b_r[2][7] , \in_b_r[2][6] , \in_b_r[2][5] , \in_b_r[2][4] ,
         \in_b_r[2][3] , \in_b_r[2][2] , \in_b_r[2][1] , \in_b_r[2][0] ,
         \in_b_r[3][11] , \in_b_r[3][10] , \in_b_r[3][9] , \in_b_r[3][8] ,
         \in_b_r[3][7] , \in_b_r[3][6] , \in_b_r[3][5] , \in_b_r[3][4] ,
         \in_b_r[3][3] , \in_b_r[3][2] , \in_b_r[3][1] , \in_b_r[3][0] ,
         \in_b_i[0][11] , \in_b_i[0][10] , \in_b_i[0][9] , \in_b_i[0][8] ,
         \in_b_i[0][7] , \in_b_i[0][6] , \in_b_i[0][5] , \in_b_i[0][4] ,
         \in_b_i[0][3] , \in_b_i[0][2] , \in_b_i[0][1] , \in_b_i[0][0] ,
         \in_b_i[1][11] , \in_b_i[1][10] , \in_b_i[1][9] , \in_b_i[1][8] ,
         \in_b_i[1][7] , \in_b_i[1][6] , \in_b_i[1][5] , \in_b_i[1][4] ,
         \in_b_i[1][3] , \in_b_i[1][2] , \in_b_i[1][1] , \in_b_i[1][0] ,
         \in_b_i[2][11] , \in_b_i[2][10] , \in_b_i[2][9] , \in_b_i[2][8] ,
         \in_b_i[2][7] , \in_b_i[2][6] , \in_b_i[2][5] , \in_b_i[2][4] ,
         \in_b_i[2][3] , \in_b_i[2][2] , \in_b_i[2][1] , \in_b_i[2][0] ,
         \in_b_i[3][11] , \in_b_i[3][10] , \in_b_i[3][9] , \in_b_i[3][8] ,
         \in_b_i[3][7] , \in_b_i[3][6] , \in_b_i[3][5] , \in_b_i[3][4] ,
         \in_b_i[3][3] , \in_b_i[3][2] , \in_b_i[3][1] , \in_b_i[3][0] ,
         w_in_a, clk;
  output \out_r[0][11] , \out_r[0][10] , \out_r[0][9] , \out_r[0][8] ,
         \out_r[0][7] , \out_r[0][6] , \out_r[0][5] , \out_r[0][4] ,
         \out_r[0][3] , \out_r[0][2] , \out_r[0][1] , \out_r[0][0] ,
         \out_r[1][11] , \out_r[1][10] , \out_r[1][9] , \out_r[1][8] ,
         \out_r[1][7] , \out_r[1][6] , \out_r[1][5] , \out_r[1][4] ,
         \out_r[1][3] , \out_r[1][2] , \out_r[1][1] , \out_r[1][0] ,
         \out_r[2][11] , \out_r[2][10] , \out_r[2][9] , \out_r[2][8] ,
         \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , \out_r[2][4] ,
         \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , \out_r[2][0] ,
         \out_r[3][11] , \out_r[3][10] , \out_r[3][9] , \out_r[3][8] ,
         \out_r[3][7] , \out_r[3][6] , \out_r[3][5] , \out_r[3][4] ,
         \out_r[3][3] , \out_r[3][2] , \out_r[3][1] , \out_r[3][0] ,
         \out_i[0][11] , \out_i[0][10] , \out_i[0][9] , \out_i[0][8] ,
         \out_i[0][7] , \out_i[0][6] , \out_i[0][5] , \out_i[0][4] ,
         \out_i[0][3] , \out_i[0][2] , \out_i[0][1] , \out_i[0][0] ,
         \out_i[1][11] , \out_i[1][10] , \out_i[1][9] , \out_i[1][8] ,
         \out_i[1][7] , \out_i[1][6] , \out_i[1][5] , \out_i[1][4] ,
         \out_i[1][3] , \out_i[1][2] , \out_i[1][1] , \out_i[1][0] ,
         \out_i[2][11] , \out_i[2][10] , \out_i[2][9] , \out_i[2][8] ,
         \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , \out_i[2][4] ,
         \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , \out_i[2][0] ,
         \out_i[3][11] , \out_i[3][10] , \out_i[3][9] , \out_i[3][8] ,
         \out_i[3][7] , \out_i[3][6] , \out_i[3][5] , \out_i[3][4] ,
         \out_i[3][3] , \out_i[3][2] , \out_i[3][1] , \out_i[3][0] ;
  wire   \in_a_r_reg[0][11] , \in_a_r_reg[0][10] , \in_a_r_reg[0][9] ,
         \in_a_r_reg[0][8] , \in_a_r_reg[0][7] , \in_a_r_reg[0][6] ,
         \in_a_r_reg[0][5] , \in_a_r_reg[0][4] , \in_a_r_reg[0][3] ,
         \in_a_r_reg[0][2] , \in_a_r_reg[0][1] , \in_a_r_reg[0][0] ,
         \in_a_r_reg[1][11] , \in_a_r_reg[1][10] , \in_a_r_reg[1][9] ,
         \in_a_r_reg[1][8] , \in_a_r_reg[1][7] , \in_a_r_reg[1][6] ,
         \in_a_r_reg[1][5] , \in_a_r_reg[1][4] , \in_a_r_reg[1][3] ,
         \in_a_r_reg[1][2] , \in_a_r_reg[1][1] , \in_a_r_reg[1][0] ,
         \in_a_r_reg[2][11] , \in_a_r_reg[2][10] , \in_a_r_reg[2][9] ,
         \in_a_r_reg[2][8] , \in_a_r_reg[2][7] , \in_a_r_reg[2][6] ,
         \in_a_r_reg[2][5] , \in_a_r_reg[2][4] , \in_a_r_reg[2][3] ,
         \in_a_r_reg[2][2] , \in_a_r_reg[2][1] , \in_a_r_reg[2][0] ,
         \in_a_r_reg[3][11] , \in_a_r_reg[3][10] , \in_a_r_reg[3][9] ,
         \in_a_r_reg[3][8] , \in_a_r_reg[3][7] , \in_a_r_reg[3][6] ,
         \in_a_r_reg[3][5] , \in_a_r_reg[3][4] , \in_a_r_reg[3][3] ,
         \in_a_r_reg[3][2] , \in_a_r_reg[3][1] , \in_a_r_reg[3][0] ,
         \in_a_i_reg[0][11] , \in_a_i_reg[0][10] , \in_a_i_reg[0][9] ,
         \in_a_i_reg[0][8] , \in_a_i_reg[0][7] , \in_a_i_reg[0][6] ,
         \in_a_i_reg[0][5] , \in_a_i_reg[0][4] , \in_a_i_reg[0][3] ,
         \in_a_i_reg[0][2] , \in_a_i_reg[0][1] , \in_a_i_reg[0][0] ,
         \in_a_i_reg[1][11] , \in_a_i_reg[1][10] , \in_a_i_reg[1][9] ,
         \in_a_i_reg[1][8] , \in_a_i_reg[1][7] , \in_a_i_reg[1][6] ,
         \in_a_i_reg[1][5] , \in_a_i_reg[1][4] , \in_a_i_reg[1][3] ,
         \in_a_i_reg[1][2] , \in_a_i_reg[1][1] , \in_a_i_reg[1][0] ,
         \in_a_i_reg[2][11] , \in_a_i_reg[2][10] , \in_a_i_reg[2][9] ,
         \in_a_i_reg[2][8] , \in_a_i_reg[2][7] , \in_a_i_reg[2][6] ,
         \in_a_i_reg[2][5] , \in_a_i_reg[2][4] , \in_a_i_reg[2][3] ,
         \in_a_i_reg[2][2] , \in_a_i_reg[2][1] , \in_a_i_reg[2][0] ,
         \in_a_i_reg[3][11] , \in_a_i_reg[3][10] , \in_a_i_reg[3][9] ,
         \in_a_i_reg[3][8] , \in_a_i_reg[3][7] , \in_a_i_reg[3][6] ,
         \in_a_i_reg[3][5] , \in_a_i_reg[3][4] , \in_a_i_reg[3][3] ,
         \in_a_i_reg[3][2] , \in_a_i_reg[3][1] , \in_a_i_reg[3][0] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n1, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115;

  DFFX1 \in_a_i_reg_reg[0][11]  ( .D(n97), .CLK(clk), .Q(\in_a_i_reg[0][11] )
         );
  DFFX1 \in_a_i_reg_reg[0][10]  ( .D(n96), .CLK(clk), .Q(\in_a_i_reg[0][10] )
         );
  DFFX1 \in_a_i_reg_reg[0][9]  ( .D(n95), .CLK(clk), .Q(\in_a_i_reg[0][9] ) );
  DFFX1 \in_a_i_reg_reg[0][8]  ( .D(n94), .CLK(clk), .Q(\in_a_i_reg[0][8] ) );
  DFFX1 \in_a_i_reg_reg[0][7]  ( .D(n93), .CLK(clk), .Q(\in_a_i_reg[0][7] ) );
  DFFX1 \in_a_i_reg_reg[0][6]  ( .D(n92), .CLK(clk), .Q(\in_a_i_reg[0][6] ) );
  DFFX1 \in_a_i_reg_reg[0][5]  ( .D(n91), .CLK(clk), .Q(\in_a_i_reg[0][5] ) );
  DFFX1 \in_a_i_reg_reg[0][4]  ( .D(n90), .CLK(clk), .Q(\in_a_i_reg[0][4] ) );
  DFFX1 \in_a_i_reg_reg[0][3]  ( .D(n89), .CLK(clk), .Q(\in_a_i_reg[0][3] ) );
  DFFX1 \in_a_i_reg_reg[0][2]  ( .D(n88), .CLK(clk), .Q(\in_a_i_reg[0][2] ) );
  DFFX1 \in_a_i_reg_reg[0][1]  ( .D(n87), .CLK(clk), .Q(\in_a_i_reg[0][1] ) );
  DFFX1 \in_a_i_reg_reg[0][0]  ( .D(n86), .CLK(clk), .Q(\in_a_i_reg[0][0] ) );
  DFFX1 \in_a_i_reg_reg[1][11]  ( .D(n85), .CLK(clk), .Q(\in_a_i_reg[1][11] )
         );
  DFFX1 \in_a_i_reg_reg[1][10]  ( .D(n84), .CLK(clk), .Q(\in_a_i_reg[1][10] )
         );
  DFFX1 \in_a_i_reg_reg[1][9]  ( .D(n83), .CLK(clk), .Q(\in_a_i_reg[1][9] ) );
  DFFX1 \in_a_i_reg_reg[1][8]  ( .D(n82), .CLK(clk), .Q(\in_a_i_reg[1][8] ) );
  DFFX1 \in_a_i_reg_reg[1][7]  ( .D(n81), .CLK(clk), .Q(\in_a_i_reg[1][7] ) );
  DFFX1 \in_a_i_reg_reg[1][6]  ( .D(n80), .CLK(clk), .Q(\in_a_i_reg[1][6] ) );
  DFFX1 \in_a_i_reg_reg[1][5]  ( .D(n79), .CLK(clk), .Q(\in_a_i_reg[1][5] ) );
  DFFX1 \in_a_i_reg_reg[1][4]  ( .D(n78), .CLK(clk), .Q(\in_a_i_reg[1][4] ) );
  DFFX1 \in_a_i_reg_reg[1][3]  ( .D(n77), .CLK(clk), .Q(\in_a_i_reg[1][3] ) );
  DFFX1 \in_a_i_reg_reg[1][2]  ( .D(n76), .CLK(clk), .Q(\in_a_i_reg[1][2] ) );
  DFFX1 \in_a_i_reg_reg[1][1]  ( .D(n75), .CLK(clk), .Q(\in_a_i_reg[1][1] ) );
  DFFX1 \in_a_i_reg_reg[1][0]  ( .D(n74), .CLK(clk), .Q(\in_a_i_reg[1][0] ) );
  DFFX1 \in_a_i_reg_reg[2][11]  ( .D(n73), .CLK(clk), .Q(\in_a_i_reg[2][11] )
         );
  DFFX1 \in_a_i_reg_reg[2][10]  ( .D(n72), .CLK(clk), .Q(\in_a_i_reg[2][10] )
         );
  DFFX1 \in_a_i_reg_reg[2][9]  ( .D(n71), .CLK(clk), .Q(\in_a_i_reg[2][9] ) );
  DFFX1 \in_a_i_reg_reg[2][8]  ( .D(n70), .CLK(clk), .Q(\in_a_i_reg[2][8] ) );
  DFFX1 \in_a_i_reg_reg[2][7]  ( .D(n69), .CLK(clk), .Q(\in_a_i_reg[2][7] ) );
  DFFX1 \in_a_i_reg_reg[2][6]  ( .D(n68), .CLK(clk), .Q(\in_a_i_reg[2][6] ) );
  DFFX1 \in_a_i_reg_reg[2][5]  ( .D(n67), .CLK(clk), .Q(\in_a_i_reg[2][5] ) );
  DFFX1 \in_a_i_reg_reg[2][4]  ( .D(n66), .CLK(clk), .Q(\in_a_i_reg[2][4] ) );
  DFFX1 \in_a_i_reg_reg[2][3]  ( .D(n65), .CLK(clk), .Q(\in_a_i_reg[2][3] ) );
  DFFX1 \in_a_i_reg_reg[2][2]  ( .D(n64), .CLK(clk), .Q(\in_a_i_reg[2][2] ) );
  DFFX1 \in_a_i_reg_reg[2][1]  ( .D(n63), .CLK(clk), .Q(\in_a_i_reg[2][1] ) );
  DFFX1 \in_a_i_reg_reg[2][0]  ( .D(n62), .CLK(clk), .Q(\in_a_i_reg[2][0] ) );
  DFFX1 \in_a_i_reg_reg[3][11]  ( .D(n61), .CLK(clk), .Q(\in_a_i_reg[3][11] )
         );
  DFFX1 \in_a_i_reg_reg[3][10]  ( .D(n60), .CLK(clk), .Q(\in_a_i_reg[3][10] )
         );
  DFFX1 \in_a_i_reg_reg[3][9]  ( .D(n59), .CLK(clk), .Q(\in_a_i_reg[3][9] ) );
  DFFX1 \in_a_i_reg_reg[3][8]  ( .D(n58), .CLK(clk), .Q(\in_a_i_reg[3][8] ) );
  DFFX1 \in_a_i_reg_reg[3][7]  ( .D(n57), .CLK(clk), .Q(\in_a_i_reg[3][7] ) );
  DFFX1 \in_a_i_reg_reg[3][6]  ( .D(n56), .CLK(clk), .Q(\in_a_i_reg[3][6] ) );
  DFFX1 \in_a_i_reg_reg[3][5]  ( .D(n55), .CLK(clk), .Q(\in_a_i_reg[3][5] ) );
  DFFX1 \in_a_i_reg_reg[3][4]  ( .D(n54), .CLK(clk), .Q(\in_a_i_reg[3][4] ) );
  DFFX1 \in_a_i_reg_reg[3][3]  ( .D(n53), .CLK(clk), .Q(\in_a_i_reg[3][3] ) );
  DFFX1 \in_a_i_reg_reg[3][2]  ( .D(n52), .CLK(clk), .Q(\in_a_i_reg[3][2] ) );
  DFFX1 \in_a_i_reg_reg[3][1]  ( .D(n51), .CLK(clk), .Q(\in_a_i_reg[3][1] ) );
  DFFX1 \in_a_i_reg_reg[3][0]  ( .D(n50), .CLK(clk), .Q(\in_a_i_reg[3][0] ) );
  DFFX1 \in_a_r_reg_reg[0][11]  ( .D(n49), .CLK(clk), .Q(\in_a_r_reg[0][11] )
         );
  DFFX1 \in_a_r_reg_reg[0][10]  ( .D(n48), .CLK(clk), .Q(\in_a_r_reg[0][10] )
         );
  DFFX1 \in_a_r_reg_reg[0][9]  ( .D(n47), .CLK(clk), .Q(\in_a_r_reg[0][9] ) );
  DFFX1 \in_a_r_reg_reg[0][8]  ( .D(n46), .CLK(clk), .Q(\in_a_r_reg[0][8] ) );
  DFFX1 \in_a_r_reg_reg[0][7]  ( .D(n45), .CLK(clk), .Q(\in_a_r_reg[0][7] ) );
  DFFX1 \in_a_r_reg_reg[0][6]  ( .D(n44), .CLK(clk), .Q(\in_a_r_reg[0][6] ) );
  DFFX1 \in_a_r_reg_reg[0][5]  ( .D(n43), .CLK(clk), .Q(\in_a_r_reg[0][5] ) );
  DFFX1 \in_a_r_reg_reg[0][4]  ( .D(n42), .CLK(clk), .Q(\in_a_r_reg[0][4] ) );
  DFFX1 \in_a_r_reg_reg[0][3]  ( .D(n41), .CLK(clk), .Q(\in_a_r_reg[0][3] ) );
  DFFX1 \in_a_r_reg_reg[0][2]  ( .D(n40), .CLK(clk), .Q(\in_a_r_reg[0][2] ) );
  DFFX1 \in_a_r_reg_reg[0][1]  ( .D(n39), .CLK(clk), .Q(\in_a_r_reg[0][1] ) );
  DFFX1 \in_a_r_reg_reg[0][0]  ( .D(n38), .CLK(clk), .Q(\in_a_r_reg[0][0] ) );
  DFFX1 \in_a_r_reg_reg[1][11]  ( .D(n37), .CLK(clk), .Q(\in_a_r_reg[1][11] )
         );
  DFFX1 \in_a_r_reg_reg[1][10]  ( .D(n36), .CLK(clk), .Q(\in_a_r_reg[1][10] )
         );
  DFFX1 \in_a_r_reg_reg[1][9]  ( .D(n35), .CLK(clk), .Q(\in_a_r_reg[1][9] ) );
  DFFX1 \in_a_r_reg_reg[1][8]  ( .D(n34), .CLK(clk), .Q(\in_a_r_reg[1][8] ) );
  DFFX1 \in_a_r_reg_reg[1][7]  ( .D(n33), .CLK(clk), .Q(\in_a_r_reg[1][7] ) );
  DFFX1 \in_a_r_reg_reg[1][6]  ( .D(n32), .CLK(clk), .Q(\in_a_r_reg[1][6] ) );
  DFFX1 \in_a_r_reg_reg[1][5]  ( .D(n31), .CLK(clk), .Q(\in_a_r_reg[1][5] ) );
  DFFX1 \in_a_r_reg_reg[1][4]  ( .D(n30), .CLK(clk), .Q(\in_a_r_reg[1][4] ) );
  DFFX1 \in_a_r_reg_reg[1][3]  ( .D(n29), .CLK(clk), .Q(\in_a_r_reg[1][3] ) );
  DFFX1 \in_a_r_reg_reg[1][2]  ( .D(n28), .CLK(clk), .Q(\in_a_r_reg[1][2] ) );
  DFFX1 \in_a_r_reg_reg[1][1]  ( .D(n27), .CLK(clk), .Q(\in_a_r_reg[1][1] ) );
  DFFX1 \in_a_r_reg_reg[1][0]  ( .D(n26), .CLK(clk), .Q(\in_a_r_reg[1][0] ) );
  DFFX1 \in_a_r_reg_reg[2][11]  ( .D(n25), .CLK(clk), .Q(\in_a_r_reg[2][11] )
         );
  DFFX1 \in_a_r_reg_reg[2][10]  ( .D(n24), .CLK(clk), .Q(\in_a_r_reg[2][10] )
         );
  DFFX1 \in_a_r_reg_reg[2][9]  ( .D(n23), .CLK(clk), .Q(\in_a_r_reg[2][9] ) );
  DFFX1 \in_a_r_reg_reg[2][8]  ( .D(n22), .CLK(clk), .Q(\in_a_r_reg[2][8] ) );
  DFFX1 \in_a_r_reg_reg[2][7]  ( .D(n21), .CLK(clk), .Q(\in_a_r_reg[2][7] ) );
  DFFX1 \in_a_r_reg_reg[2][6]  ( .D(n20), .CLK(clk), .Q(\in_a_r_reg[2][6] ) );
  DFFX1 \in_a_r_reg_reg[2][5]  ( .D(n19), .CLK(clk), .Q(\in_a_r_reg[2][5] ) );
  DFFX1 \in_a_r_reg_reg[2][4]  ( .D(n18), .CLK(clk), .Q(\in_a_r_reg[2][4] ) );
  DFFX1 \in_a_r_reg_reg[2][3]  ( .D(n17), .CLK(clk), .Q(\in_a_r_reg[2][3] ) );
  DFFX1 \in_a_r_reg_reg[2][2]  ( .D(n16), .CLK(clk), .Q(\in_a_r_reg[2][2] ) );
  DFFX1 \in_a_r_reg_reg[2][1]  ( .D(n15), .CLK(clk), .Q(\in_a_r_reg[2][1] ) );
  DFFX1 \in_a_r_reg_reg[2][0]  ( .D(n14), .CLK(clk), .Q(\in_a_r_reg[2][0] ) );
  DFFX1 \in_a_r_reg_reg[3][11]  ( .D(n13), .CLK(clk), .Q(\in_a_r_reg[3][11] )
         );
  DFFX1 \in_a_r_reg_reg[3][10]  ( .D(n12), .CLK(clk), .Q(\in_a_r_reg[3][10] )
         );
  DFFX1 \in_a_r_reg_reg[3][9]  ( .D(n11), .CLK(clk), .Q(\in_a_r_reg[3][9] ) );
  DFFX1 \in_a_r_reg_reg[3][8]  ( .D(n10), .CLK(clk), .Q(\in_a_r_reg[3][8] ) );
  DFFX1 \in_a_r_reg_reg[3][7]  ( .D(n9), .CLK(clk), .Q(\in_a_r_reg[3][7] ) );
  DFFX1 \in_a_r_reg_reg[3][6]  ( .D(n8), .CLK(clk), .Q(\in_a_r_reg[3][6] ) );
  DFFX1 \in_a_r_reg_reg[3][5]  ( .D(n7), .CLK(clk), .Q(\in_a_r_reg[3][5] ) );
  DFFX1 \in_a_r_reg_reg[3][4]  ( .D(n6), .CLK(clk), .Q(\in_a_r_reg[3][4] ) );
  DFFX1 \in_a_r_reg_reg[3][3]  ( .D(n5), .CLK(clk), .Q(\in_a_r_reg[3][3] ) );
  DFFX1 \in_a_r_reg_reg[3][2]  ( .D(n4), .CLK(clk), .Q(\in_a_r_reg[3][2] ) );
  DFFX1 \in_a_r_reg_reg[3][1]  ( .D(n3), .CLK(clk), .Q(\in_a_r_reg[3][1] ) );
  DFFX1 \in_a_r_reg_reg[3][0]  ( .D(n2), .CLK(clk), .Q(\in_a_r_reg[3][0] ) );
  AO22X1 U3 ( .IN1(\in_a_r_reg[3][1] ), .IN2(n102), .IN3(\in_a_r[3][1] ), 
        .IN4(n1), .Q(n3) );
  AO22X1 U4 ( .IN1(\in_a_r_reg[3][2] ), .IN2(n103), .IN3(\in_a_r[3][2] ), 
        .IN4(n1), .Q(n4) );
  AO22X1 U5 ( .IN1(\in_a_r_reg[3][3] ), .IN2(n103), .IN3(\in_a_r[3][3] ), 
        .IN4(n1), .Q(n5) );
  AO22X1 U6 ( .IN1(\in_a_r_reg[3][4] ), .IN2(n103), .IN3(\in_a_r[3][4] ), 
        .IN4(n1), .Q(n6) );
  AO22X1 U7 ( .IN1(\in_a_r_reg[3][5] ), .IN2(n103), .IN3(\in_a_r[3][5] ), 
        .IN4(n98), .Q(n7) );
  AO22X1 U8 ( .IN1(\in_a_r_reg[3][6] ), .IN2(n103), .IN3(\in_a_r[3][6] ), 
        .IN4(n98), .Q(n8) );
  AO22X1 U9 ( .IN1(\in_a_r_reg[3][7] ), .IN2(n103), .IN3(\in_a_r[3][7] ), 
        .IN4(n98), .Q(n9) );
  AO22X1 U10 ( .IN1(\in_a_r_reg[3][8] ), .IN2(n103), .IN3(\in_a_r[3][8] ), 
        .IN4(n98), .Q(n10) );
  AO22X1 U11 ( .IN1(\in_a_r_reg[3][9] ), .IN2(n104), .IN3(\in_a_r[3][9] ), 
        .IN4(n98), .Q(n11) );
  AO22X1 U12 ( .IN1(\in_a_r_reg[3][10] ), .IN2(n104), .IN3(\in_a_r[3][10] ), 
        .IN4(n98), .Q(n12) );
  AO22X1 U13 ( .IN1(\in_a_r_reg[3][11] ), .IN2(n104), .IN3(\in_a_r[3][11] ), 
        .IN4(n98), .Q(n13) );
  AO22X1 U15 ( .IN1(\in_a_r_reg[2][1] ), .IN2(n104), .IN3(\in_a_r[2][1] ), 
        .IN4(n98), .Q(n15) );
  AO22X1 U16 ( .IN1(\in_a_r_reg[2][2] ), .IN2(n104), .IN3(\in_a_r[2][2] ), 
        .IN4(n98), .Q(n16) );
  AO22X1 U17 ( .IN1(\in_a_r_reg[2][3] ), .IN2(n104), .IN3(\in_a_r[2][3] ), 
        .IN4(n98), .Q(n17) );
  AO22X1 U18 ( .IN1(\in_a_r_reg[2][4] ), .IN2(n104), .IN3(\in_a_r[2][4] ), 
        .IN4(n98), .Q(n18) );
  AO22X1 U19 ( .IN1(\in_a_r_reg[2][5] ), .IN2(n105), .IN3(\in_a_r[2][5] ), 
        .IN4(n98), .Q(n19) );
  AO22X1 U20 ( .IN1(\in_a_r_reg[2][6] ), .IN2(n105), .IN3(\in_a_r[2][6] ), 
        .IN4(n98), .Q(n20) );
  AO22X1 U21 ( .IN1(\in_a_r_reg[2][7] ), .IN2(n105), .IN3(\in_a_r[2][7] ), 
        .IN4(n98), .Q(n21) );
  AO22X1 U22 ( .IN1(\in_a_r_reg[2][8] ), .IN2(n105), .IN3(\in_a_r[2][8] ), 
        .IN4(n98), .Q(n22) );
  AO22X1 U23 ( .IN1(\in_a_r_reg[2][9] ), .IN2(n105), .IN3(\in_a_r[2][9] ), 
        .IN4(n98), .Q(n23) );
  AO22X1 U24 ( .IN1(\in_a_r_reg[2][10] ), .IN2(n105), .IN3(\in_a_r[2][10] ), 
        .IN4(n98), .Q(n24) );
  AO22X1 U25 ( .IN1(\in_a_r_reg[2][11] ), .IN2(n105), .IN3(\in_a_r[2][11] ), 
        .IN4(n98), .Q(n25) );
  AO22X1 U27 ( .IN1(\in_a_r_reg[1][1] ), .IN2(n106), .IN3(\in_a_r[1][1] ), 
        .IN4(n98), .Q(n27) );
  AO22X1 U28 ( .IN1(\in_a_r_reg[1][2] ), .IN2(n106), .IN3(\in_a_r[1][2] ), 
        .IN4(n98), .Q(n28) );
  AO22X1 U29 ( .IN1(\in_a_r_reg[1][3] ), .IN2(n106), .IN3(\in_a_r[1][3] ), 
        .IN4(n98), .Q(n29) );
  AO22X1 U30 ( .IN1(\in_a_r_reg[1][4] ), .IN2(n106), .IN3(\in_a_r[1][4] ), 
        .IN4(n98), .Q(n30) );
  AO22X1 U31 ( .IN1(\in_a_r_reg[1][5] ), .IN2(n106), .IN3(\in_a_r[1][5] ), 
        .IN4(n98), .Q(n31) );
  AO22X1 U32 ( .IN1(\in_a_r_reg[1][6] ), .IN2(n106), .IN3(\in_a_r[1][6] ), 
        .IN4(n98), .Q(n32) );
  AO22X1 U33 ( .IN1(\in_a_r_reg[1][7] ), .IN2(n106), .IN3(\in_a_r[1][7] ), 
        .IN4(n99), .Q(n33) );
  AO22X1 U34 ( .IN1(\in_a_r_reg[1][8] ), .IN2(n107), .IN3(\in_a_r[1][8] ), 
        .IN4(n99), .Q(n34) );
  AO22X1 U35 ( .IN1(\in_a_r_reg[1][9] ), .IN2(n107), .IN3(\in_a_r[1][9] ), 
        .IN4(n99), .Q(n35) );
  AO22X1 U36 ( .IN1(\in_a_r_reg[1][10] ), .IN2(n107), .IN3(\in_a_r[1][10] ), 
        .IN4(n99), .Q(n36) );
  AO22X1 U37 ( .IN1(\in_a_r_reg[1][11] ), .IN2(n107), .IN3(\in_a_r[1][11] ), 
        .IN4(n99), .Q(n37) );
  AO22X1 U40 ( .IN1(\in_a_r_reg[0][2] ), .IN2(n107), .IN3(\in_a_r[0][2] ), 
        .IN4(n99), .Q(n40) );
  AO22X1 U41 ( .IN1(\in_a_r_reg[0][3] ), .IN2(n107), .IN3(\in_a_r[0][3] ), 
        .IN4(n99), .Q(n41) );
  AO22X1 U42 ( .IN1(\in_a_r_reg[0][4] ), .IN2(n107), .IN3(\in_a_r[0][4] ), 
        .IN4(n99), .Q(n42) );
  AO22X1 U43 ( .IN1(\in_a_r_reg[0][5] ), .IN2(n108), .IN3(\in_a_r[0][5] ), 
        .IN4(n99), .Q(n43) );
  AO22X1 U44 ( .IN1(\in_a_r_reg[0][6] ), .IN2(n108), .IN3(\in_a_r[0][6] ), 
        .IN4(n99), .Q(n44) );
  AO22X1 U45 ( .IN1(\in_a_r_reg[0][7] ), .IN2(n108), .IN3(\in_a_r[0][7] ), 
        .IN4(n99), .Q(n45) );
  AO22X1 U46 ( .IN1(\in_a_r_reg[0][8] ), .IN2(n108), .IN3(\in_a_r[0][8] ), 
        .IN4(n99), .Q(n46) );
  AO22X1 U47 ( .IN1(\in_a_r_reg[0][9] ), .IN2(n108), .IN3(\in_a_r[0][9] ), 
        .IN4(n99), .Q(n47) );
  AO22X1 U48 ( .IN1(\in_a_r_reg[0][10] ), .IN2(n108), .IN3(\in_a_r[0][10] ), 
        .IN4(n99), .Q(n48) );
  AO22X1 U49 ( .IN1(\in_a_r_reg[0][11] ), .IN2(n108), .IN3(\in_a_r[0][11] ), 
        .IN4(n99), .Q(n49) );
  AO22X1 U51 ( .IN1(\in_a_i_reg[3][1] ), .IN2(n109), .IN3(\in_a_i[3][1] ), 
        .IN4(n99), .Q(n51) );
  AO22X1 U52 ( .IN1(\in_a_i_reg[3][2] ), .IN2(n109), .IN3(\in_a_i[3][2] ), 
        .IN4(n99), .Q(n52) );
  AO22X1 U53 ( .IN1(\in_a_i_reg[3][3] ), .IN2(n109), .IN3(\in_a_i[3][3] ), 
        .IN4(n99), .Q(n53) );
  AO22X1 U54 ( .IN1(\in_a_i_reg[3][4] ), .IN2(n109), .IN3(\in_a_i[3][4] ), 
        .IN4(n99), .Q(n54) );
  AO22X1 U55 ( .IN1(\in_a_i_reg[3][5] ), .IN2(n109), .IN3(\in_a_i[3][5] ), 
        .IN4(n99), .Q(n55) );
  AO22X1 U56 ( .IN1(\in_a_i_reg[3][6] ), .IN2(n109), .IN3(\in_a_i[3][6] ), 
        .IN4(n99), .Q(n56) );
  AO22X1 U57 ( .IN1(\in_a_i_reg[3][7] ), .IN2(n109), .IN3(\in_a_i[3][7] ), 
        .IN4(n99), .Q(n57) );
  AO22X1 U58 ( .IN1(\in_a_i_reg[3][8] ), .IN2(n110), .IN3(\in_a_i[3][8] ), 
        .IN4(n99), .Q(n58) );
  AO22X1 U59 ( .IN1(\in_a_i_reg[3][9] ), .IN2(n110), .IN3(\in_a_i[3][9] ), 
        .IN4(n99), .Q(n59) );
  AO22X1 U60 ( .IN1(\in_a_i_reg[3][10] ), .IN2(n110), .IN3(\in_a_i[3][10] ), 
        .IN4(n100), .Q(n60) );
  AO22X1 U61 ( .IN1(\in_a_i_reg[3][11] ), .IN2(n110), .IN3(\in_a_i[3][11] ), 
        .IN4(n100), .Q(n61) );
  AO22X1 U63 ( .IN1(\in_a_i_reg[2][1] ), .IN2(n110), .IN3(\in_a_i[2][1] ), 
        .IN4(n100), .Q(n63) );
  AO22X1 U64 ( .IN1(\in_a_i_reg[2][2] ), .IN2(n110), .IN3(\in_a_i[2][2] ), 
        .IN4(n100), .Q(n64) );
  AO22X1 U65 ( .IN1(\in_a_i_reg[2][3] ), .IN2(n110), .IN3(\in_a_i[2][3] ), 
        .IN4(n100), .Q(n65) );
  AO22X1 U66 ( .IN1(\in_a_i_reg[2][4] ), .IN2(n111), .IN3(\in_a_i[2][4] ), 
        .IN4(n100), .Q(n66) );
  AO22X1 U67 ( .IN1(\in_a_i_reg[2][5] ), .IN2(n111), .IN3(\in_a_i[2][5] ), 
        .IN4(n100), .Q(n67) );
  AO22X1 U68 ( .IN1(\in_a_i_reg[2][6] ), .IN2(n111), .IN3(\in_a_i[2][6] ), 
        .IN4(n100), .Q(n68) );
  AO22X1 U69 ( .IN1(\in_a_i_reg[2][7] ), .IN2(n111), .IN3(\in_a_i[2][7] ), 
        .IN4(n100), .Q(n69) );
  AO22X1 U70 ( .IN1(\in_a_i_reg[2][8] ), .IN2(n111), .IN3(\in_a_i[2][8] ), 
        .IN4(n100), .Q(n70) );
  AO22X1 U71 ( .IN1(\in_a_i_reg[2][9] ), .IN2(n111), .IN3(\in_a_i[2][9] ), 
        .IN4(n100), .Q(n71) );
  AO22X1 U72 ( .IN1(\in_a_i_reg[2][10] ), .IN2(n111), .IN3(\in_a_i[2][10] ), 
        .IN4(n100), .Q(n72) );
  AO22X1 U73 ( .IN1(\in_a_i_reg[2][11] ), .IN2(n112), .IN3(\in_a_i[2][11] ), 
        .IN4(n100), .Q(n73) );
  AO22X1 U75 ( .IN1(\in_a_i_reg[1][1] ), .IN2(n112), .IN3(\in_a_i[1][1] ), 
        .IN4(n100), .Q(n75) );
  AO22X1 U76 ( .IN1(\in_a_i_reg[1][2] ), .IN2(n112), .IN3(\in_a_i[1][2] ), 
        .IN4(n100), .Q(n76) );
  AO22X1 U77 ( .IN1(\in_a_i_reg[1][3] ), .IN2(n112), .IN3(\in_a_i[1][3] ), 
        .IN4(n100), .Q(n77) );
  AO22X1 U78 ( .IN1(\in_a_i_reg[1][4] ), .IN2(n112), .IN3(\in_a_i[1][4] ), 
        .IN4(n100), .Q(n78) );
  AO22X1 U79 ( .IN1(\in_a_i_reg[1][5] ), .IN2(n112), .IN3(\in_a_i[1][5] ), 
        .IN4(n100), .Q(n79) );
  AO22X1 U80 ( .IN1(\in_a_i_reg[1][6] ), .IN2(n112), .IN3(\in_a_i[1][6] ), 
        .IN4(n100), .Q(n80) );
  AO22X1 U81 ( .IN1(\in_a_i_reg[1][7] ), .IN2(n113), .IN3(\in_a_i[1][7] ), 
        .IN4(n100), .Q(n81) );
  AO22X1 U82 ( .IN1(\in_a_i_reg[1][8] ), .IN2(n113), .IN3(\in_a_i[1][8] ), 
        .IN4(n100), .Q(n82) );
  AO22X1 U83 ( .IN1(\in_a_i_reg[1][9] ), .IN2(n113), .IN3(\in_a_i[1][9] ), 
        .IN4(n100), .Q(n83) );
  AO22X1 U84 ( .IN1(\in_a_i_reg[1][10] ), .IN2(n113), .IN3(\in_a_i[1][10] ), 
        .IN4(n100), .Q(n84) );
  AO22X1 U85 ( .IN1(\in_a_i_reg[1][11] ), .IN2(n113), .IN3(\in_a_i[1][11] ), 
        .IN4(n100), .Q(n85) );
  AO22X1 U88 ( .IN1(\in_a_i_reg[0][2] ), .IN2(n113), .IN3(\in_a_i[0][2] ), 
        .IN4(n101), .Q(n88) );
  AO22X1 U89 ( .IN1(\in_a_i_reg[0][3] ), .IN2(n113), .IN3(\in_a_i[0][3] ), 
        .IN4(n101), .Q(n89) );
  AO22X1 U90 ( .IN1(\in_a_i_reg[0][4] ), .IN2(n114), .IN3(\in_a_i[0][4] ), 
        .IN4(n101), .Q(n90) );
  AO22X1 U91 ( .IN1(\in_a_i_reg[0][5] ), .IN2(n114), .IN3(\in_a_i[0][5] ), 
        .IN4(n101), .Q(n91) );
  AO22X1 U92 ( .IN1(\in_a_i_reg[0][6] ), .IN2(n114), .IN3(\in_a_i[0][6] ), 
        .IN4(n101), .Q(n92) );
  AO22X1 U93 ( .IN1(\in_a_i_reg[0][7] ), .IN2(n114), .IN3(\in_a_i[0][7] ), 
        .IN4(n101), .Q(n93) );
  AO22X1 U94 ( .IN1(\in_a_i_reg[0][8] ), .IN2(n114), .IN3(\in_a_i[0][8] ), 
        .IN4(n101), .Q(n94) );
  AO22X1 U95 ( .IN1(\in_a_i_reg[0][9] ), .IN2(n114), .IN3(\in_a_i[0][9] ), 
        .IN4(n101), .Q(n95) );
  AO22X1 U96 ( .IN1(\in_a_i_reg[0][10] ), .IN2(n114), .IN3(\in_a_i[0][10] ), 
        .IN4(n101), .Q(n96) );
  AO22X1 U97 ( .IN1(\in_a_i_reg[0][11] ), .IN2(n114), .IN3(\in_a_i[0][11] ), 
        .IN4(n101), .Q(n97) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_7 sub_r_0 ( .a({\in_a_r_reg[0][11] , 
        \in_a_r_reg[0][10] , \in_a_r_reg[0][9] , \in_a_r_reg[0][8] , 
        \in_a_r_reg[0][7] , \in_a_r_reg[0][6] , \in_a_r_reg[0][5] , 
        \in_a_r_reg[0][4] , \in_a_r_reg[0][3] , \in_a_r_reg[0][2] , 
        \in_a_r_reg[0][1] , \in_a_r_reg[0][0] }), .b({\in_b_r[0][11] , 
        \in_b_r[0][10] , \in_b_r[0][9] , \in_b_r[0][8] , \in_b_r[0][7] , 
        \in_b_r[0][6] , \in_b_r[0][5] , \in_b_r[0][4] , \in_b_r[0][3] , 
        \in_b_r[0][2] , \in_b_r[0][1] , \in_b_r[0][0] }), .\output ({
        \out_r[0][11] , \out_r[0][10] , \out_r[0][9] , \out_r[0][8] , 
        \out_r[0][7] , \out_r[0][6] , \out_r[0][5] , \out_r[0][4] , 
        \out_r[0][3] , \out_r[0][2] , \out_r[0][1] , \out_r[0][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_6 sub_i_0 ( .a({\in_a_i_reg[0][11] , 
        \in_a_i_reg[0][10] , \in_a_i_reg[0][9] , \in_a_i_reg[0][8] , 
        \in_a_i_reg[0][7] , \in_a_i_reg[0][6] , \in_a_i_reg[0][5] , 
        \in_a_i_reg[0][4] , \in_a_i_reg[0][3] , \in_a_i_reg[0][2] , 
        \in_a_i_reg[0][1] , \in_a_i_reg[0][0] }), .b({\in_b_i[0][11] , 
        \in_b_i[0][10] , \in_b_i[0][9] , \in_b_i[0][8] , \in_b_i[0][7] , 
        \in_b_i[0][6] , \in_b_i[0][5] , \in_b_i[0][4] , \in_b_i[0][3] , 
        \in_b_i[0][2] , \in_b_i[0][1] , \in_b_i[0][0] }), .\output ({
        \out_i[0][11] , \out_i[0][10] , \out_i[0][9] , \out_i[0][8] , 
        \out_i[0][7] , \out_i[0][6] , \out_i[0][5] , \out_i[0][4] , 
        \out_i[0][3] , \out_i[0][2] , \out_i[0][1] , \out_i[0][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_5 sub_r_1 ( .a({\in_a_r_reg[1][11] , 
        \in_a_r_reg[1][10] , \in_a_r_reg[1][9] , \in_a_r_reg[1][8] , 
        \in_a_r_reg[1][7] , \in_a_r_reg[1][6] , \in_a_r_reg[1][5] , 
        \in_a_r_reg[1][4] , \in_a_r_reg[1][3] , \in_a_r_reg[1][2] , 
        \in_a_r_reg[1][1] , \in_a_r_reg[1][0] }), .b({\in_b_r[1][11] , 
        \in_b_r[1][10] , \in_b_r[1][9] , \in_b_r[1][8] , \in_b_r[1][7] , 
        \in_b_r[1][6] , \in_b_r[1][5] , \in_b_r[1][4] , \in_b_r[1][3] , 
        \in_b_r[1][2] , \in_b_r[1][1] , \in_b_r[1][0] }), .\output ({
        \out_r[1][11] , \out_r[1][10] , \out_r[1][9] , \out_r[1][8] , 
        \out_r[1][7] , \out_r[1][6] , \out_r[1][5] , \out_r[1][4] , 
        \out_r[1][3] , \out_r[1][2] , \out_r[1][1] , \out_r[1][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_4 sub_i_1 ( .a({\in_a_i_reg[1][11] , 
        \in_a_i_reg[1][10] , \in_a_i_reg[1][9] , \in_a_i_reg[1][8] , 
        \in_a_i_reg[1][7] , \in_a_i_reg[1][6] , \in_a_i_reg[1][5] , 
        \in_a_i_reg[1][4] , \in_a_i_reg[1][3] , \in_a_i_reg[1][2] , 
        \in_a_i_reg[1][1] , \in_a_i_reg[1][0] }), .b({\in_b_i[1][11] , 
        \in_b_i[1][10] , \in_b_i[1][9] , \in_b_i[1][8] , \in_b_i[1][7] , 
        \in_b_i[1][6] , \in_b_i[1][5] , \in_b_i[1][4] , \in_b_i[1][3] , 
        \in_b_i[1][2] , \in_b_i[1][1] , \in_b_i[1][0] }), .\output ({
        \out_i[1][11] , \out_i[1][10] , \out_i[1][9] , \out_i[1][8] , 
        \out_i[1][7] , \out_i[1][6] , \out_i[1][5] , \out_i[1][4] , 
        \out_i[1][3] , \out_i[1][2] , \out_i[1][1] , \out_i[1][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_3 sub_r_2 ( .a({\in_a_r_reg[2][11] , 
        \in_a_r_reg[2][10] , \in_a_r_reg[2][9] , \in_a_r_reg[2][8] , 
        \in_a_r_reg[2][7] , \in_a_r_reg[2][6] , \in_a_r_reg[2][5] , 
        \in_a_r_reg[2][4] , \in_a_r_reg[2][3] , \in_a_r_reg[2][2] , 
        \in_a_r_reg[2][1] , \in_a_r_reg[2][0] }), .b({\in_b_r[2][11] , 
        \in_b_r[2][10] , \in_b_r[2][9] , \in_b_r[2][8] , \in_b_r[2][7] , 
        \in_b_r[2][6] , \in_b_r[2][5] , \in_b_r[2][4] , \in_b_r[2][3] , 
        \in_b_r[2][2] , \in_b_r[2][1] , \in_b_r[2][0] }), .\output ({
        \out_r[2][11] , \out_r[2][10] , \out_r[2][9] , \out_r[2][8] , 
        \out_r[2][7] , \out_r[2][6] , \out_r[2][5] , \out_r[2][4] , 
        \out_r[2][3] , \out_r[2][2] , \out_r[2][1] , \out_r[2][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_2 sub_i_2 ( .a({\in_a_i_reg[2][11] , 
        \in_a_i_reg[2][10] , \in_a_i_reg[2][9] , \in_a_i_reg[2][8] , 
        \in_a_i_reg[2][7] , \in_a_i_reg[2][6] , \in_a_i_reg[2][5] , 
        \in_a_i_reg[2][4] , \in_a_i_reg[2][3] , \in_a_i_reg[2][2] , 
        \in_a_i_reg[2][1] , \in_a_i_reg[2][0] }), .b({\in_b_i[2][11] , 
        \in_b_i[2][10] , \in_b_i[2][9] , \in_b_i[2][8] , \in_b_i[2][7] , 
        \in_b_i[2][6] , \in_b_i[2][5] , \in_b_i[2][4] , \in_b_i[2][3] , 
        \in_b_i[2][2] , \in_b_i[2][1] , \in_b_i[2][0] }), .\output ({
        \out_i[2][11] , \out_i[2][10] , \out_i[2][9] , \out_i[2][8] , 
        \out_i[2][7] , \out_i[2][6] , \out_i[2][5] , \out_i[2][4] , 
        \out_i[2][3] , \out_i[2][2] , \out_i[2][1] , \out_i[2][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_1 sub_r_3 ( .a({\in_a_r_reg[3][11] , 
        \in_a_r_reg[3][10] , \in_a_r_reg[3][9] , \in_a_r_reg[3][8] , 
        \in_a_r_reg[3][7] , \in_a_r_reg[3][6] , \in_a_r_reg[3][5] , 
        \in_a_r_reg[3][4] , \in_a_r_reg[3][3] , \in_a_r_reg[3][2] , 
        \in_a_r_reg[3][1] , \in_a_r_reg[3][0] }), .b({\in_b_r[3][11] , 
        \in_b_r[3][10] , \in_b_r[3][9] , \in_b_r[3][8] , \in_b_r[3][7] , 
        \in_b_r[3][6] , \in_b_r[3][5] , \in_b_r[3][4] , \in_b_r[3][3] , 
        \in_b_r[3][2] , \in_b_r[3][1] , \in_b_r[3][0] }), .\output ({
        \out_r[3][11] , \out_r[3][10] , \out_r[3][9] , \out_r[3][8] , 
        \out_r[3][7] , \out_r[3][6] , \out_r[3][5] , \out_r[3][4] , 
        \out_r[3][3] , \out_r[3][2] , \out_r[3][1] , \out_r[3][0] }) );
  add_sub_WORD_WIDTH12_OPERATION0_USE_SAT1_0 sub_i_3 ( .a({\in_a_i_reg[3][11] , 
        \in_a_i_reg[3][10] , \in_a_i_reg[3][9] , \in_a_i_reg[3][8] , 
        \in_a_i_reg[3][7] , \in_a_i_reg[3][6] , \in_a_i_reg[3][5] , 
        \in_a_i_reg[3][4] , \in_a_i_reg[3][3] , \in_a_i_reg[3][2] , 
        \in_a_i_reg[3][1] , \in_a_i_reg[3][0] }), .b({\in_b_i[3][11] , 
        \in_b_i[3][10] , \in_b_i[3][9] , \in_b_i[3][8] , \in_b_i[3][7] , 
        \in_b_i[3][6] , \in_b_i[3][5] , \in_b_i[3][4] , \in_b_i[3][3] , 
        \in_b_i[3][2] , \in_b_i[3][1] , \in_b_i[3][0] }), .\output ({
        \out_i[3][11] , \out_i[3][10] , \out_i[3][9] , \out_i[3][8] , 
        \out_i[3][7] , \out_i[3][6] , \out_i[3][5] , \out_i[3][4] , 
        \out_i[3][3] , \out_i[3][2] , \out_i[3][1] , \out_i[3][0] }) );
  INVX0 U2 ( .INP(n102), .ZN(n99) );
  INVX0 U14 ( .INP(n102), .ZN(n100) );
  INVX0 U26 ( .INP(n102), .ZN(n1) );
  NBUFFX2 U38 ( .INP(n115), .Z(n102) );
  NBUFFX2 U39 ( .INP(n107), .Z(n104) );
  NBUFFX2 U50 ( .INP(n108), .Z(n105) );
  NBUFFX2 U62 ( .INP(n110), .Z(n106) );
  NBUFFX2 U74 ( .INP(n115), .Z(n107) );
  NBUFFX2 U86 ( .INP(n115), .Z(n108) );
  NBUFFX2 U87 ( .INP(n111), .Z(n109) );
  NBUFFX2 U98 ( .INP(n115), .Z(n110) );
  NBUFFX2 U99 ( .INP(n115), .Z(n111) );
  NBUFFX2 U100 ( .INP(n115), .Z(n112) );
  NBUFFX2 U101 ( .INP(n115), .Z(n113) );
  NBUFFX2 U102 ( .INP(n115), .Z(n114) );
  NBUFFX2 U103 ( .INP(n113), .Z(n103) );
  INVX0 U104 ( .INP(n102), .ZN(n98) );
  INVX0 U105 ( .INP(n102), .ZN(n101) );
  INVX0 U106 ( .INP(w_in_a), .ZN(n115) );
  MUX21X1 U107 ( .IN1(\in_a_i_reg[3][0] ), .IN2(\in_a_i[3][0] ), .S(n1), .Q(
        n50) );
  MUX21X1 U108 ( .IN1(\in_a_r_reg[3][0] ), .IN2(\in_a_r[3][0] ), .S(n1), .Q(n2) );
  MUX21X1 U109 ( .IN1(\in_a_i_reg[2][0] ), .IN2(\in_a_i[2][0] ), .S(n1), .Q(
        n62) );
  MUX21X1 U110 ( .IN1(\in_a_r_reg[2][0] ), .IN2(\in_a_r[2][0] ), .S(n1), .Q(
        n14) );
  MUX21X1 U111 ( .IN1(\in_a_i_reg[1][0] ), .IN2(\in_a_i[1][0] ), .S(n1), .Q(
        n74) );
  MUX21X1 U112 ( .IN1(\in_a_r_reg[1][0] ), .IN2(\in_a_r[1][0] ), .S(n1), .Q(
        n26) );
  MUX21X1 U113 ( .IN1(\in_a_i_reg[0][0] ), .IN2(\in_a_i[0][0] ), .S(n1), .Q(
        n86) );
  MUX21X1 U114 ( .IN1(\in_a_i_reg[0][1] ), .IN2(\in_a_i[0][1] ), .S(n1), .Q(
        n87) );
  MUX21X1 U115 ( .IN1(\in_a_r_reg[0][0] ), .IN2(\in_a_r[0][0] ), .S(n1), .Q(
        n38) );
  MUX21X1 U116 ( .IN1(\in_a_r_reg[0][1] ), .IN2(\in_a_r[0][1] ), .S(n1), .Q(
        n39) );
endmodule


module mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_DW01_inc_0 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;

  wire   [12:2] carry;

  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  XOR2X1 U1 ( .IN1(carry[12]), .IN2(A[12]), .Q(SUM[12]) );
endmodule


module mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_DW_mult_tc_0 ( a, b, 
        product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n25, n27, n28, n29, n30, n31, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n146, n147, n148, n149, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n202, n203, n204, n205, n206, n207, n208, n209, n210, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534;

  FADDX1 U4 ( .A(n25), .B(n152), .CI(n4), .CO(n3), .S(product[22]) );
  FADDX1 U5 ( .A(n27), .B(n430), .CI(n5), .CO(n4), .S(product[21]) );
  FADDX1 U6 ( .A(n29), .B(n28), .CI(n6), .CO(n5), .S(product[20]) );
  FADDX1 U7 ( .A(n33), .B(n30), .CI(n7), .CO(n6), .S(product[19]) );
  FADDX1 U8 ( .A(n37), .B(n34), .CI(n8), .CO(n7), .S(product[18]) );
  FADDX1 U9 ( .A(n43), .B(n38), .CI(n9), .CO(n8), .S(product[17]) );
  FADDX1 U10 ( .A(n49), .B(n44), .CI(n10), .CO(n9), .S(product[16]) );
  FADDX1 U11 ( .A(n57), .B(n50), .CI(n11), .CO(n10), .S(product[15]) );
  FADDX1 U12 ( .A(n65), .B(n58), .CI(n12), .CO(n11), .S(product[14]) );
  FADDX1 U13 ( .A(n66), .B(n75), .CI(n13), .CO(n12), .S(product[13]) );
  FADDX1 U14 ( .A(n76), .B(n85), .CI(n14), .CO(n13), .S(product[12]) );
  FADDX1 U15 ( .A(n86), .B(n95), .CI(n15), .CO(n14), .S(product[11]) );
  FADDX1 U17 ( .A(n104), .B(n111), .CI(n17), .CO(n16), .S(product[9]) );
  FADDX1 U27 ( .A(n153), .B(n164), .CI(n31), .CO(n27), .S(n28) );
  FADDX1 U28 ( .A(n428), .B(n154), .CI(n35), .CO(n29), .S(n30) );
  FADDX1 U30 ( .A(n36), .B(n41), .CI(n39), .CO(n33), .S(n34) );
  FADDX1 U31 ( .A(n165), .B(n176), .CI(n155), .CO(n35), .S(n36) );
  FADDX1 U32 ( .A(n40), .B(n47), .CI(n45), .CO(n37), .S(n38) );
  FADDX1 U33 ( .A(n156), .B(n166), .CI(n426), .CO(n39), .S(n40) );
  FADDX1 U35 ( .A(n46), .B(n48), .CI(n51), .CO(n43), .S(n44) );
  FADDX1 U36 ( .A(n55), .B(n167), .CI(n53), .CO(n45), .S(n46) );
  FADDX1 U37 ( .A(n157), .B(n188), .CI(n177), .CO(n47), .S(n48) );
  FADDX1 U38 ( .A(n52), .B(n54), .CI(n59), .CO(n49), .S(n50) );
  FADDX1 U39 ( .A(n63), .B(n424), .CI(n61), .CO(n51), .S(n52) );
  FADDX1 U40 ( .A(n158), .B(n168), .CI(n178), .CO(n53), .S(n54) );
  FADDX1 U42 ( .A(n60), .B(n69), .CI(n67), .CO(n57), .S(n58) );
  FADDX1 U43 ( .A(n64), .B(n71), .CI(n62), .CO(n59), .S(n60) );
  FADDX1 U44 ( .A(n169), .B(n73), .CI(n179), .CO(n61), .S(n62) );
  FADDX1 U45 ( .A(n159), .B(n200), .CI(n189), .CO(n63), .S(n64) );
  FADDX1 U46 ( .A(n77), .B(n79), .CI(n68), .CO(n65), .S(n66) );
  FADDX1 U47 ( .A(n72), .B(n81), .CI(n70), .CO(n67), .S(n68) );
  FADDX1 U48 ( .A(n421), .B(n180), .CI(n83), .CO(n69), .S(n70) );
  FADDX1 U49 ( .A(n190), .B(n170), .CI(n160), .CO(n71), .S(n72) );
  FADDX1 U51 ( .A(n87), .B(n80), .CI(n78), .CO(n75), .S(n76) );
  FADDX1 U52 ( .A(n82), .B(n84), .CI(n89), .CO(n77), .S(n78) );
  FADDX1 U53 ( .A(n93), .B(n181), .CI(n91), .CO(n79), .S(n80) );
  FADDX1 U54 ( .A(n161), .B(n191), .CI(n171), .CO(n81), .S(n82) );
  FADDX1 U57 ( .A(n97), .B(n90), .CI(n88), .CO(n85), .S(n86) );
  FADDX1 U58 ( .A(n99), .B(n101), .CI(n92), .CO(n87), .S(n88) );
  FADDX1 U59 ( .A(n172), .B(n192), .CI(n94), .CO(n89), .S(n90) );
  FADDX1 U60 ( .A(n182), .B(n146), .CI(n202), .CO(n91), .S(n92) );
  HADDX1 U61 ( .A0(n213), .B0(n162), .C1(n93), .SO(n94) );
  FADDX1 U62 ( .A(n105), .B(n100), .CI(n98), .CO(n95), .S(n96) );
  FADDX1 U63 ( .A(n102), .B(n109), .CI(n107), .CO(n97), .S(n98) );
  FADDX1 U64 ( .A(n183), .B(n173), .CI(n193), .CO(n99), .S(n100) );
  FADDX1 U65 ( .A(n214), .B(n163), .CI(n203), .CO(n101), .S(n102) );
  FADDX1 U66 ( .A(n113), .B(n108), .CI(n106), .CO(n103), .S(n104) );
  FADDX1 U67 ( .A(n110), .B(n204), .CI(n115), .CO(n105), .S(n106) );
  FADDX1 U68 ( .A(n147), .B(n184), .CI(n194), .CO(n107), .S(n108) );
  HADDX1 U69 ( .A0(n215), .B0(n174), .C1(n109), .SO(n110) );
  FADDX1 U70 ( .A(n116), .B(n119), .CI(n114), .CO(n111), .S(n112) );
  FADDX1 U71 ( .A(n185), .B(n195), .CI(n121), .CO(n113), .S(n114) );
  FADDX1 U72 ( .A(n216), .B(n175), .CI(n205), .CO(n115), .S(n116) );
  FADDX1 U73 ( .A(n125), .B(n122), .CI(n120), .CO(n117), .S(n118) );
  FADDX1 U74 ( .A(n148), .B(n206), .CI(n196), .CO(n119), .S(n120) );
  HADDX1 U75 ( .A0(n217), .B0(n186), .C1(n121), .SO(n122) );
  FADDX1 U76 ( .A(n129), .B(n197), .CI(n126), .CO(n123), .S(n124) );
  FADDX1 U77 ( .A(n207), .B(n187), .CI(n218), .CO(n125), .S(n126) );
  FADDX1 U78 ( .A(n149), .B(n198), .CI(n130), .CO(n127), .S(n128) );
  HADDX1 U79 ( .A0(n219), .B0(n208), .C1(n129), .SO(n130) );
  FADDX1 U80 ( .A(n220), .B(n199), .CI(n209), .CO(n131), .S(n132) );
  HADDX1 U81 ( .A0(n221), .B0(n210), .C1(n133), .SO(n134) );
  INVX0 U309 ( .INP(b[9]), .ZN(n400) );
  INVX0 U310 ( .INP(n400), .ZN(n401) );
  INVX0 U311 ( .INP(b[1]), .ZN(n402) );
  INVX0 U312 ( .INP(n402), .ZN(n403) );
  DELLN1X2 U313 ( .INP(b[6]), .Z(n404) );
  INVX0 U314 ( .INP(b[3]), .ZN(n405) );
  INVX0 U315 ( .INP(n405), .ZN(n406) );
  FADDX1 U316 ( .A(n118), .B(n123), .CI(n19), .CO(n18), .S(product[7]) );
  FADDX1 U317 ( .A(n112), .B(n117), .CI(n18), .CO(n17), .S(product[8]) );
  FADDX1 U318 ( .A(n96), .B(n103), .CI(n16), .CO(n15), .S(product[10]) );
  INVX0 U319 ( .INP(b[8]), .ZN(n407) );
  INVX0 U320 ( .INP(n407), .ZN(n408) );
  DELLN1X2 U321 ( .INP(b[5]), .Z(n409) );
  XOR2X2 U322 ( .IN1(b[6]), .IN2(a[1]), .Q(n459) );
  DELLN1X2 U323 ( .INP(b[4]), .Z(n410) );
  DELLN1X2 U324 ( .INP(b[2]), .Z(n411) );
  XOR2X2 U325 ( .IN1(n409), .IN2(n415), .Q(n469) );
  XOR2X2 U326 ( .IN1(b[5]), .IN2(a[1]), .Q(n458) );
  INVX0 U327 ( .INP(a[11]), .ZN(n412) );
  INVX1 U328 ( .INP(n412), .ZN(n413) );
  AND2X2 U329 ( .IN1(n516), .IN2(n534), .Q(n453) );
  XOR2X2 U330 ( .IN1(a[11]), .IN2(a[10]), .Q(n534) );
  AND2X2 U331 ( .IN1(n422), .IN2(n490), .Q(n438) );
  XOR2X2 U332 ( .IN1(n408), .IN2(n418), .Q(n514) );
  XOR2X2 U333 ( .IN1(n408), .IN2(n417), .Q(n503) );
  XOR2X2 U334 ( .IN1(n408), .IN2(n416), .Q(n482) );
  XOR2X2 U335 ( .IN1(n408), .IN2(n415), .Q(n472) );
  XOR2X2 U336 ( .IN1(n410), .IN2(n413), .Q(n521) );
  XOR2X2 U337 ( .IN1(n410), .IN2(n418), .Q(n510) );
  XOR2X2 U338 ( .IN1(n410), .IN2(n417), .Q(n499) );
  XOR2X2 U339 ( .IN1(n410), .IN2(n416), .Q(n478) );
  XOR2X2 U340 ( .IN1(n410), .IN2(n415), .Q(n468) );
  XOR2X2 U341 ( .IN1(b[4]), .IN2(a[1]), .Q(n457) );
  XOR2X2 U342 ( .IN1(n406), .IN2(a[1]), .Q(n455) );
  XOR2X2 U343 ( .IN1(n406), .IN2(n415), .Q(n467) );
  XOR2X2 U344 ( .IN1(n406), .IN2(n416), .Q(n477) );
  XOR2X2 U345 ( .IN1(n406), .IN2(n417), .Q(n498) );
  XOR2X2 U346 ( .IN1(n406), .IN2(n418), .Q(n509) );
  XOR2X2 U347 ( .IN1(n406), .IN2(n413), .Q(n520) );
  XOR2X2 U348 ( .IN1(n411), .IN2(n413), .Q(n519) );
  XOR2X2 U349 ( .IN1(n411), .IN2(n418), .Q(n508) );
  XOR2X2 U350 ( .IN1(n411), .IN2(n417), .Q(n497) );
  XOR2X2 U351 ( .IN1(n411), .IN2(n416), .Q(n476) );
  XOR2X2 U352 ( .IN1(n411), .IN2(n415), .Q(n466) );
  XOR2X2 U353 ( .IN1(b[2]), .IN2(a[1]), .Q(n456) );
  XOR2X2 U354 ( .IN1(n403), .IN2(n413), .Q(n517) );
  XOR2X2 U355 ( .IN1(n403), .IN2(n418), .Q(n506) );
  XOR2X2 U356 ( .IN1(n403), .IN2(n417), .Q(n495) );
  XOR2X2 U357 ( .IN1(n403), .IN2(n416), .Q(n474) );
  XOR2X2 U358 ( .IN1(n403), .IN2(n415), .Q(n464) );
  INVX0 U359 ( .INP(n25), .ZN(n430) );
  INVX0 U360 ( .INP(n3), .ZN(product[23]) );
  INVX0 U361 ( .INP(n55), .ZN(n424) );
  INVX0 U362 ( .INP(n473), .ZN(n425) );
  INVX0 U363 ( .INP(n494), .ZN(n427) );
  INVX0 U364 ( .INP(n134), .ZN(n420) );
  INVX0 U365 ( .INP(n505), .ZN(n429) );
  INVX0 U366 ( .INP(n516), .ZN(n431) );
  INVX0 U367 ( .INP(n73), .ZN(n421) );
  INVX0 U368 ( .INP(n437), .ZN(n422) );
  INVX0 U369 ( .INP(n31), .ZN(n428) );
  INVX0 U370 ( .INP(n41), .ZN(n426) );
  INVX0 U371 ( .INP(n414), .ZN(n432) );
  DELLN1X2 U372 ( .INP(a[7]), .Z(n417) );
  DELLN1X2 U373 ( .INP(a[5]), .Z(n416) );
  DELLN1X2 U374 ( .INP(a[3]), .Z(n415) );
  AND2X1 U375 ( .IN1(n494), .IN2(n530), .Q(n447) );
  AND2X1 U376 ( .IN1(n473), .IN2(n528), .Q(n444) );
  DELLN1X2 U377 ( .INP(a[9]), .Z(n418) );
  AND2X1 U378 ( .IN1(n505), .IN2(n532), .Q(n450) );
  INVX0 U379 ( .INP(a[1]), .ZN(n423) );
  INVX0 U380 ( .INP(n403), .ZN(n433) );
  DELLN1X2 U381 ( .INP(b[0]), .Z(n414) );
  XNOR2X1 U382 ( .IN1(n434), .IN2(n435), .Q(n84) );
  NAND2X0 U383 ( .IN1(n435), .IN2(n434), .QN(n83) );
  AOI22X1 U384 ( .IN1(n436), .IN2(n437), .IN3(n438), .IN4(n439), .QN(n434) );
  OA21X1 U385 ( .IN1(n440), .IN2(a[0]), .IN3(n441), .Q(n435) );
  AO22X1 U386 ( .IN1(n442), .IN2(n437), .IN3(n438), .IN4(n436), .Q(n73) );
  XOR2X1 U387 ( .IN1(b[10]), .IN2(n415), .Q(n436) );
  AO22X1 U388 ( .IN1(n443), .IN2(n425), .IN3(n444), .IN4(n445), .Q(n55) );
  AO22X1 U389 ( .IN1(n446), .IN2(n427), .IN3(n447), .IN4(n448), .Q(n41) );
  AO22X1 U390 ( .IN1(n449), .IN2(n429), .IN3(n450), .IN4(n451), .Q(n31) );
  AO22X1 U391 ( .IN1(n452), .IN2(n431), .IN3(n453), .IN4(n454), .Q(n25) );
  AO22X1 U392 ( .IN1(a[0]), .IN2(n455), .IN3(n440), .IN4(n456), .Q(n221) );
  AO22X1 U393 ( .IN1(a[0]), .IN2(n457), .IN3(n440), .IN4(n455), .Q(n220) );
  AO22X1 U394 ( .IN1(a[0]), .IN2(n458), .IN3(n440), .IN4(n457), .Q(n219) );
  AO22X1 U395 ( .IN1(a[0]), .IN2(n459), .IN3(n440), .IN4(n458), .Q(n218) );
  AO22X1 U396 ( .IN1(a[0]), .IN2(n460), .IN3(n440), .IN4(n459), .Q(n217) );
  AO22X1 U397 ( .IN1(a[0]), .IN2(n461), .IN3(n440), .IN4(n460), .Q(n216) );
  XOR2X1 U398 ( .IN1(b[7]), .IN2(a[1]), .Q(n460) );
  AO22X1 U399 ( .IN1(a[0]), .IN2(n462), .IN3(n440), .IN4(n461), .Q(n215) );
  XOR2X1 U400 ( .IN1(n408), .IN2(a[1]), .Q(n461) );
  AO22X1 U401 ( .IN1(a[0]), .IN2(n463), .IN3(n440), .IN4(n462), .Q(n214) );
  XOR2X1 U402 ( .IN1(n401), .IN2(a[1]), .Q(n462) );
  AO22X1 U403 ( .IN1(a[0]), .IN2(n441), .IN3(n440), .IN4(n463), .Q(n213) );
  XOR2X1 U404 ( .IN1(b[10]), .IN2(a[1]), .Q(n463) );
  XNOR2X1 U405 ( .IN1(b[11]), .IN2(n423), .Q(n441) );
  AO22X1 U406 ( .IN1(n464), .IN2(n437), .IN3(n438), .IN4(n465), .Q(n210) );
  XOR2X1 U407 ( .IN1(n414), .IN2(n415), .Q(n465) );
  AO22X1 U408 ( .IN1(n466), .IN2(n437), .IN3(n438), .IN4(n464), .Q(n209) );
  AO22X1 U409 ( .IN1(n467), .IN2(n437), .IN3(n438), .IN4(n466), .Q(n208) );
  AO22X1 U410 ( .IN1(n468), .IN2(n437), .IN3(n438), .IN4(n467), .Q(n207) );
  AO22X1 U411 ( .IN1(n469), .IN2(n437), .IN3(n438), .IN4(n468), .Q(n206) );
  AO22X1 U412 ( .IN1(n470), .IN2(n437), .IN3(n438), .IN4(n469), .Q(n205) );
  AO22X1 U413 ( .IN1(n471), .IN2(n437), .IN3(n438), .IN4(n470), .Q(n204) );
  XOR2X1 U414 ( .IN1(n404), .IN2(n415), .Q(n470) );
  AO22X1 U415 ( .IN1(n472), .IN2(n437), .IN3(n438), .IN4(n471), .Q(n203) );
  XOR2X1 U416 ( .IN1(b[7]), .IN2(n415), .Q(n471) );
  AO22X1 U417 ( .IN1(n439), .IN2(n437), .IN3(n438), .IN4(n472), .Q(n202) );
  XOR2X1 U418 ( .IN1(n401), .IN2(n415), .Q(n439) );
  OAI21X1 U419 ( .IN1(n437), .IN2(n438), .IN3(n442), .QN(n200) );
  XOR2X1 U420 ( .IN1(b[11]), .IN2(n415), .Q(n442) );
  NOR2X0 U421 ( .IN1(n473), .IN2(n432), .QN(n199) );
  AO22X1 U422 ( .IN1(n474), .IN2(n425), .IN3(n444), .IN4(n475), .Q(n198) );
  XOR2X1 U423 ( .IN1(n414), .IN2(n416), .Q(n475) );
  AO22X1 U424 ( .IN1(n476), .IN2(n425), .IN3(n444), .IN4(n474), .Q(n197) );
  AO22X1 U425 ( .IN1(n477), .IN2(n425), .IN3(n444), .IN4(n476), .Q(n196) );
  AO22X1 U426 ( .IN1(n478), .IN2(n425), .IN3(n444), .IN4(n477), .Q(n195) );
  AO22X1 U427 ( .IN1(n479), .IN2(n425), .IN3(n444), .IN4(n478), .Q(n194) );
  AO22X1 U428 ( .IN1(n480), .IN2(n425), .IN3(n444), .IN4(n479), .Q(n193) );
  XOR2X1 U429 ( .IN1(n409), .IN2(n416), .Q(n479) );
  AO22X1 U430 ( .IN1(n481), .IN2(n425), .IN3(n444), .IN4(n480), .Q(n192) );
  XOR2X1 U431 ( .IN1(n404), .IN2(n416), .Q(n480) );
  AO22X1 U432 ( .IN1(n482), .IN2(n425), .IN3(n444), .IN4(n481), .Q(n191) );
  XOR2X1 U433 ( .IN1(b[7]), .IN2(n416), .Q(n481) );
  AO22X1 U434 ( .IN1(n483), .IN2(n425), .IN3(n444), .IN4(n482), .Q(n190) );
  AO222X1 U435 ( .IN1(n484), .IN2(n124), .IN3(n484), .IN4(n127), .IN5(n127), 
        .IN6(n124), .Q(n19) );
  AO222X1 U436 ( .IN1(n485), .IN2(n128), .IN3(n485), .IN4(n131), .IN5(n131), 
        .IN6(n128), .Q(n484) );
  AO222X1 U437 ( .IN1(n486), .IN2(n132), .IN3(n486), .IN4(n133), .IN5(n133), 
        .IN6(n132), .Q(n485) );
  OAI222X1 U438 ( .IN1(n487), .IN2(n420), .IN3(n488), .IN4(n487), .IN5(n488), 
        .IN6(n420), .QN(n486) );
  AOI22X1 U439 ( .IN1(n489), .IN2(n415), .IN3(n438), .IN4(n415), .QN(n488) );
  XOR2X1 U440 ( .IN1(n415), .IN2(a[2]), .Q(n490) );
  NOR2X0 U441 ( .IN1(n414), .IN2(n422), .QN(n489) );
  MUX21X1 U442 ( .IN1(n491), .IN2(n492), .S(n414), .Q(n487) );
  NAND2X0 U443 ( .IN1(n437), .IN2(n493), .QN(n492) );
  XOR2X1 U444 ( .IN1(a[2]), .IN2(a[1]), .Q(n437) );
  NAND3X0 U445 ( .IN1(n493), .IN2(n433), .IN3(a[1]), .QN(n491) );
  AO22X1 U446 ( .IN1(a[0]), .IN2(n456), .IN3(n440), .IN4(n433), .Q(n493) );
  NOR2X0 U447 ( .IN1(n423), .IN2(a[0]), .QN(n440) );
  AO22X1 U448 ( .IN1(n445), .IN2(n425), .IN3(n444), .IN4(n483), .Q(n189) );
  XOR2X1 U449 ( .IN1(n401), .IN2(n416), .Q(n483) );
  XOR2X1 U450 ( .IN1(b[10]), .IN2(n416), .Q(n445) );
  OAI21X1 U451 ( .IN1(n425), .IN2(n444), .IN3(n443), .QN(n188) );
  XOR2X1 U452 ( .IN1(b[11]), .IN2(n416), .Q(n443) );
  NOR2X0 U453 ( .IN1(n494), .IN2(n432), .QN(n187) );
  AO22X1 U454 ( .IN1(n495), .IN2(n427), .IN3(n447), .IN4(n496), .Q(n186) );
  XOR2X1 U455 ( .IN1(n414), .IN2(n417), .Q(n496) );
  AO22X1 U456 ( .IN1(n497), .IN2(n427), .IN3(n447), .IN4(n495), .Q(n185) );
  AO22X1 U457 ( .IN1(n498), .IN2(n427), .IN3(n447), .IN4(n497), .Q(n184) );
  AO22X1 U458 ( .IN1(n499), .IN2(n427), .IN3(n447), .IN4(n498), .Q(n183) );
  AO22X1 U459 ( .IN1(n500), .IN2(n427), .IN3(n447), .IN4(n499), .Q(n182) );
  AO22X1 U460 ( .IN1(n501), .IN2(n427), .IN3(n447), .IN4(n500), .Q(n181) );
  XOR2X1 U461 ( .IN1(n409), .IN2(n417), .Q(n500) );
  AO22X1 U462 ( .IN1(n502), .IN2(n427), .IN3(n447), .IN4(n501), .Q(n180) );
  XOR2X1 U463 ( .IN1(n404), .IN2(n417), .Q(n501) );
  AO22X1 U464 ( .IN1(n503), .IN2(n427), .IN3(n447), .IN4(n502), .Q(n179) );
  XOR2X1 U465 ( .IN1(b[7]), .IN2(n417), .Q(n502) );
  AO22X1 U466 ( .IN1(n504), .IN2(n427), .IN3(n447), .IN4(n503), .Q(n178) );
  AO22X1 U467 ( .IN1(n448), .IN2(n427), .IN3(n447), .IN4(n504), .Q(n177) );
  XOR2X1 U468 ( .IN1(n401), .IN2(n417), .Q(n504) );
  XOR2X1 U469 ( .IN1(b[10]), .IN2(n417), .Q(n448) );
  OAI21X1 U470 ( .IN1(n427), .IN2(n447), .IN3(n446), .QN(n176) );
  XOR2X1 U471 ( .IN1(b[11]), .IN2(n417), .Q(n446) );
  NOR2X0 U472 ( .IN1(n505), .IN2(n432), .QN(n175) );
  AO22X1 U473 ( .IN1(n506), .IN2(n429), .IN3(n450), .IN4(n507), .Q(n174) );
  XOR2X1 U474 ( .IN1(n414), .IN2(n418), .Q(n507) );
  AO22X1 U475 ( .IN1(n508), .IN2(n429), .IN3(n450), .IN4(n506), .Q(n173) );
  AO22X1 U476 ( .IN1(n509), .IN2(n429), .IN3(n450), .IN4(n508), .Q(n172) );
  AO22X1 U477 ( .IN1(n510), .IN2(n429), .IN3(n450), .IN4(n509), .Q(n171) );
  AO22X1 U478 ( .IN1(n511), .IN2(n429), .IN3(n450), .IN4(n510), .Q(n170) );
  AO22X1 U479 ( .IN1(n512), .IN2(n429), .IN3(n450), .IN4(n511), .Q(n169) );
  XOR2X1 U480 ( .IN1(n409), .IN2(n418), .Q(n511) );
  AO22X1 U481 ( .IN1(n513), .IN2(n429), .IN3(n450), .IN4(n512), .Q(n168) );
  XOR2X1 U482 ( .IN1(n404), .IN2(n418), .Q(n512) );
  AO22X1 U483 ( .IN1(n514), .IN2(n429), .IN3(n450), .IN4(n513), .Q(n167) );
  XOR2X1 U484 ( .IN1(b[7]), .IN2(n418), .Q(n513) );
  AO22X1 U485 ( .IN1(n515), .IN2(n429), .IN3(n450), .IN4(n514), .Q(n166) );
  AO22X1 U486 ( .IN1(n451), .IN2(n429), .IN3(n450), .IN4(n515), .Q(n165) );
  XOR2X1 U487 ( .IN1(n401), .IN2(n418), .Q(n515) );
  XOR2X1 U488 ( .IN1(b[10]), .IN2(n418), .Q(n451) );
  OAI21X1 U489 ( .IN1(n429), .IN2(n450), .IN3(n449), .QN(n164) );
  XOR2X1 U490 ( .IN1(b[11]), .IN2(n418), .Q(n449) );
  NOR2X0 U491 ( .IN1(n516), .IN2(n432), .QN(n163) );
  AO22X1 U492 ( .IN1(n517), .IN2(n431), .IN3(n453), .IN4(n518), .Q(n162) );
  XOR2X1 U493 ( .IN1(n414), .IN2(n413), .Q(n518) );
  AO22X1 U494 ( .IN1(n519), .IN2(n431), .IN3(n453), .IN4(n517), .Q(n161) );
  AO22X1 U495 ( .IN1(n520), .IN2(n431), .IN3(n453), .IN4(n519), .Q(n160) );
  AO22X1 U496 ( .IN1(n521), .IN2(n431), .IN3(n453), .IN4(n520), .Q(n159) );
  AO22X1 U497 ( .IN1(n522), .IN2(n431), .IN3(n453), .IN4(n521), .Q(n158) );
  AO22X1 U498 ( .IN1(n523), .IN2(n431), .IN3(n453), .IN4(n522), .Q(n157) );
  XOR2X1 U499 ( .IN1(n409), .IN2(n413), .Q(n522) );
  AO22X1 U500 ( .IN1(n524), .IN2(n431), .IN3(n453), .IN4(n523), .Q(n156) );
  XOR2X1 U501 ( .IN1(n404), .IN2(n413), .Q(n523) );
  AO22X1 U502 ( .IN1(n525), .IN2(n431), .IN3(n453), .IN4(n524), .Q(n155) );
  XOR2X1 U503 ( .IN1(b[7]), .IN2(n413), .Q(n524) );
  AO22X1 U504 ( .IN1(n526), .IN2(n431), .IN3(n453), .IN4(n525), .Q(n154) );
  XOR2X1 U505 ( .IN1(n408), .IN2(n413), .Q(n525) );
  AO22X1 U506 ( .IN1(n454), .IN2(n431), .IN3(n453), .IN4(n526), .Q(n153) );
  XOR2X1 U507 ( .IN1(n401), .IN2(n413), .Q(n526) );
  XOR2X1 U508 ( .IN1(b[10]), .IN2(n413), .Q(n454) );
  OAI21X1 U509 ( .IN1(n431), .IN2(n453), .IN3(n452), .QN(n152) );
  XOR2X1 U510 ( .IN1(b[11]), .IN2(n413), .Q(n452) );
  AO22X1 U511 ( .IN1(n527), .IN2(n416), .IN3(n444), .IN4(n416), .Q(n149) );
  XOR2X1 U512 ( .IN1(n416), .IN2(a[4]), .Q(n528) );
  NOR2X0 U513 ( .IN1(n414), .IN2(n473), .QN(n527) );
  XNOR2X1 U514 ( .IN1(a[4]), .IN2(n415), .Q(n473) );
  AO22X1 U515 ( .IN1(n529), .IN2(n417), .IN3(n447), .IN4(n417), .Q(n148) );
  XOR2X1 U516 ( .IN1(n417), .IN2(a[6]), .Q(n530) );
  NOR2X0 U517 ( .IN1(n414), .IN2(n494), .QN(n529) );
  XNOR2X1 U518 ( .IN1(a[6]), .IN2(n416), .Q(n494) );
  AO22X1 U519 ( .IN1(n531), .IN2(n418), .IN3(n450), .IN4(n418), .Q(n147) );
  XOR2X1 U520 ( .IN1(n418), .IN2(a[8]), .Q(n532) );
  NOR2X0 U521 ( .IN1(n414), .IN2(n505), .QN(n531) );
  XNOR2X1 U522 ( .IN1(a[8]), .IN2(n417), .Q(n505) );
  AO22X1 U523 ( .IN1(n533), .IN2(n413), .IN3(n453), .IN4(n413), .Q(n146) );
  NOR2X0 U524 ( .IN1(n414), .IN2(n516), .QN(n533) );
  XNOR2X1 U525 ( .IN1(a[10]), .IN2(n418), .Q(n516) );
endmodule


module mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1 ( in_a, in_b, clk, 
        \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [11:0] \output ;
  input clk;
  wire   n3, n4, n5, n6, n1, n2, n7, n8, n9, n10, n11, n12, n13;
  wire   [23:7] pre_out;
  wire   [23:7] pre_out_reg;
  wire   [11:0] rnd_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  DFFX1 \pre_out_reg_reg[23]  ( .D(pre_out[23]), .CLK(clk), .Q(pre_out_reg[23]), .QN(n7) );
  DFFX1 \pre_out_reg_reg[22]  ( .D(pre_out[22]), .CLK(clk), .Q(pre_out_reg[22]), .QN(n2) );
  DFFX1 \pre_out_reg_reg[21]  ( .D(pre_out[21]), .CLK(clk), .Q(pre_out_reg[21]), .QN(n3) );
  DFFX1 \pre_out_reg_reg[20]  ( .D(pre_out[20]), .CLK(clk), .Q(n1), .QN(n4) );
  DFFX1 \pre_out_reg_reg[19]  ( .D(pre_out[19]), .CLK(clk), .Q(pre_out_reg[19]), .QN(n5) );
  DFFX1 \pre_out_reg_reg[18]  ( .D(pre_out[18]), .CLK(clk), .Q(pre_out_reg[18]) );
  DFFX1 \pre_out_reg_reg[17]  ( .D(pre_out[17]), .CLK(clk), .Q(pre_out_reg[17]) );
  DFFX1 \pre_out_reg_reg[16]  ( .D(pre_out[16]), .CLK(clk), .Q(pre_out_reg[16]) );
  DFFX1 \pre_out_reg_reg[15]  ( .D(pre_out[15]), .CLK(clk), .Q(pre_out_reg[15]) );
  DFFX1 \pre_out_reg_reg[14]  ( .D(pre_out[14]), .CLK(clk), .Q(pre_out_reg[14]) );
  DFFX1 \pre_out_reg_reg[13]  ( .D(pre_out[13]), .CLK(clk), .Q(pre_out_reg[13]) );
  DFFX1 \pre_out_reg_reg[12]  ( .D(pre_out[12]), .CLK(clk), .Q(pre_out_reg[12]) );
  DFFX1 \pre_out_reg_reg[11]  ( .D(pre_out[11]), .CLK(clk), .Q(pre_out_reg[11]) );
  DFFX1 \pre_out_reg_reg[10]  ( .D(pre_out[10]), .CLK(clk), .Q(pre_out_reg[10]) );
  DFFX1 \pre_out_reg_reg[9]  ( .D(pre_out[9]), .CLK(clk), .Q(pre_out_reg[9])
         );
  DFFX1 \pre_out_reg_reg[8]  ( .D(pre_out[8]), .CLK(clk), .Q(pre_out_reg[8])
         );
  DFFX1 \pre_out_reg_reg[7]  ( .D(pre_out[7]), .CLK(clk), .Q(pre_out_reg[7])
         );
  AO21X1 U8 ( .IN1(rnd_out[9]), .IN2(n6), .IN3(n10), .Q(\output [9]) );
  AO21X1 U9 ( .IN1(rnd_out[8]), .IN2(n6), .IN3(n10), .Q(\output [8]) );
  AO21X1 U10 ( .IN1(rnd_out[7]), .IN2(n6), .IN3(n10), .Q(\output [7]) );
  AO21X1 U11 ( .IN1(rnd_out[6]), .IN2(n6), .IN3(n10), .Q(\output [6]) );
  AO21X1 U12 ( .IN1(rnd_out[5]), .IN2(n6), .IN3(n10), .Q(\output [5]) );
  AO21X1 U13 ( .IN1(rnd_out[4]), .IN2(n6), .IN3(n10), .Q(\output [4]) );
  AO21X1 U14 ( .IN1(rnd_out[3]), .IN2(n6), .IN3(n10), .Q(\output [3]) );
  AO21X1 U15 ( .IN1(rnd_out[2]), .IN2(n6), .IN3(n10), .Q(\output [2]) );
  AO21X1 U16 ( .IN1(rnd_out[1]), .IN2(n6), .IN3(n10), .Q(\output [1]) );
  AO21X1 U18 ( .IN1(rnd_out[10]), .IN2(n6), .IN3(n10), .Q(\output [10]) );
  AO21X1 U19 ( .IN1(rnd_out[0]), .IN2(n6), .IN3(n10), .Q(\output [0]) );
  mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_DW01_inc_0 add_48_round ( .A(
        pre_out_reg[19:7]), .SUM({rnd_out, SYNOPSYS_UNCONNECTED__0}) );
  mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1_DW_mult_tc_0 mult_37 ( .a({
        in_a[11:2], n9, in_a[0]}), .b(in_b), .product({pre_out, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7}) );
  INVX0 U3 ( .INP(in_a[1]), .ZN(n8) );
  INVX1 U4 ( .INP(n8), .ZN(n9) );
  INVX0 U5 ( .INP(n13), .ZN(n6) );
  AND2X1 U6 ( .IN1(n13), .IN2(n7), .Q(n10) );
  NAND4X0 U7 ( .IN1(n4), .IN2(n3), .IN3(n5), .IN4(n2), .QN(n12) );
  NAND4X0 U17 ( .IN1(pre_out_reg[21]), .IN2(pre_out_reg[22]), .IN3(n1), .IN4(
        pre_out_reg[19]), .QN(n11) );
  MUX21X1 U20 ( .IN1(n12), .IN2(n11), .S(pre_out_reg[23]), .Q(n13) );
  MUX21X1 U21 ( .IN1(pre_out_reg[23]), .IN2(rnd_out[11]), .S(n6), .Q(
        \output [11]) );
endmodule



    module shifter_WORD_WIDTH12_LOG_WORD_WIDTH4_SMALLER_POW2_WW16_MAX_LEFT8_MAX_RIGHT3 ( 
        \input , \output , direction, amount );
  input [11:0] \input ;
  output [11:0] \output ;
  input [3:0] amount;
  input direction;
  wire   N2, N3, N4, N5, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143;
  assign N2 = amount[0];
  assign N3 = amount[1];
  assign N4 = amount[2];
  assign N5 = amount[3];

  AND4X4 U2 ( .IN1(n4), .IN2(n140), .IN3(n25), .IN4(n45), .Q(n1) );
  INVX0 U3 ( .INP(n119), .ZN(n2) );
  AO22X2 U4 ( .IN1(n2), .IN2(\input [0]), .IN3(n40), .IN4(n41), .Q(N28) );
  MUX21X1 U5 ( .IN1(n68), .IN2(n63), .S(n12), .Q(n55) );
  AND2X4 U6 ( .IN1(n85), .IN2(n24), .Q(n28) );
  AND3X1 U7 ( .IN1(n28), .IN2(n138), .IN3(n22), .Q(n8) );
  MUX21X1 U8 ( .IN1(n96), .IN2(n97), .S(n18), .Q(n84) );
  INVX0 U9 ( .INP(n8), .ZN(n136) );
  DELLN2X2 U10 ( .INP(n25), .Z(n3) );
  INVX0 U11 ( .INP(N5), .ZN(n4) );
  DELLN2X2 U12 ( .INP(n36), .Z(n5) );
  NAND2X0 U13 ( .IN1(n76), .IN2(n77), .QN(n75) );
  AO22X1 U14 ( .IN1(\input [4]), .IN2(n24), .IN3(N4), .IN4(\input [0]), .Q(n63) );
  OR2X4 U15 ( .IN1(n68), .IN2(n139), .Q(n65) );
  INVX0 U16 ( .INP(n1), .ZN(n6) );
  INVX0 U17 ( .INP(n6), .ZN(n7) );
  AO22X1 U18 ( .IN1(N15), .IN2(n142), .IN3(N27), .IN4(n143), .Q(\output [3])
         );
  OAI221X1 U19 ( .IN1(n69), .IN2(n57), .IN3(n48), .IN4(n70), .IN5(n71), .QN(
        N22) );
  INVX0 U20 ( .INP(n16), .ZN(n9) );
  OR2X1 U21 ( .IN1(n72), .IN2(n13), .Q(n66) );
  AO22X1 U22 ( .IN1(\input [6]), .IN2(n25), .IN3(n17), .IN4(\input [2]), .Q(
        n72) );
  OR2X1 U23 ( .IN1(N2), .IN2(n63), .Q(n51) );
  NAND3X1 U24 ( .IN1(n30), .IN2(\input [2]), .IN3(n22), .QN(n108) );
  NAND2X0 U25 ( .IN1(\input [4]), .IN2(n39), .QN(n110) );
  AO22X2 U26 ( .IN1(n40), .IN2(n67), .IN3(n62), .IN4(n55), .Q(N23) );
  NAND2X0 U27 ( .IN1(n65), .IN2(n66), .QN(n70) );
  AND2X2 U28 ( .IN1(n85), .IN2(n38), .Q(n19) );
  INVX0 U29 ( .INP(n40), .ZN(n10) );
  INVX0 U30 ( .INP(n10), .ZN(n11) );
  INVX0 U31 ( .INP(n137), .ZN(n12) );
  INVX0 U32 ( .INP(n137), .ZN(n13) );
  DELLN1X2 U33 ( .INP(N5), .Z(n14) );
  INVX0 U34 ( .INP(n20), .ZN(n15) );
  MUX21X2 U35 ( .IN1(n91), .IN2(n92), .S(n14), .Q(n90) );
  INVX0 U36 ( .INP(N4), .ZN(n16) );
  INVX0 U37 ( .INP(n16), .ZN(n17) );
  NAND2X0 U38 ( .IN1(n102), .IN2(n4), .QN(n101) );
  NAND2X0 U39 ( .IN1(\input [0]), .IN2(n8), .QN(n34) );
  NAND2X0 U40 ( .IN1(\input [10]), .IN2(n8), .QN(n79) );
  INVX0 U41 ( .INP(n139), .ZN(n141) );
  INVX0 U42 ( .INP(n3), .ZN(n18) );
  MUX21X2 U43 ( .IN1(\input [11]), .IN2(\input [7]), .S(n18), .Q(n32) );
  MUX21X2 U44 ( .IN1(n98), .IN2(n87), .S(n18), .Q(n95) );
  MUX21X1 U45 ( .IN1(n36), .IN2(n52), .S(n139), .Q(n42) );
  INVX0 U46 ( .INP(n45), .ZN(n20) );
  OA221X1 U47 ( .IN1(n21), .IN2(n43), .IN3(n44), .IN4(n15), .IN5(n28), .Q(N27)
         );
  NAND2X0 U48 ( .IN1(n61), .IN2(n60), .QN(N24) );
  NBUFFX4 U49 ( .INP(N3), .Z(n21) );
  INVX0 U50 ( .INP(N3), .ZN(n22) );
  INVX0 U51 ( .INP(n28), .ZN(n23) );
  INVX0 U52 ( .INP(N4), .ZN(n24) );
  INVX0 U53 ( .INP(N4), .ZN(n25) );
  AND2X4 U54 ( .IN1(n14), .IN2(n15), .Q(n31) );
  MUX21X2 U55 ( .IN1(n74), .IN2(n103), .S(n20), .Q(n102) );
  MUX21X2 U56 ( .IN1(n133), .IN2(n33), .S(n20), .Q(n132) );
  OAI221X2 U57 ( .IN1(n87), .IN2(n115), .IN3(n21), .IN4(n116), .IN5(n117), 
        .QN(N14) );
  AND2X1 U58 ( .IN1(n76), .IN2(n77), .Q(n26) );
  INVX0 U59 ( .INP(n119), .ZN(n39) );
  INVX0 U60 ( .INP(n48), .ZN(n62) );
  AND2X1 U61 ( .IN1(n139), .IN2(n31), .Q(n27) );
  AND3X1 U62 ( .IN1(n21), .IN2(n12), .IN3(n28), .Q(n29) );
  INVX0 U63 ( .INP(direction), .ZN(n143) );
  AND3X1 U64 ( .IN1(n38), .IN2(n138), .IN3(n4), .Q(n30) );
  INVX0 U65 ( .INP(n42), .ZN(n41) );
  INVX0 U66 ( .INP(n52), .ZN(n88) );
  INVX0 U67 ( .INP(n34), .ZN(N30) );
  INVX0 U68 ( .INP(\input [2]), .ZN(n59) );
  AND2X1 U69 ( .IN1(n47), .IN2(n46), .Q(n43) );
  INVX0 U70 ( .INP(n5), .ZN(n74) );
  NOR2X0 U71 ( .IN1(n33), .IN2(n136), .QN(N7) );
  NOR2X0 U72 ( .IN1(n131), .IN2(n132), .QN(N9) );
  INVX0 U73 ( .INP(n64), .ZN(n103) );
  INVX0 U74 ( .INP(n79), .ZN(n135) );
  NAND4X0 U75 ( .IN1(n31), .IN2(\input [0]), .IN3(n3), .IN4(n138), .QN(n71) );
  INVX0 U76 ( .INP(n33), .ZN(n128) );
  INVX0 U77 ( .INP(n94), .ZN(n73) );
  INVX0 U78 ( .INP(\input [3]), .ZN(n58) );
  NAND2X0 U79 ( .IN1(\input [3]), .IN2(n39), .QN(n106) );
  NAND2X0 U80 ( .IN1(\input [1]), .IN2(n8), .QN(n105) );
  INVX0 U81 ( .INP(\input [7]), .ZN(n123) );
  INVX0 U82 ( .INP(\input [5]), .ZN(n87) );
  INVX0 U83 ( .INP(\input [6]), .ZN(n86) );
  INVX0 U84 ( .INP(\input [11]), .ZN(n33) );
  NOR2X0 U85 ( .IN1(n141), .IN2(n64), .QN(n92) );
  INVX0 U86 ( .INP(n78), .ZN(n130) );
  INVX0 U87 ( .INP(\input [9]), .ZN(n98) );
  INVX0 U88 ( .INP(\input [8]), .ZN(n96) );
  INVX0 U89 ( .INP(\input [4]), .ZN(n97) );
  INVX0 U90 ( .INP(\input [10]), .ZN(n134) );
  NOR3X0 U91 ( .IN1(n35), .IN2(n20), .IN3(n14), .QN(N29) );
  MUX21X1 U92 ( .IN1(n36), .IN2(n37), .S(n12), .Q(n35) );
  OA22X1 U93 ( .IN1(\input [0]), .IN2(n139), .IN3(\input [1]), .IN4(n12), .Q(
        n44) );
  OAI21X1 U94 ( .IN1(n42), .IN2(n48), .IN3(n49), .QN(N26) );
  NAND3X0 U95 ( .IN1(n56), .IN2(n50), .IN3(n51), .QN(n49) );
  NAND4X0 U96 ( .IN1(n19), .IN2(n47), .IN3(n46), .IN4(n20), .QN(n53) );
  NAND2X1 U97 ( .IN1(n139), .IN2(n58), .QN(n46) );
  NAND3X0 U98 ( .IN1(n62), .IN2(n50), .IN3(n51), .QN(n61) );
  NAND3X0 U99 ( .IN1(n65), .IN2(n66), .IN3(n40), .QN(n60) );
  AO222X1 U100 ( .IN1(n73), .IN2(n11), .IN3(n74), .IN4(n27), .IN5(n62), .IN6(
        n67), .Q(N21) );
  MUX21X1 U101 ( .IN1(n75), .IN2(n72), .S(n13), .Q(n67) );
  NAND4X0 U102 ( .IN1(n78), .IN2(n79), .IN3(n80), .IN4(n81), .QN(N20) );
  OA22X1 U103 ( .IN1(n82), .IN2(n83), .IN3(n69), .IN4(n48), .Q(n81) );
  MUX21X1 U104 ( .IN1(n84), .IN2(n26), .S(n141), .Q(n69) );
  MUX21X1 U105 ( .IN1(n86), .IN2(n87), .S(n141), .Q(n82) );
  NAND2X1 U106 ( .IN1(n88), .IN2(n27), .QN(n80) );
  AO222X1 U107 ( .IN1(n7), .IN2(\input [10]), .IN3(n73), .IN4(n62), .IN5(n90), 
        .IN6(n15), .Q(N19) );
  MUX21X1 U108 ( .IN1(n32), .IN2(n93), .S(n141), .Q(n91) );
  MUX21X1 U109 ( .IN1(n95), .IN2(n84), .S(n141), .Q(n94) );
  NAND2X1 U110 ( .IN1(n34), .IN2(n99), .QN(N18) );
  MUX21X1 U111 ( .IN1(n100), .IN2(n101), .S(n141), .Q(n99) );
  NAND2X1 U112 ( .IN1(n88), .IN2(n62), .QN(n100) );
  NAND4X0 U113 ( .IN1(n107), .IN2(n104), .IN3(n106), .IN4(n105), .QN(N17) );
  NAND4X0 U114 ( .IN1(n108), .IN2(n109), .IN3(n110), .IN4(n111), .QN(N16) );
  NAND4X0 U115 ( .IN1(n19), .IN2(n20), .IN3(\input [5]), .IN4(n12), .QN(n111)
         );
  AO221X1 U116 ( .IN1(\input [5]), .IN2(n2), .IN3(n89), .IN4(\input [4]), 
        .IN5(n112), .Q(N15) );
  NAND4X0 U117 ( .IN1(n19), .IN2(n21), .IN3(\input [6]), .IN4(n12), .QN(n114)
         );
  NAND4X0 U118 ( .IN1(n22), .IN2(n28), .IN3(\input [3]), .IN4(n138), .QN(n113)
         );
  OA22X1 U119 ( .IN1(n22), .IN2(n118), .IN3(n119), .IN4(n86), .Q(n117) );
  NAND4X0 U120 ( .IN1(n4), .IN2(n25), .IN3(n140), .IN4(\input [7]), .QN(n118)
         );
  NAND2X1 U121 ( .IN1(n30), .IN2(\input [4]), .QN(n116) );
  NAND3X0 U122 ( .IN1(n120), .IN2(n121), .IN3(n122), .QN(N13) );
  OA22X1 U123 ( .IN1(n119), .IN2(n123), .IN3(n86), .IN4(n115), .Q(n122) );
  NAND4X0 U124 ( .IN1(n19), .IN2(n21), .IN3(\input [8]), .IN4(n13), .QN(n121)
         );
  NAND4X0 U125 ( .IN1(n19), .IN2(n22), .IN3(\input [5]), .IN4(n139), .QN(n120)
         );
  AO221X1 U126 ( .IN1(\input [8]), .IN2(n2), .IN3(n89), .IN4(\input [7]), 
        .IN5(n124), .Q(N12) );
  NAND4X0 U127 ( .IN1(n19), .IN2(n21), .IN3(\input [9]), .IN4(n13), .QN(n126)
         );
  NAND4X0 U128 ( .IN1(n19), .IN2(n22), .IN3(\input [6]), .IN4(n139), .QN(n125)
         );
  AO221X1 U129 ( .IN1(\input [8]), .IN2(n1), .IN3(\input [7]), .IN4(n8), .IN5(
        n127), .Q(N11) );
  AO22X1 U130 ( .IN1(\input [9]), .IN2(n39), .IN3(n29), .IN4(\input [10]), .Q(
        n127) );
  AO221X1 U131 ( .IN1(n29), .IN2(n128), .IN3(\input [10]), .IN4(n2), .IN5(n129), .Q(N10) );
  AO21X1 U132 ( .IN1(\input [8]), .IN2(n8), .IN3(n130), .Q(n129) );
  NAND4X0 U133 ( .IN1(n85), .IN2(n38), .IN3(n138), .IN4(N3), .QN(n119) );
  MUX21X1 U134 ( .IN1(n98), .IN2(n134), .S(n141), .Q(n133) );
  OA22X1 U135 ( .IN1(n20), .IN2(n23), .IN3(n141), .IN4(n23), .Q(n131) );
  AO21X1 U136 ( .IN1(n7), .IN2(n128), .IN3(n135), .Q(N8) );
  NAND4X0 U137 ( .IN1(n4), .IN2(n140), .IN3(n25), .IN4(n45), .QN(n115) );
  INVX0 U138 ( .INP(n137), .ZN(n140) );
  INVX0 U139 ( .INP(N2), .ZN(n137) );
  NAND2X0 U140 ( .IN1(n40), .IN2(n55), .QN(n54) );
  INVX0 U141 ( .INP(N3), .ZN(n45) );
  NAND2X0 U142 ( .IN1(n4), .IN2(n45), .QN(n57) );
  NAND2X0 U143 ( .IN1(\input [3]), .IN2(n25), .QN(n64) );
  NAND2X0 U144 ( .IN1(\input [1]), .IN2(n25), .QN(n36) );
  NAND2X0 U145 ( .IN1(\input [2]), .IN2(n24), .QN(n52) );
  NAND2X0 U146 ( .IN1(\input [7]), .IN2(n24), .QN(n76) );
  NAND2X0 U147 ( .IN1(\input [3]), .IN2(n17), .QN(n77) );
  NAND2X0 U148 ( .IN1(\input [0]), .IN2(n38), .QN(n37) );
  NOR2X0 U149 ( .IN1(n3), .IN2(n86), .QN(n93) );
  NAND2X0 U150 ( .IN1(n18), .IN2(n11), .QN(n83) );
  NAND2X0 U151 ( .IN1(n53), .IN2(n54), .QN(N25) );
  NAND2X0 U152 ( .IN1(n113), .IN2(n114), .QN(n112) );
  NAND2X0 U153 ( .IN1(n13), .IN2(n59), .QN(n47) );
  INVX0 U154 ( .INP(n57), .ZN(n40) );
  INVX0 U155 ( .INP(n115), .ZN(n89) );
  INVX0 U156 ( .INP(N4), .ZN(n38) );
  INVX0 U157 ( .INP(N5), .ZN(n85) );
  NAND2X0 U158 ( .IN1(n29), .IN2(\input [4]), .QN(n107) );
  NAND2X0 U159 ( .IN1(n4), .IN2(N3), .QN(n48) );
  INVX0 U160 ( .INP(N2), .ZN(n138) );
  INVX0 U161 ( .INP(N2), .ZN(n139) );
  AO22X1 U162 ( .IN1(\input [5]), .IN2(n38), .IN3(n9), .IN4(\input [1]), .Q(
        n68) );
  NAND2X0 U163 ( .IN1(n140), .IN2(n64), .QN(n50) );
  NAND2X0 U164 ( .IN1(n125), .IN2(n126), .QN(n124) );
  NAND2X0 U165 ( .IN1(\input [9]), .IN2(n7), .QN(n78) );
  NAND2X0 U166 ( .IN1(\input [2]), .IN2(n1), .QN(n104) );
  NAND2X0 U167 ( .IN1(\input [3]), .IN2(n89), .QN(n109) );
  INVX0 U168 ( .INP(n57), .ZN(n56) );
  INVX0 U169 ( .INP(n143), .ZN(n142) );
  MUX21X1 U170 ( .IN1(N30), .IN2(N18), .S(n142), .Q(\output [0]) );
  AO22X1 U171 ( .IN1(N29), .IN2(n143), .IN3(n142), .IN4(N17), .Q(\output [1])
         );
  AO22X1 U172 ( .IN1(N28), .IN2(n143), .IN3(N16), .IN4(n142), .Q(\output [2])
         );
  AO22X1 U173 ( .IN1(N26), .IN2(n143), .IN3(N14), .IN4(n142), .Q(\output [4])
         );
  AO22X1 U174 ( .IN1(n143), .IN2(N25), .IN3(N13), .IN4(n142), .Q(\output [5])
         );
  AO22X1 U175 ( .IN1(n143), .IN2(N24), .IN3(N12), .IN4(n142), .Q(\output [6])
         );
  AO22X1 U176 ( .IN1(N23), .IN2(n143), .IN3(N11), .IN4(n142), .Q(\output [7])
         );
  MUX21X1 U177 ( .IN1(N22), .IN2(N10), .S(n142), .Q(\output [8]) );
  MUX21X1 U178 ( .IN1(N21), .IN2(N9), .S(n142), .Q(\output [9]) );
  MUX21X1 U179 ( .IN1(N20), .IN2(N8), .S(n142), .Q(\output [10]) );
  MUX21X1 U180 ( .IN1(N19), .IN2(N7), .S(n142), .Q(\output [11]) );
endmodule



    module shifter_WORD_WIDTH12_LOG_WORD_WIDTH4_SMALLER_POW2_WW16_MAX_LEFT4_MAX_RIGHT2 ( 
        \input , \output , direction, amount );
  input [11:0] \input ;
  output [11:0] \output ;
  input [3:0] amount;
  input direction;
  wire   N2, N3, N4, N5, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118;
  assign N2 = amount[0];
  assign N3 = amount[1];
  assign N4 = amount[2];
  assign N5 = amount[3];

  NAND2X0 U2 ( .IN1(N2), .IN2(n19), .QN(n110) );
  NAND2X0 U3 ( .IN1(n29), .IN2(n23), .QN(n36) );
  NAND2X0 U4 ( .IN1(n11), .IN2(n29), .QN(n45) );
  NAND2X0 U5 ( .IN1(n29), .IN2(n61), .QN(n74) );
  NAND2X0 U6 ( .IN1(n29), .IN2(n83), .QN(n66) );
  NAND2X0 U7 ( .IN1(n1), .IN2(n29), .QN(n22) );
  NAND2X0 U8 ( .IN1(n19), .IN2(n29), .QN(n113) );
  NAND2X0 U9 ( .IN1(N3), .IN2(n29), .QN(n99) );
  MUX21X1 U10 ( .IN1(N19), .IN2(N7), .S(n117), .Q(\output [11]) );
  AO22X1 U11 ( .IN1(N24), .IN2(n118), .IN3(N12), .IN4(n117), .Q(\output [6])
         );
  OAI222X1 U12 ( .IN1(n15), .IN2(n68), .IN3(n34), .IN4(n57), .IN5(n7), .IN6(
        n103), .QN(N13) );
  AND2X4 U13 ( .IN1(N3), .IN2(n17), .Q(n1) );
  AND2X4 U14 ( .IN1(N2), .IN2(n10), .Q(n2) );
  AND2X4 U15 ( .IN1(N4), .IN2(n73), .Q(n3) );
  AND3X1 U16 ( .IN1(n87), .IN2(n85), .IN3(n86), .Q(n4) );
  MUX21X2 U17 ( .IN1(N13), .IN2(N25), .S(n118), .Q(\output [5]) );
  NAND3X1 U18 ( .IN1(n48), .IN2(n102), .IN3(n49), .QN(N24) );
  NAND3X1 U19 ( .IN1(n12), .IN2(N2), .IN3(\input [4]), .QN(n54) );
  OR2X1 U20 ( .IN1(n29), .IN2(\input [1]), .Q(n25) );
  NAND2X0 U21 ( .IN1(\input [3]), .IN2(n1), .QN(n5) );
  NAND2X0 U22 ( .IN1(N4), .IN2(n78), .QN(n33) );
  AO22X1 U23 ( .IN1(n117), .IN2(N14), .IN3(N26), .IN4(n118), .Q(\output [4])
         );
  NAND3X0 U24 ( .IN1(n63), .IN2(n64), .IN3(n65), .QN(N22) );
  AO22X1 U25 ( .IN1(N21), .IN2(n118), .IN3(N9), .IN4(n117), .Q(\output [9]) );
  AO22X1 U26 ( .IN1(n118), .IN2(N23), .IN3(N11), .IN4(n117), .Q(\output [7])
         );
  NAND2X0 U27 ( .IN1(n4), .IN2(n84), .QN(N19) );
  NAND2X0 U28 ( .IN1(n13), .IN2(n98), .QN(n85) );
  NAND2X0 U29 ( .IN1(n104), .IN2(n14), .QN(n86) );
  INVX0 U30 ( .INP(n58), .ZN(n6) );
  INVX0 U31 ( .INP(n6), .ZN(n7) );
  NAND3X1 U32 ( .IN1(n93), .IN2(n92), .IN3(\input [1]), .QN(n90) );
  MUX21X2 U33 ( .IN1(N17), .IN2(N29), .S(n118), .Q(\output [1]) );
  MUX21X2 U34 ( .IN1(N27), .IN2(N15), .S(n117), .Q(\output [3]) );
  NAND2X0 U35 ( .IN1(\input [3]), .IN2(n1), .QN(n43) );
  NAND3X4 U36 ( .IN1(n36), .IN2(n25), .IN3(n1), .QN(n30) );
  NAND2X0 U37 ( .IN1(n9), .IN2(n25), .QN(n24) );
  MUX21X2 U38 ( .IN1(n28), .IN2(n16), .S(N2), .Q(n27) );
  AND2X4 U39 ( .IN1(n6), .IN2(n17), .Q(n8) );
  NAND3X2 U40 ( .IN1(n10), .IN2(n29), .IN3(\input [7]), .QN(n70) );
  NAND2X0 U41 ( .IN1(N2), .IN2(n58), .QN(n67) );
  NAND3X1 U42 ( .IN1(n12), .IN2(n29), .IN3(\input [5]), .QN(n55) );
  NAND2X0 U43 ( .IN1(n2), .IN2(\input [6]), .QN(n72) );
  NAND2X0 U44 ( .IN1(n3), .IN2(\input [5]), .QN(n71) );
  NAND3X1 U45 ( .IN1(\input [0]), .IN2(n78), .IN3(n92), .QN(n91) );
  NAND2X0 U46 ( .IN1(\input [11]), .IN2(n100), .QN(n87) );
  INVX0 U47 ( .INP(n22), .ZN(n101) );
  INVX0 U48 ( .INP(n113), .ZN(n108) );
  INVX0 U49 ( .INP(n15), .ZN(n100) );
  NOR2X0 U50 ( .IN1(n110), .IN2(n83), .QN(n107) );
  INVX0 U51 ( .INP(n49), .ZN(n106) );
  INVX0 U52 ( .INP(n25), .ZN(n20) );
  INVX0 U53 ( .INP(n110), .ZN(n98) );
  INVX0 U54 ( .INP(n34), .ZN(n50) );
  INVX0 U55 ( .INP(n77), .ZN(n59) );
  INVX0 U56 ( .INP(N2), .ZN(n29) );
  NOR2X0 U57 ( .IN1(n15), .IN2(n16), .QN(N30) );
  NOR2X0 U58 ( .IN1(n83), .IN2(n99), .QN(n105) );
  INVX0 U59 ( .INP(n92), .ZN(n95) );
  NOR2X0 U60 ( .IN1(n33), .IN2(n28), .QN(n42) );
  INVX0 U61 ( .INP(n45), .ZN(n44) );
  INVX0 U62 ( .INP(\input [1]), .ZN(n28) );
  INVX0 U63 ( .INP(n47), .ZN(n46) );
  INVX0 U64 ( .INP(\input [8]), .ZN(n83) );
  INVX0 U65 ( .INP(n33), .ZN(n62) );
  INVX0 U66 ( .INP(\input [0]), .ZN(n16) );
  INVX0 U67 ( .INP(\input [6]), .ZN(n57) );
  INVX0 U68 ( .INP(\input [4]), .ZN(n51) );
  INVX0 U69 ( .INP(n27), .ZN(n18) );
  INVX0 U70 ( .INP(n99), .ZN(n104) );
  AND2X1 U71 ( .IN1(n17), .IN2(n19), .Q(n9) );
  NAND3X1 U72 ( .IN1(\input [2]), .IN2(N2), .IN3(n1), .QN(n40) );
  INVX0 U73 ( .INP(n86), .ZN(n109) );
  INVX0 U74 ( .INP(n94), .ZN(n93) );
  INVX0 U75 ( .INP(n97), .ZN(n78) );
  INVX0 U76 ( .INP(\input [2]), .ZN(n23) );
  INVX0 U77 ( .INP(\input [3]), .ZN(n35) );
  AND2X1 U78 ( .IN1(N3), .IN2(n73), .Q(n10) );
  NAND3X0 U79 ( .IN1(n1), .IN2(n92), .IN3(\input [2]), .QN(n89) );
  INVX0 U80 ( .INP(n114), .ZN(n17) );
  INVX0 U81 ( .INP(N4), .ZN(n61) );
  INVX0 U82 ( .INP(N3), .ZN(n19) );
  NOR2X0 U83 ( .IN1(n113), .IN2(n114), .QN(n111) );
  INVX0 U84 ( .INP(direction), .ZN(n118) );
  INVX0 U85 ( .INP(n80), .ZN(n112) );
  AND2X1 U86 ( .IN1(n59), .IN2(n60), .Q(n11) );
  AND3X1 U87 ( .IN1(N3), .IN2(n61), .IN3(n60), .Q(n12) );
  INVX0 U88 ( .INP(n87), .ZN(N7) );
  INVX0 U89 ( .INP(n85), .ZN(n115) );
  INVX0 U90 ( .INP(n81), .ZN(n116) );
  AND2X1 U91 ( .IN1(\input [10]), .IN2(n17), .Q(n13) );
  AND2X1 U92 ( .IN1(\input [9]), .IN2(n17), .Q(n14) );
  INVX0 U93 ( .INP(N5), .ZN(n60) );
  AND3X1 U94 ( .IN1(n17), .IN2(n18), .IN3(n19), .Q(N29) );
  OAI222X1 U95 ( .IN1(n20), .IN2(n21), .IN3(n16), .IN4(n22), .IN5(n23), .IN6(
        n24), .QN(N28) );
  NAND2X1 U96 ( .IN1(n9), .IN2(N2), .QN(n21) );
  AO22X1 U97 ( .IN1(n26), .IN2(n9), .IN3(n1), .IN4(n18), .Q(N27) );
  OA22X1 U98 ( .IN1(\input [3]), .IN2(N2), .IN3(\input [2]), .IN4(n29), .Q(n26) );
  NAND3X0 U99 ( .IN1(n30), .IN2(n31), .IN3(n32), .QN(N26) );
  OA22X1 U100 ( .IN1(n16), .IN2(n33), .IN3(n34), .IN4(n35), .Q(n32) );
  NAND4X0 U101 ( .IN1(n37), .IN2(n38), .IN3(n39), .IN4(n40), .QN(N25) );
  OA222X1 U102 ( .IN1(n22), .IN2(n51), .IN3(n35), .IN4(n52), .IN5(n23), .IN6(
        n33), .Q(n48) );
  NAND4X0 U103 ( .IN1(n56), .IN2(n54), .IN3(n55), .IN4(n53), .QN(N23) );
  OA22X1 U104 ( .IN1(n47), .IN2(n57), .IN3(n45), .IN4(n7), .Q(n56) );
  NAND2X1 U105 ( .IN1(n11), .IN2(N2), .QN(n47) );
  NAND2X1 U106 ( .IN1(\input [3]), .IN2(n62), .QN(n53) );
  NAND4X0 U107 ( .IN1(n67), .IN2(n66), .IN3(n19), .IN4(n17), .QN(n64) );
  OA22X1 U108 ( .IN1(n33), .IN2(n51), .IN3(n52), .IN4(n68), .Q(n63) );
  NAND2X1 U109 ( .IN1(N2), .IN2(n1), .QN(n52) );
  NAND4X0 U110 ( .IN1(n72), .IN2(n70), .IN3(n71), .IN4(n69), .QN(N21) );
  OA21X1 U111 ( .IN1(n74), .IN2(n75), .IN3(n76), .Q(n69) );
  NAND4X0 U112 ( .IN1(n59), .IN2(N2), .IN3(n73), .IN4(\input [8]), .QN(n76) );
  NAND3X0 U113 ( .IN1(n73), .IN2(n19), .IN3(\input [9]), .QN(n75) );
  AO21X1 U114 ( .IN1(n60), .IN2(n61), .IN3(n78), .Q(n73) );
  NAND4X0 U115 ( .IN1(n79), .IN2(n82), .IN3(n81), .IN4(n80), .QN(N20) );
  NAND3X0 U116 ( .IN1(n66), .IN2(n67), .IN3(n1), .QN(n82) );
  OA21X1 U117 ( .IN1(n33), .IN2(n58), .IN3(n88), .Q(n84) );
  NAND4X0 U118 ( .IN1(N2), .IN2(N3), .IN3(\input [8]), .IN4(n17), .QN(n88) );
  NAND3X0 U119 ( .IN1(n89), .IN2(n90), .IN3(n91), .QN(N18) );
  OA221X1 U120 ( .IN1(n97), .IN2(n28), .IN3(n23), .IN4(n94), .IN5(n43), .Q(n96) );
  NAND2X1 U121 ( .IN1(n98), .IN2(n60), .QN(n94) );
  NAND2X1 U122 ( .IN1(n99), .IN2(n77), .QN(n92) );
  NAND2X1 U123 ( .IN1(n19), .IN2(n61), .QN(n77) );
  AO222X1 U124 ( .IN1(\input [4]), .IN2(n50), .IN3(\input [3]), .IN4(n100), 
        .IN5(n101), .IN6(\input [5]), .Q(N15) );
  NAND3X0 U125 ( .IN1(n65), .IN2(n102), .IN3(n31), .QN(N14) );
  NAND2X1 U126 ( .IN1(n104), .IN2(n17), .QN(n103) );
  AO221X1 U127 ( .IN1(n105), .IN2(n17), .IN3(n8), .IN4(n98), .IN5(n106), .Q(
        N12) );
  AO221X1 U128 ( .IN1(n107), .IN2(n17), .IN3(n8), .IN4(n108), .IN5(n109), .Q(
        N11) );
  AO221X1 U129 ( .IN1(n111), .IN2(\input [8]), .IN3(n104), .IN4(n13), .IN5(
        n112), .Q(N10) );
  NAND2X1 U130 ( .IN1(n14), .IN2(n98), .QN(n80) );
  AO221X1 U131 ( .IN1(\input [11]), .IN2(n101), .IN3(n14), .IN4(n108), .IN5(
        n115), .Q(N9) );
  AO21X1 U132 ( .IN1(\input [11]), .IN2(n50), .IN3(n116), .Q(N8) );
  NAND2X1 U133 ( .IN1(n13), .IN2(n108), .QN(n81) );
  NAND2X1 U134 ( .IN1(n98), .IN2(n17), .QN(n34) );
  NAND2X1 U135 ( .IN1(n60), .IN2(n61), .QN(n114) );
  NAND2X1 U136 ( .IN1(n78), .IN2(n61), .QN(n15) );
  NAND2X1 U137 ( .IN1(n108), .IN2(n60), .QN(n97) );
  NAND2X0 U138 ( .IN1(n100), .IN2(\input [6]), .QN(n49) );
  NAND2X0 U139 ( .IN1(n101), .IN2(\input [6]), .QN(n65) );
  NAND2X0 U140 ( .IN1(n62), .IN2(\input [6]), .QN(n79) );
  NAND2X0 U141 ( .IN1(n50), .IN2(\input [5]), .QN(n102) );
  NAND2X0 U142 ( .IN1(n44), .IN2(\input [5]), .QN(n38) );
  AO222X1 U143 ( .IN1(\input [2]), .IN2(n100), .IN3(\input [3]), .IN4(n50), 
        .IN5(\input [4]), .IN6(n101), .Q(N16) );
  NAND2X0 U144 ( .IN1(n100), .IN2(\input [4]), .QN(n31) );
  NAND2X0 U145 ( .IN1(n46), .IN2(\input [4]), .QN(n37) );
  NOR2X0 U146 ( .IN1(n95), .IN2(n96), .QN(N17) );
  NOR2X0 U147 ( .IN1(N2), .IN2(n5), .QN(n41) );
  NOR2X0 U148 ( .IN1(n41), .IN2(n42), .QN(n39) );
  INVX0 U149 ( .INP(\input [7]), .ZN(n58) );
  INVX0 U150 ( .INP(\input [5]), .ZN(n68) );
  AO22X2 U151 ( .IN1(N22), .IN2(n118), .IN3(N10), .IN4(n117), .Q(\output [8])
         );
  MUX21X2 U152 ( .IN1(N20), .IN2(N8), .S(n117), .Q(\output [10]) );
  AO22X2 U153 ( .IN1(N16), .IN2(n117), .IN3(N28), .IN4(n118), .Q(\output [2])
         );
  INVX0 U154 ( .INP(n118), .ZN(n117) );
  AO22X1 U155 ( .IN1(N30), .IN2(n118), .IN3(N18), .IN4(n117), .Q(\output [0])
         );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2_DW01_inc_2 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;
  wire   n1, n2, n5, n7, n8, n10, n12, n13, n14, n15, n19, n20, n21, n22, n23,
         n24, n25, n26, n28, n29, n32, n33, n35, n36, n37, n38, n39, n69, n70,
         n71, n72, n73, n74, n75;
  assign n5 = A[11];
  assign n8 = A[10];
  assign n12 = A[9];
  assign n15 = A[8];
  assign n26 = A[5];
  assign n29 = A[4];
  assign n33 = A[3];
  assign n38 = A[1];

  XOR2X1 U1 ( .IN1(n2), .IN2(n1), .Q(SUM[12]) );
  XOR2X1 U13 ( .IN1(n13), .IN2(n14), .Q(SUM[9]) );
  XNOR2X1 U22 ( .IN1(n21), .IN2(n20), .Q(SUM[7]) );
  XOR2X1 U27 ( .IN1(n23), .IN2(n22), .Q(SUM[6]) );
  XNOR2X1 U48 ( .IN1(n39), .IN2(A[0]), .Q(SUM[1]) );
  AND2X1 U54 ( .IN1(n70), .IN2(A[6]), .Q(n21) );
  AND2X1 U55 ( .IN1(n38), .IN2(A[0]), .Q(n69) );
  NOR2X0 U56 ( .IN1(n25), .IN2(n32), .QN(n70) );
  AND4X1 U57 ( .IN1(n12), .IN2(n15), .IN3(n19), .IN4(n70), .Q(n71) );
  AND4X1 U58 ( .IN1(n12), .IN2(n15), .IN3(n19), .IN4(n24), .Q(n10) );
  AND2X1 U59 ( .IN1(n24), .IN2(n19), .Q(n72) );
  AND2X4 U60 ( .IN1(A[2]), .IN2(n74), .Q(n73) );
  AND2X1 U61 ( .IN1(A[6]), .IN2(A[7]), .Q(n19) );
  AND2X1 U62 ( .IN1(n33), .IN2(n69), .Q(n74) );
  AND2X1 U63 ( .IN1(A[2]), .IN2(n69), .Q(n35) );
  XOR2X2 U64 ( .IN1(n36), .IN2(n37), .Q(SUM[2]) );
  NAND2X0 U65 ( .IN1(A[2]), .IN2(n74), .QN(n32) );
  XOR2X1 U66 ( .IN1(n8), .IN2(n71), .Q(SUM[10]) );
  INVX0 U67 ( .INP(n70), .ZN(n23) );
  NAND2X0 U68 ( .IN1(n38), .IN2(A[0]), .QN(n37) );
  INVX0 U69 ( .INP(n38), .ZN(n39) );
  XOR2X1 U70 ( .IN1(n29), .IN2(n73), .Q(SUM[4]) );
  XNOR2X1 U71 ( .IN1(n26), .IN2(n28), .Q(SUM[5]) );
  XNOR2X1 U72 ( .IN1(n7), .IN2(n5), .Q(SUM[11]) );
  AND2X1 U73 ( .IN1(n8), .IN2(n5), .Q(n75) );
  XOR2X1 U74 ( .IN1(n33), .IN2(n35), .Q(SUM[3]) );
  INVX0 U75 ( .INP(n12), .ZN(n13) );
  INVX0 U76 ( .INP(A[6]), .ZN(n22) );
  XOR2X1 U77 ( .IN1(n15), .IN2(n72), .Q(SUM[8]) );
  INVX0 U78 ( .INP(A[7]), .ZN(n20) );
  INVX0 U79 ( .INP(A[12]), .ZN(n1) );
  NAND2X0 U80 ( .IN1(n15), .IN2(n72), .QN(n14) );
  NOR2X0 U81 ( .IN1(n25), .IN2(n32), .QN(n24) );
  NAND2X0 U82 ( .IN1(n75), .IN2(n71), .QN(n2) );
  NAND2X0 U83 ( .IN1(n8), .IN2(n10), .QN(n7) );
  NAND2X0 U84 ( .IN1(n73), .IN2(n29), .QN(n28) );
  NAND2X0 U85 ( .IN1(n26), .IN2(n29), .QN(n25) );
  INVX0 U86 ( .INP(A[2]), .ZN(n36) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2_DW_mult_tc_6 ( a, b, 
        product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n18, n19, n21,
         n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n33, n34, n35, n36,
         n37, n39, n41, n43, n44, n45, n46, n52, n54, n55, n56, n57, n58, n59,
         n60, n61, n63, n64, n65, n68, n69, n70, n74, n75, n76, n77, n78, n79,
         n80, n81, n84, n85, n86, n87, n88, n89, n92, n93, n94, n95, n97, n98,
         n100, n101, n102, n103, n104, n105, n107, n108, n112, n114, n115,
         n116, n120, n121, n125, n127, n128, n129, n130, n131, n132, n134,
         n135, n136, n137, n138, n139, n141, n143, n149, n150, n153, n154,
         n156, n157, n158, n161, n162, n164, n167, n168, n170, n171, n175,
         n176, n177, n178, n180, n181, n183, n184, n185, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962;

  AOI21X1 U6 ( .IN1(n1), .IN2(n21), .IN3(n22), .QN(product[23]) );
  OAI21X1 U8 ( .IN1(n23), .IN2(n639), .IN3(n24), .QN(n22) );
  AOI21X1 U10 ( .IN1(n622), .IN2(n25), .IN3(n26), .QN(n24) );
  OAI21X1 U12 ( .IN1(n27), .IN2(n37), .IN3(n28), .QN(n26) );
  OAI21X1 U20 ( .IN1(n32), .IN2(n2), .IN3(n33), .QN(n31) );
  AOI21X1 U22 ( .IN1(n34), .IN2(n59), .IN3(n35), .QN(n33) );
  AOI21X1 U26 ( .IN1(n692), .IN2(n962), .IN3(n39), .QN(n37) );
  OAI21X1 U36 ( .IN1(n45), .IN2(n639), .IN3(n46), .QN(n44) );
  AOI21X1 U38 ( .IN1(n59), .IN2(n961), .IN3(n692), .QN(n46) );
  OAI21X1 U50 ( .IN1(n56), .IN2(n2), .IN3(n57), .QN(n55) );
  OAI21X1 U54 ( .IN1(n60), .IN2(n68), .IN3(n61), .QN(n59) );
  XOR2X1 U59 ( .IN1(n69), .IN2(n8), .Q(product[18]) );
  OAI21X1 U62 ( .IN1(n65), .IN2(n639), .IN3(n621), .QN(n64) );
  XOR2X1 U69 ( .IN1(n78), .IN2(n9), .Q(product[17]) );
  AOI21X1 U70 ( .IN1(n1), .IN2(n70), .IN3(n797), .QN(n69) );
  AOI21X1 U74 ( .IN1(n74), .IN2(n87), .IN3(n75), .QN(n2) );
  OAI21X1 U76 ( .IN1(n84), .IN2(n76), .IN3(n77), .QN(n75) );
  AOI21X1 U82 ( .IN1(n1), .IN2(n79), .IN3(n80), .QN(n78) );
  OAI21X1 U98 ( .IN1(n98), .IN2(n92), .IN3(n93), .QN(n87) );
  AOI21X1 U104 ( .IN1(n1), .IN2(n95), .IN3(n685), .QN(n94) );
  AOI21X1 U114 ( .IN1(n102), .IN2(n115), .IN3(n103), .QN(n101) );
  OAI21X1 U116 ( .IN1(n112), .IN2(n104), .IN3(n105), .QN(n103) );
  OAI21X1 U124 ( .IN1(n673), .IN2(n785), .IN3(n112), .QN(n108) );
  OAI21X1 U138 ( .IN1(n678), .IN2(n120), .IN3(n121), .QN(n115) );
  AOI21X1 U153 ( .IN1(n137), .IN2(n129), .IN3(n130), .QN(n128) );
  OAI21X1 U155 ( .IN1(n135), .IN2(n131), .IN3(n132), .QN(n130) );
  OAI21X1 U168 ( .IN1(n150), .IN2(n138), .IN3(n139), .QN(n137) );
  AOI21X1 U170 ( .IN1(n949), .IN2(n952), .IN3(n141), .QN(n139) );
  FADDX1 U204 ( .A(n408), .B(n419), .CI(n191), .CO(n187), .S(n188) );
  FADDX1 U205 ( .A(n192), .B(n197), .CI(n195), .CO(n189), .S(n190) );
  FADDX1 U206 ( .A(n431), .B(n420), .CI(n409), .CO(n191), .S(n192) );
  FADDX1 U207 ( .A(n196), .B(n203), .CI(n201), .CO(n193), .S(n194) );
  FADDX1 U208 ( .A(n205), .B(n410), .CI(n198), .CO(n195), .S(n196) );
  FADDX1 U209 ( .A(n421), .B(n432), .CI(n443), .CO(n197), .S(n198) );
  FADDX1 U212 ( .A(n411), .B(n455), .CI(n206), .CO(n203), .S(n204) );
  FADDX1 U213 ( .A(n422), .B(n433), .CI(n444), .CO(n205), .S(n206) );
  FADDX1 U217 ( .A(n456), .B(n467), .CI(n412), .CO(n213), .S(n214) );
  FADDX1 U218 ( .A(n434), .B(n445), .CI(n423), .CO(n215), .S(n216) );
  FADDX1 U221 ( .A(n226), .B(n239), .CI(n237), .CO(n221), .S(n222) );
  FADDX1 U223 ( .A(n435), .B(n457), .CI(n413), .CO(n225), .S(n226) );
  FADDX1 U224 ( .A(n446), .B(n424), .CI(n468), .CO(n227), .S(n228) );
  FADDX1 U230 ( .A(n458), .B(n436), .CI(n447), .CO(n239), .S(n240) );
  FADDX1 U234 ( .A(n267), .B(n269), .CI(n252), .CO(n247), .S(n248) );
  FADDX1 U238 ( .A(n470), .B(n415), .CI(n448), .CO(n255), .S(n256) );
  FADDX1 U251 ( .A(n305), .B(n288), .CI(n286), .CO(n281), .S(n282) );
  FADDX1 U257 ( .A(n439), .B(n505), .CI(n417), .CO(n293), .S(n294) );
  XNOR2X1 U258 ( .IN1(n516), .IN2(n428), .Q(n296) );
  FADDX1 U260 ( .A(n319), .B(n302), .CI(n300), .CO(n297), .S(n298) );
  HADDX1 U269 ( .A0(n528), .B0(n429), .C1(n315), .SO(n316) );
  FADDX1 U275 ( .A(n463), .B(n507), .CI(n334), .CO(n327), .S(n328) );
  HADDX1 U278 ( .A0(n430), .B0(n540), .C1(n333), .SO(n334) );
  FADDX1 U283 ( .A(n486), .B(n497), .CI(n350), .CO(n343), .S(n344) );
  HADDX1 U286 ( .A0(n442), .B0(n541), .C1(n349), .SO(n350) );
  FADDX1 U291 ( .A(n531), .B(n465), .CI(n509), .CO(n359), .S(n360) );
  FADDX1 U295 ( .A(n372), .B(n374), .CI(n381), .CO(n367), .S(n368) );
  FADDX1 U300 ( .A(n382), .B(n389), .CI(n380), .CO(n377), .S(n378) );
  FADDX1 U302 ( .A(n489), .B(n386), .CI(n533), .CO(n381), .S(n382) );
  FADDX1 U303 ( .A(n544), .B(n511), .CI(n478), .CO(n383), .S(n384) );
  HADDX1 U304 ( .A0(n522), .B0(n500), .C1(n385), .SO(n386) );
  FADDX1 U305 ( .A(n392), .B(n397), .CI(n390), .CO(n387), .S(n388) );
  FADDX1 U306 ( .A(n545), .B(n399), .CI(n490), .CO(n389), .S(n390) );
  HADDX1 U308 ( .A0(n501), .B0(n523), .C1(n393), .SO(n394) );
  FADDX1 U309 ( .A(n403), .B(n400), .CI(n398), .CO(n395), .S(n396) );
  FADDX1 U310 ( .A(n535), .B(n502), .CI(n513), .CO(n397), .S(n398) );
  HADDX1 U311 ( .A0(n524), .B0(n546), .C1(n399), .SO(n400) );
  FADDX1 U312 ( .A(n514), .B(n547), .CI(n404), .CO(n401), .S(n402) );
  HADDX1 U313 ( .A0(n525), .B0(n536), .C1(n403), .SO(n404) );
  HADDX1 U314 ( .A0(n548), .B0(n526), .C1(n405), .SO(n406) );
  OR2X1 U323 ( .IN1(n677), .IN2(n558), .Q(n415) );
  OR2X1 U324 ( .IN1(n562), .IN2(n559), .Q(n416) );
  OR2X1 U325 ( .IN1(n560), .IN2(n677), .Q(n417) );
  OR2X1 U326 ( .IN1(n562), .IN2(n561), .Q(n418) );
  OR2X1 U327 ( .IN1(n550), .IN2(n705), .Q(n419) );
  OR2X1 U363 ( .IN1(n714), .IN2(n550), .Q(n455) );
  OR2X1 U411 ( .IN1(n550), .IN2(n570), .Q(n503) );
  OR2X1 U423 ( .IN1(n571), .IN2(n550), .Q(n515) );
  OR2X1 U435 ( .IN1(n550), .IN2(n572), .Q(n527) );
  NAND3X0 U484 ( .IN1(n787), .IN2(n789), .IN3(n788), .QN(n619) );
  INVX0 U485 ( .INP(n68), .ZN(n620) );
  INVX0 U486 ( .INP(n620), .ZN(n621) );
  NAND3X1 U487 ( .IN1(n944), .IN2(n945), .IN3(n946), .QN(n245) );
  AND2X4 U488 ( .IN1(a[6]), .IN2(n676), .Q(n468) );
  OAI21X1 U489 ( .IN1(n60), .IN2(n68), .IN3(n61), .QN(n622) );
  NAND3X0 U490 ( .IN1(n944), .IN2(n945), .IN3(n946), .QN(n623) );
  NAND3X0 U491 ( .IN1(n848), .IN2(n849), .IN3(n696), .QN(n709) );
  NAND3X4 U492 ( .IN1(n902), .IN2(n903), .IN3(n904), .QN(n798) );
  INVX0 U493 ( .INP(n306), .ZN(n624) );
  INVX0 U494 ( .INP(n624), .ZN(n625) );
  NAND2X0 U495 ( .IN1(n315), .IN2(n296), .QN(n750) );
  NAND2X0 U496 ( .IN1(n313), .IN2(n315), .QN(n752) );
  XOR2X2 U497 ( .IN1(n796), .IN2(n257), .Q(n238) );
  AND2X1 U498 ( .IN1(n676), .IN2(n707), .Q(n528) );
  AND3X4 U499 ( .IN1(n928), .IN2(n927), .IN3(n929), .Q(n670) );
  XNOR3X1 U500 ( .IN1(n311), .IN2(n626), .IN3(n294), .Q(n286) );
  XNOR3X1 U501 ( .IN1(n450), .IN2(n527), .IN3(n494), .Q(n626) );
  INVX0 U502 ( .INP(n551), .ZN(n627) );
  INVX0 U503 ( .INP(n627), .ZN(n628) );
  INVX0 U504 ( .INP(n636), .ZN(n629) );
  NAND3X2 U505 ( .IN1(n888), .IN2(n890), .IN3(n889), .QN(n331) );
  NAND3X1 U506 ( .IN1(n918), .IN2(n916), .IN3(n917), .QN(n683) );
  INVX0 U507 ( .INP(n694), .ZN(n630) );
  XOR2X1 U508 ( .IN1(n337), .IN2(n322), .Q(n631) );
  XOR2X1 U509 ( .IN1(n631), .IN2(n320), .Q(n318) );
  NAND2X0 U510 ( .IN1(n322), .IN2(n320), .QN(n632) );
  NAND2X0 U511 ( .IN1(n337), .IN2(n320), .QN(n633) );
  NAND2X0 U512 ( .IN1(n337), .IN2(n322), .QN(n634) );
  NAND3X0 U513 ( .IN1(n632), .IN2(n634), .IN3(n633), .QN(n317) );
  NAND3X1 U514 ( .IN1(n851), .IN2(n853), .IN3(n852), .QN(n337) );
  XOR2X2 U515 ( .IN1(n943), .IN2(n263), .Q(n246) );
  NAND2X0 U516 ( .IN1(n515), .IN2(n493), .QN(n759) );
  NAND2X0 U517 ( .IN1(n515), .IN2(n416), .QN(n758) );
  INVX0 U518 ( .INP(b[0]), .ZN(n561) );
  NAND3X0 U519 ( .IN1(n870), .IN2(n871), .IN3(n872), .QN(n309) );
  NAND3X0 U520 ( .IN1(n743), .IN2(n744), .IN3(n745), .QN(n271) );
  OR2X1 U521 ( .IN1(n772), .IN2(n550), .Q(n479) );
  NAND3X0 U522 ( .IN1(n809), .IN2(n810), .IN3(n811), .QN(n373) );
  OR2X1 U523 ( .IN1(n556), .IN2(n677), .Q(n413) );
  XOR2X1 U524 ( .IN1(n821), .IN2(n369), .Q(n354) );
  NAND3X0 U525 ( .IN1(n933), .IN2(n934), .IN3(n935), .QN(n329) );
  XOR3X1 U526 ( .IN1(n518), .IN2(n441), .IN3(n529), .Q(n332) );
  OR2X1 U527 ( .IN1(n555), .IN2(n677), .Q(n412) );
  OAI21X1 U528 ( .IN1(n776), .IN2(n89), .IN3(n640), .QN(n80) );
  INVX0 U529 ( .INP(n27), .ZN(n171) );
  AOI21X1 U530 ( .IN1(n1), .IN2(n86), .IN3(n722), .QN(n85) );
  XNOR2X1 U531 ( .IN1(n861), .IN2(n14), .Q(product[12]) );
  INVX0 U532 ( .INP(n150), .ZN(n149) );
  AND2X4 U533 ( .IN1(n318), .IN2(n335), .Q(n635) );
  INVX0 U534 ( .INP(n560), .ZN(n636) );
  INVX0 U535 ( .INP(n636), .ZN(n637) );
  NAND2X0 U536 ( .IN1(n86), .IN2(n641), .QN(n638) );
  AOI21X1 U537 ( .IN1(n74), .IN2(n87), .IN3(n75), .QN(n639) );
  DELLN1X2 U538 ( .INP(n84), .Z(n640) );
  AND2X4 U539 ( .IN1(a[10]), .IN2(b[0]), .Q(n430) );
  XOR2X1 U540 ( .IN1(n370), .IN2(n379), .Q(n838) );
  NOR2X0 U541 ( .IN1(n820), .IN2(n81), .QN(n641) );
  XOR2X2 U542 ( .IN1(n746), .IN2(n271), .Q(n642) );
  NAND2X0 U543 ( .IN1(n328), .IN2(n326), .QN(n643) );
  XOR2X1 U544 ( .IN1(n866), .IN2(n280), .Q(n278) );
  INVX0 U545 ( .INP(n128), .ZN(n644) );
  NAND2X0 U546 ( .IN1(n425), .IN2(n480), .QN(n907) );
  AND2X1 U547 ( .IN1(n713), .IN2(n715), .Q(n460) );
  XNOR3X1 U548 ( .IN1(n645), .IN2(n248), .IN3(n246), .Q(n244) );
  AND3X1 U549 ( .IN1(n918), .IN2(n916), .IN3(n917), .Q(n645) );
  INVX0 U550 ( .INP(n676), .ZN(n646) );
  XOR2X1 U551 ( .IN1(n236), .IN2(n249), .Q(n898) );
  NAND2X0 U552 ( .IN1(n370), .IN2(n368), .QN(n840) );
  XOR3X1 U553 ( .IN1(n450), .IN2(n527), .IN3(n494), .Q(n647) );
  NAND2X0 U554 ( .IN1(n343), .IN2(n326), .QN(n648) );
  XOR2X1 U555 ( .IN1(n887), .IN2(n332), .Q(n326) );
  DELLN1X2 U556 ( .INP(n143), .Z(n649) );
  NOR2X0 U557 ( .IN1(n260), .IN2(n277), .QN(n650) );
  NOR2X0 U558 ( .IN1(n564), .IN2(n703), .QN(n651) );
  XOR3X1 U559 ( .IN1(n655), .IN2(n487), .IN3(n364), .Q(n358) );
  NAND2X0 U560 ( .IN1(n364), .IN2(n375), .QN(n652) );
  NAND2X0 U561 ( .IN1(n487), .IN2(n375), .QN(n653) );
  NAND2X0 U562 ( .IN1(n487), .IN2(n364), .QN(n654) );
  NAND3X0 U563 ( .IN1(n652), .IN2(n654), .IN3(n653), .QN(n357) );
  AND2X1 U564 ( .IN1(n510), .IN2(n499), .Q(n655) );
  XOR2X2 U565 ( .IN1(n359), .IN2(n357), .Q(n844) );
  HADDX1 U566 ( .A0(n498), .B0(n454), .C1(n363), .SO(n364) );
  XOR3X1 U567 ( .IN1(n210), .IN2(n221), .IN3(n219), .Q(n208) );
  NAND2X0 U568 ( .IN1(n219), .IN2(n210), .QN(n656) );
  NAND2X0 U569 ( .IN1(n221), .IN2(n210), .QN(n657) );
  NAND2X0 U570 ( .IN1(n221), .IN2(n219), .QN(n658) );
  NAND3X0 U571 ( .IN1(n656), .IN2(n658), .IN3(n657), .QN(n207) );
  INVX0 U572 ( .INP(a[1]), .ZN(n659) );
  XOR2X2 U573 ( .IN1(n953), .IN2(n954), .Q(product[20]) );
  XOR2X1 U574 ( .IN1(n314), .IN2(n681), .Q(n936) );
  XOR3X1 U575 ( .IN1(n213), .IN2(n215), .IN3(n204), .Q(n202) );
  XOR2X1 U576 ( .IN1(n211), .IN2(n209), .Q(n660) );
  XOR2X2 U577 ( .IN1(n660), .IN2(n202), .Q(n200) );
  NAND2X1 U578 ( .IN1(n213), .IN2(n215), .QN(n661) );
  NAND2X0 U579 ( .IN1(n213), .IN2(n204), .QN(n662) );
  NAND2X0 U580 ( .IN1(n215), .IN2(n204), .QN(n663) );
  NAND3X0 U581 ( .IN1(n661), .IN2(n662), .IN3(n663), .QN(n201) );
  NAND2X0 U582 ( .IN1(n211), .IN2(n209), .QN(n664) );
  NAND2X0 U583 ( .IN1(n211), .IN2(n202), .QN(n665) );
  NAND2X0 U584 ( .IN1(n209), .IN2(n202), .QN(n666) );
  NAND3X0 U585 ( .IN1(n664), .IN2(n665), .IN3(n666), .QN(n199) );
  XOR3X1 U586 ( .IN1(n327), .IN2(n312), .IN3(n310), .Q(n304) );
  NAND2X0 U587 ( .IN1(n310), .IN2(n327), .QN(n667) );
  NAND2X0 U588 ( .IN1(n312), .IN2(n327), .QN(n668) );
  NAND2X0 U589 ( .IN1(n312), .IN2(n310), .QN(n669) );
  NAND3X0 U590 ( .IN1(n667), .IN2(n669), .IN3(n668), .QN(n303) );
  XOR2X2 U591 ( .IN1(n284), .IN2(n303), .Q(n926) );
  AO21X1 U592 ( .IN1(n54), .IN2(n922), .IN3(n55), .Q(n953) );
  XOR2X2 U593 ( .IN1(n85), .IN2(n10), .Q(product[16]) );
  NAND3X0 U594 ( .IN1(n884), .IN2(n886), .IN3(n885), .QN(n671) );
  INVX0 U595 ( .INP(a[3]), .ZN(n672) );
  NOR2X0 U596 ( .IN1(n278), .IN2(n297), .QN(n673) );
  INVX0 U597 ( .INP(n685), .ZN(n674) );
  XOR2X2 U598 ( .IN1(n94), .IN2(n11), .Q(product[15]) );
  INVX0 U599 ( .INP(b[9]), .ZN(n675) );
  INVX0 U600 ( .INP(n551), .ZN(n676) );
  INVX0 U601 ( .INP(a[11]), .ZN(n677) );
  NAND2X0 U602 ( .IN1(n318), .IN2(n335), .QN(n678) );
  INVX0 U603 ( .INP(n713), .ZN(n679) );
  OR2X1 U604 ( .IN1(n199), .IN2(n194), .Q(n680) );
  NAND3X0 U605 ( .IN1(n890), .IN2(n889), .IN3(n888), .QN(n681) );
  INVX0 U606 ( .INP(b[3]), .ZN(n682) );
  INVX0 U607 ( .INP(b[2]), .ZN(n684) );
  AND2X4 U608 ( .IN1(n244), .IN2(n259), .Q(n685) );
  INVX0 U609 ( .INP(b[5]), .ZN(n686) );
  INVX0 U610 ( .INP(n700), .ZN(n687) );
  INVX0 U611 ( .INP(n698), .ZN(n688) );
  INVX0 U612 ( .INP(n450), .ZN(n689) );
  INVX0 U613 ( .INP(n689), .ZN(n690) );
  NOR2X0 U614 ( .IN1(n243), .IN2(n230), .QN(n691) );
  AND2X1 U615 ( .IN1(n193), .IN2(n190), .Q(n692) );
  NAND2X0 U616 ( .IN1(n517), .IN2(n440), .QN(n817) );
  INVX0 U617 ( .INP(n670), .ZN(n693) );
  OR2X1 U618 ( .IN1(n557), .IN2(n677), .Q(n414) );
  INVX0 U619 ( .INP(n564), .ZN(n694) );
  INVX0 U620 ( .INP(n694), .ZN(n695) );
  NAND2X0 U621 ( .IN1(n346), .IN2(n357), .QN(n696) );
  INVX0 U622 ( .INP(n704), .ZN(n697) );
  INVX0 U623 ( .INP(n571), .ZN(n698) );
  INVX0 U624 ( .INP(n698), .ZN(n699) );
  INVX0 U625 ( .INP(n551), .ZN(n700) );
  INVX0 U626 ( .INP(n700), .ZN(n701) );
  NOR2X0 U627 ( .IN1(n298), .IN2(n317), .QN(n702) );
  INVX0 U628 ( .INP(b[4]), .ZN(n703) );
  INVX0 U629 ( .INP(n563), .ZN(n704) );
  INVX0 U630 ( .INP(n704), .ZN(n705) );
  INVX0 U631 ( .INP(n707), .ZN(n706) );
  INVX0 U632 ( .INP(n572), .ZN(n707) );
  INVX0 U633 ( .INP(n707), .ZN(n708) );
  INVX0 U634 ( .INP(b[6]), .ZN(n710) );
  INVX0 U635 ( .INP(a[4]), .ZN(n711) );
  INVX0 U636 ( .INP(a[6]), .ZN(n712) );
  INVX0 U637 ( .INP(n566), .ZN(n713) );
  INVX0 U638 ( .INP(n713), .ZN(n714) );
  INVX0 U639 ( .INP(n555), .ZN(n715) );
  NAND2X0 U640 ( .IN1(n479), .IN2(n228), .QN(n792) );
  XOR2X2 U641 ( .IN1(n256), .IN2(n254), .Q(n746) );
  XOR3X1 U642 ( .IN1(n459), .IN2(n481), .IN3(n437), .Q(n254) );
  NAND2X1 U643 ( .IN1(n437), .IN2(n459), .QN(n716) );
  NAND2X0 U644 ( .IN1(n481), .IN2(n459), .QN(n717) );
  NAND2X0 U645 ( .IN1(n481), .IN2(n437), .QN(n718) );
  NAND3X0 U646 ( .IN1(n716), .IN2(n718), .IN3(n717), .QN(n253) );
  INVX0 U647 ( .INP(n301), .ZN(n719) );
  INVX0 U648 ( .INP(n719), .ZN(n720) );
  INVX0 U649 ( .INP(b[7]), .ZN(n721) );
  INVX0 U650 ( .INP(n89), .ZN(n722) );
  XOR2X1 U651 ( .IN1(n273), .IN2(n275), .Q(n723) );
  XOR2X1 U652 ( .IN1(n723), .IN2(n258), .Q(n252) );
  NAND2X0 U653 ( .IN1(n275), .IN2(n258), .QN(n724) );
  NAND2X0 U654 ( .IN1(n273), .IN2(n258), .QN(n725) );
  NAND2X1 U655 ( .IN1(n273), .IN2(n275), .QN(n726) );
  NAND3X0 U656 ( .IN1(n724), .IN2(n726), .IN3(n725), .QN(n251) );
  XOR3X1 U657 ( .IN1(n492), .IN2(n503), .IN3(n426), .Q(n258) );
  NAND2X0 U658 ( .IN1(n426), .IN2(n492), .QN(n727) );
  NAND2X0 U659 ( .IN1(n503), .IN2(n492), .QN(n728) );
  NAND2X0 U660 ( .IN1(n503), .IN2(n426), .QN(n729) );
  NAND3X0 U661 ( .IN1(n727), .IN2(n729), .IN3(n728), .QN(n257) );
  XOR2X2 U662 ( .IN1(n926), .IN2(n720), .Q(n280) );
  NAND2X0 U663 ( .IN1(n418), .IN2(n440), .QN(n819) );
  XOR2X1 U664 ( .IN1(n482), .IN2(n449), .Q(n730) );
  XOR2X1 U665 ( .IN1(n730), .IN2(n293), .Q(n270) );
  NAND2X0 U666 ( .IN1(n449), .IN2(n293), .QN(n731) );
  NAND2X0 U667 ( .IN1(n482), .IN2(n293), .QN(n732) );
  NAND2X1 U668 ( .IN1(n482), .IN2(n449), .QN(n733) );
  NAND3X0 U669 ( .IN1(n731), .IN2(n733), .IN3(n732), .QN(n269) );
  XOR3X1 U670 ( .IN1(n354), .IN2(n356), .IN3(n367), .Q(n352) );
  NAND2X1 U671 ( .IN1(n367), .IN2(n356), .QN(n734) );
  NAND2X0 U672 ( .IN1(n354), .IN2(n356), .QN(n735) );
  NAND2X0 U673 ( .IN1(n354), .IN2(n367), .QN(n736) );
  NAND3X0 U674 ( .IN1(n734), .IN2(n736), .IN3(n735), .QN(n351) );
  XOR3X1 U675 ( .IN1(n521), .IN2(n376), .IN3(n466), .Q(n372) );
  NAND2X0 U676 ( .IN1(n466), .IN2(n521), .QN(n737) );
  NAND2X0 U677 ( .IN1(n376), .IN2(n521), .QN(n738) );
  NAND2X0 U678 ( .IN1(n376), .IN2(n466), .QN(n739) );
  NAND3X0 U679 ( .IN1(n737), .IN2(n739), .IN3(n738), .QN(n371) );
  XOR2X1 U680 ( .IN1(n812), .IN2(n373), .Q(n356) );
  HADDX1 U681 ( .A0(n510), .B0(n499), .C1(n375), .SO(n376) );
  XOR2X2 U682 ( .IN1(n362), .IN2(n371), .Q(n812) );
  XNOR2X2 U683 ( .IN1(n127), .IN2(n16), .Q(product[10]) );
  XOR3X1 U684 ( .IN1(n472), .IN2(n483), .IN3(n461), .Q(n290) );
  NAND2X0 U685 ( .IN1(n461), .IN2(n472), .QN(n740) );
  NAND2X0 U686 ( .IN1(n483), .IN2(n472), .QN(n741) );
  NAND2X0 U687 ( .IN1(n483), .IN2(n461), .QN(n742) );
  NAND3X0 U688 ( .IN1(n740), .IN2(n742), .IN3(n741), .QN(n289) );
  XOR3X1 U689 ( .IN1(n460), .IN2(n471), .IN3(n295), .Q(n272) );
  NAND2X0 U690 ( .IN1(n460), .IN2(n471), .QN(n743) );
  NAND2X1 U691 ( .IN1(n460), .IN2(n295), .QN(n744) );
  NAND2X0 U692 ( .IN1(n471), .IN2(n295), .QN(n745) );
  XOR2X2 U693 ( .IN1(n746), .IN2(n271), .Q(n250) );
  NAND2X0 U694 ( .IN1(n256), .IN2(n254), .QN(n747) );
  NAND2X0 U695 ( .IN1(n256), .IN2(n271), .QN(n748) );
  NAND2X0 U696 ( .IN1(n254), .IN2(n271), .QN(n749) );
  NAND3X0 U697 ( .IN1(n747), .IN2(n748), .IN3(n749), .QN(n249) );
  XNOR2X2 U698 ( .IN1(n862), .IN2(n15), .Q(product[11]) );
  XOR3X1 U699 ( .IN1(n296), .IN2(n313), .IN3(n315), .Q(n288) );
  NAND2X1 U700 ( .IN1(n313), .IN2(n296), .QN(n751) );
  NAND3X0 U701 ( .IN1(n750), .IN2(n752), .IN3(n751), .QN(n287) );
  XOR3X1 U702 ( .IN1(n285), .IN2(n287), .IN3(n268), .Q(n264) );
  OR2X4 U703 ( .IN1(n675), .IN2(n677), .Q(n409) );
  XNOR2X2 U704 ( .IN1(n1), .IN2(n12), .Q(product[14]) );
  INVX0 U705 ( .INP(a[8]), .ZN(n753) );
  XOR3X1 U706 ( .IN1(n473), .IN2(n333), .IN3(n484), .Q(n308) );
  NAND2X1 U707 ( .IN1(n484), .IN2(n473), .QN(n754) );
  NAND2X0 U708 ( .IN1(n333), .IN2(n473), .QN(n755) );
  NAND2X0 U709 ( .IN1(n333), .IN2(n484), .QN(n756) );
  NAND3X0 U710 ( .IN1(n754), .IN2(n756), .IN3(n755), .QN(n307) );
  XOR3X1 U711 ( .IN1(n416), .IN2(n515), .IN3(n493), .Q(n274) );
  NAND2X1 U712 ( .IN1(n493), .IN2(n416), .QN(n757) );
  NAND3X0 U713 ( .IN1(n757), .IN2(n759), .IN3(n758), .QN(n273) );
  OR2X4 U714 ( .IN1(n677), .IN2(n701), .Q(n408) );
  XOR2X1 U715 ( .IN1(n838), .IN2(n368), .Q(n366) );
  XOR3X1 U716 ( .IN1(n338), .IN2(n340), .IN3(n353), .Q(n336) );
  NAND2X1 U717 ( .IN1(n353), .IN2(n340), .QN(n760) );
  NAND2X0 U718 ( .IN1(n338), .IN2(n340), .QN(n761) );
  NAND2X0 U719 ( .IN1(n338), .IN2(n353), .QN(n762) );
  NAND3X0 U720 ( .IN1(n760), .IN2(n762), .IN3(n761), .QN(n335) );
  XOR2X1 U721 ( .IN1(n844), .IN2(n346), .Q(n340) );
  XOR2X1 U722 ( .IN1(n850), .IN2(n355), .Q(n338) );
  OR2X1 U723 ( .IN1(n550), .IN2(n711), .Q(n491) );
  XOR3X1 U724 ( .IN1(n453), .IN2(n475), .IN3(n530), .Q(n348) );
  NAND2X0 U725 ( .IN1(n475), .IN2(n530), .QN(n763) );
  NAND2X0 U726 ( .IN1(n453), .IN2(n530), .QN(n764) );
  NAND2X0 U727 ( .IN1(n453), .IN2(n475), .QN(n765) );
  NAND3X0 U728 ( .IN1(n763), .IN2(n765), .IN3(n764), .QN(n347) );
  INVX0 U729 ( .INP(b[8]), .ZN(n766) );
  INVX0 U730 ( .INP(b[8]), .ZN(n767) );
  XOR2X1 U731 ( .IN1(n488), .IN2(n385), .Q(n768) );
  XOR2X1 U732 ( .IN1(n768), .IN2(n383), .Q(n370) );
  NAND2X0 U733 ( .IN1(n385), .IN2(n383), .QN(n769) );
  NAND2X0 U734 ( .IN1(n488), .IN2(n383), .QN(n770) );
  NAND2X1 U735 ( .IN1(n488), .IN2(n385), .QN(n771) );
  NAND3X0 U736 ( .IN1(n769), .IN2(n771), .IN3(n770), .QN(n369) );
  INVX0 U737 ( .INP(a[5]), .ZN(n772) );
  OR2X4 U738 ( .IN1(n516), .IN2(n428), .Q(n295) );
  XOR2X2 U739 ( .IN1(n842), .IN2(n947), .Q(product[9]) );
  XOR3X1 U740 ( .IN1(n427), .IN2(n651), .IN3(n504), .Q(n276) );
  NAND2X1 U741 ( .IN1(n504), .IN2(n427), .QN(n773) );
  NAND2X0 U742 ( .IN1(n651), .IN2(n427), .QN(n774) );
  NAND2X0 U743 ( .IN1(n651), .IN2(n504), .QN(n775) );
  NAND3X0 U744 ( .IN1(n773), .IN2(n775), .IN3(n774), .QN(n275) );
  XOR2X1 U745 ( .IN1(n276), .IN2(n274), .Q(n857) );
  INVX0 U746 ( .INP(n177), .ZN(n776) );
  XOR3X1 U747 ( .IN1(n216), .IN2(n227), .IN3(n214), .Q(n212) );
  XOR2X2 U748 ( .IN1(n223), .IN2(n225), .Q(n777) );
  XOR2X2 U749 ( .IN1(n777), .IN2(n212), .Q(n210) );
  NAND2X0 U750 ( .IN1(n216), .IN2(n227), .QN(n778) );
  NAND2X0 U751 ( .IN1(n216), .IN2(n214), .QN(n779) );
  NAND2X0 U752 ( .IN1(n227), .IN2(n214), .QN(n780) );
  NAND3X0 U753 ( .IN1(n778), .IN2(n779), .IN3(n780), .QN(n211) );
  NAND2X0 U754 ( .IN1(n223), .IN2(n225), .QN(n781) );
  NAND2X0 U755 ( .IN1(n223), .IN2(n212), .QN(n782) );
  NAND2X0 U756 ( .IN1(n225), .IN2(n212), .QN(n783) );
  NAND3X0 U757 ( .IN1(n781), .IN2(n782), .IN3(n783), .QN(n209) );
  INVX0 U758 ( .INP(a[8]), .ZN(n784) );
  XOR2X2 U759 ( .IN1(n957), .IN2(n958), .Q(product[21]) );
  OA21X1 U760 ( .IN1(n678), .IN2(n702), .IN3(n121), .Q(n785) );
  XOR2X1 U761 ( .IN1(n289), .IN2(n272), .Q(n786) );
  XOR2X2 U762 ( .IN1(n786), .IN2(n270), .Q(n266) );
  NAND2X0 U763 ( .IN1(n272), .IN2(n270), .QN(n787) );
  NAND2X0 U764 ( .IN1(n289), .IN2(n270), .QN(n788) );
  NAND2X0 U765 ( .IN1(n289), .IN2(n272), .QN(n789) );
  NAND3X0 U766 ( .IN1(n787), .IN2(n789), .IN3(n788), .QN(n265) );
  XOR2X1 U767 ( .IN1(n265), .IN2(n250), .Q(n943) );
  XOR3X1 U768 ( .IN1(n241), .IN2(n479), .IN3(n228), .Q(n224) );
  NAND2X0 U769 ( .IN1(n228), .IN2(n241), .QN(n790) );
  NAND2X0 U770 ( .IN1(n479), .IN2(n241), .QN(n791) );
  NAND3X0 U771 ( .IN1(n790), .IN2(n792), .IN3(n791), .QN(n223) );
  XOR3X1 U772 ( .IN1(n469), .IN2(n414), .IN3(n491), .Q(n242) );
  NAND2X0 U773 ( .IN1(n491), .IN2(n469), .QN(n793) );
  NAND2X0 U774 ( .IN1(n414), .IN2(n469), .QN(n794) );
  NAND2X1 U775 ( .IN1(n414), .IN2(n491), .QN(n795) );
  NAND3X0 U776 ( .IN1(n793), .IN2(n795), .IN3(n794), .QN(n241) );
  XOR3X1 U777 ( .IN1(n266), .IN2(n283), .IN3(n281), .Q(n262) );
  XOR2X1 U778 ( .IN1(n480), .IN2(n425), .Q(n796) );
  AO21X1 U779 ( .IN1(n641), .IN2(n722), .IN3(n75), .Q(n797) );
  XOR3X1 U780 ( .IN1(n391), .IN2(n393), .IN3(n384), .Q(n380) );
  NAND2X0 U781 ( .IN1(n384), .IN2(n391), .QN(n799) );
  NAND2X0 U782 ( .IN1(n393), .IN2(n391), .QN(n800) );
  NAND2X0 U783 ( .IN1(n393), .IN2(n384), .QN(n801) );
  NAND3X0 U784 ( .IN1(n799), .IN2(n801), .IN3(n800), .QN(n379) );
  XOR2X1 U785 ( .IN1(n512), .IN2(n534), .Q(n802) );
  XOR2X1 U786 ( .IN1(n802), .IN2(n394), .Q(n392) );
  NAND2X0 U787 ( .IN1(n534), .IN2(n394), .QN(n803) );
  NAND2X0 U788 ( .IN1(n512), .IN2(n394), .QN(n804) );
  NAND2X0 U789 ( .IN1(n512), .IN2(n534), .QN(n805) );
  NAND3X0 U790 ( .IN1(n803), .IN2(n805), .IN3(n804), .QN(n391) );
  NAND2X0 U791 ( .IN1(n248), .IN2(n246), .QN(n932) );
  XOR3X1 U792 ( .IN1(n542), .IN2(n476), .IN3(n520), .Q(n362) );
  NAND2X0 U793 ( .IN1(n520), .IN2(n476), .QN(n806) );
  NAND2X0 U794 ( .IN1(n542), .IN2(n476), .QN(n807) );
  NAND2X0 U795 ( .IN1(n542), .IN2(n520), .QN(n808) );
  NAND3X0 U796 ( .IN1(n806), .IN2(n808), .IN3(n807), .QN(n361) );
  XOR3X1 U797 ( .IN1(n543), .IN2(n532), .IN3(n477), .Q(n374) );
  NAND2X0 U798 ( .IN1(n477), .IN2(n532), .QN(n809) );
  NAND2X0 U799 ( .IN1(n477), .IN2(n543), .QN(n810) );
  NAND2X1 U800 ( .IN1(n532), .IN2(n543), .QN(n811) );
  NAND2X0 U801 ( .IN1(n362), .IN2(n371), .QN(n813) );
  NAND2X0 U802 ( .IN1(n362), .IN2(n373), .QN(n814) );
  NAND2X0 U803 ( .IN1(n371), .IN2(n373), .QN(n815) );
  NAND3X0 U804 ( .IN1(n813), .IN2(n814), .IN3(n815), .QN(n355) );
  OR2X1 U805 ( .IN1(n298), .IN2(n317), .Q(n816) );
  XOR3X1 U806 ( .IN1(n517), .IN2(n418), .IN3(n440), .Q(n314) );
  NAND2X0 U807 ( .IN1(n418), .IN2(n517), .QN(n818) );
  NAND3X0 U808 ( .IN1(n817), .IN2(n819), .IN3(n818), .QN(n313) );
  NOR2X0 U809 ( .IN1(n217), .IN2(n208), .QN(n820) );
  XOR2X1 U810 ( .IN1(n360), .IN2(n358), .Q(n821) );
  NAND2X0 U811 ( .IN1(n358), .IN2(n369), .QN(n822) );
  NAND2X0 U812 ( .IN1(n360), .IN2(n369), .QN(n823) );
  NAND2X0 U813 ( .IN1(n360), .IN2(n358), .QN(n824) );
  NAND3X0 U814 ( .IN1(n822), .IN2(n824), .IN3(n823), .QN(n353) );
  XOR3X1 U815 ( .IN1(n623), .IN2(n247), .IN3(n232), .Q(n230) );
  NAND2X0 U816 ( .IN1(n232), .IN2(n245), .QN(n825) );
  NAND2X0 U817 ( .IN1(n247), .IN2(n245), .QN(n826) );
  NAND2X0 U818 ( .IN1(n247), .IN2(n232), .QN(n827) );
  NAND3X0 U819 ( .IN1(n825), .IN2(n827), .IN3(n826), .QN(n229) );
  XOR2X1 U820 ( .IN1(n898), .IN2(n234), .Q(n232) );
  XOR3X1 U821 ( .IN1(n235), .IN2(n224), .IN3(n222), .Q(n220) );
  XOR2X1 U822 ( .IN1(n233), .IN2(n231), .Q(n828) );
  XOR2X2 U823 ( .IN1(n828), .IN2(n220), .Q(n218) );
  NAND2X0 U824 ( .IN1(n235), .IN2(n224), .QN(n829) );
  NAND2X0 U825 ( .IN1(n235), .IN2(n222), .QN(n830) );
  NAND2X0 U826 ( .IN1(n224), .IN2(n222), .QN(n831) );
  NAND3X0 U827 ( .IN1(n829), .IN2(n830), .IN3(n831), .QN(n219) );
  NAND2X0 U828 ( .IN1(n233), .IN2(n798), .QN(n832) );
  NAND2X0 U829 ( .IN1(n233), .IN2(n220), .QN(n833) );
  NAND2X0 U830 ( .IN1(n798), .IN2(n220), .QN(n834) );
  NAND3X0 U831 ( .IN1(n832), .IN2(n833), .IN3(n834), .QN(n217) );
  XOR3X1 U832 ( .IN1(n255), .IN2(n242), .IN3(n240), .Q(n236) );
  NAND2X1 U833 ( .IN1(n242), .IN2(n255), .QN(n835) );
  NAND2X0 U834 ( .IN1(n240), .IN2(n255), .QN(n836) );
  NAND2X0 U835 ( .IN1(n240), .IN2(n242), .QN(n837) );
  NAND3X0 U836 ( .IN1(n835), .IN2(n837), .IN3(n836), .QN(n235) );
  NAND2X0 U837 ( .IN1(n379), .IN2(n368), .QN(n839) );
  NAND2X0 U838 ( .IN1(n370), .IN2(n379), .QN(n841) );
  NAND3X0 U839 ( .IN1(n839), .IN2(n841), .IN3(n840), .QN(n365) );
  OA21X1 U840 ( .IN1(n134), .IN2(n136), .IN3(n135), .Q(n842) );
  XOR3X1 U841 ( .IN1(n361), .IN2(n363), .IN3(n348), .Q(n843) );
  XOR2X2 U842 ( .IN1(n136), .IN2(n18), .Q(product[8]) );
  XOR3X1 U843 ( .IN1(n519), .IN2(n508), .IN3(n464), .Q(n346) );
  NAND2X0 U844 ( .IN1(n519), .IN2(n508), .QN(n845) );
  NAND2X0 U845 ( .IN1(n519), .IN2(n464), .QN(n846) );
  NAND2X0 U846 ( .IN1(n508), .IN2(n464), .QN(n847) );
  NAND3X0 U847 ( .IN1(n845), .IN2(n846), .IN3(n847), .QN(n345) );
  NAND2X0 U848 ( .IN1(n359), .IN2(n357), .QN(n848) );
  NAND2X0 U849 ( .IN1(n359), .IN2(n346), .QN(n849) );
  NAND3X0 U850 ( .IN1(n849), .IN2(n696), .IN3(n848), .QN(n339) );
  XOR2X1 U851 ( .IN1(n344), .IN2(n342), .Q(n850) );
  NAND2X0 U852 ( .IN1(n843), .IN2(n355), .QN(n851) );
  NAND2X0 U853 ( .IN1(n344), .IN2(n355), .QN(n852) );
  NAND2X0 U854 ( .IN1(n344), .IN2(n843), .QN(n853) );
  NAND2X0 U855 ( .IN1(n690), .IN2(n527), .QN(n854) );
  NAND2X0 U856 ( .IN1(n690), .IN2(n494), .QN(n855) );
  NAND2X1 U857 ( .IN1(n527), .IN2(n494), .QN(n856) );
  NAND3X0 U858 ( .IN1(n854), .IN2(n855), .IN3(n856), .QN(n291) );
  XOR2X2 U859 ( .IN1(n857), .IN2(n291), .Q(n268) );
  NAND2X0 U860 ( .IN1(n276), .IN2(n274), .QN(n858) );
  NAND2X0 U861 ( .IN1(n276), .IN2(n291), .QN(n859) );
  NAND2X0 U862 ( .IN1(n274), .IN2(n291), .QN(n860) );
  NAND3X0 U863 ( .IN1(n858), .IN2(n859), .IN3(n860), .QN(n267) );
  AO21X1 U864 ( .IN1(n127), .IN2(n114), .IN3(n115), .Q(n861) );
  AO21X1 U865 ( .IN1(n644), .IN2(n183), .IN3(n635), .Q(n862) );
  XOR3X1 U866 ( .IN1(n347), .IN2(n330), .IN3(n345), .Q(n324) );
  NAND2X0 U867 ( .IN1(n345), .IN2(n347), .QN(n863) );
  NAND2X0 U868 ( .IN1(n330), .IN2(n347), .QN(n864) );
  NAND2X1 U869 ( .IN1(n330), .IN2(n345), .QN(n865) );
  NAND3X0 U870 ( .IN1(n863), .IN2(n865), .IN3(n864), .QN(n323) );
  NAND2X0 U871 ( .IN1(n323), .IN2(n304), .QN(n897) );
  XOR2X1 U872 ( .IN1(n324), .IN2(n339), .Q(n911) );
  XOR2X1 U873 ( .IN1(n282), .IN2(n299), .Q(n866) );
  NAND2X0 U874 ( .IN1(n299), .IN2(n280), .QN(n867) );
  NAND2X0 U875 ( .IN1(n282), .IN2(n280), .QN(n868) );
  NAND2X0 U876 ( .IN1(n282), .IN2(n299), .QN(n869) );
  NAND3X0 U877 ( .IN1(n867), .IN2(n868), .IN3(n869), .QN(n277) );
  XOR3X1 U878 ( .IN1(n462), .IN2(n495), .IN3(n316), .Q(n310) );
  NAND2X0 U879 ( .IN1(n462), .IN2(n495), .QN(n870) );
  NAND2X1 U880 ( .IN1(n462), .IN2(n316), .QN(n871) );
  NAND2X0 U881 ( .IN1(n495), .IN2(n316), .QN(n872) );
  XOR2X1 U882 ( .IN1(n307), .IN2(n290), .Q(n873) );
  XOR2X2 U883 ( .IN1(n873), .IN2(n309), .Q(n284) );
  NAND2X0 U884 ( .IN1(n307), .IN2(n290), .QN(n874) );
  NAND2X0 U885 ( .IN1(n307), .IN2(n309), .QN(n875) );
  NAND2X0 U886 ( .IN1(n290), .IN2(n309), .QN(n876) );
  NAND3X0 U887 ( .IN1(n874), .IN2(n875), .IN3(n876), .QN(n283) );
  OR2X4 U888 ( .IN1(n554), .IN2(n677), .Q(n411) );
  NAND2X0 U889 ( .IN1(n294), .IN2(n311), .QN(n877) );
  NAND2X0 U890 ( .IN1(n647), .IN2(n311), .QN(n878) );
  NAND2X0 U891 ( .IN1(n647), .IN2(n294), .QN(n879) );
  NAND3X0 U892 ( .IN1(n877), .IN2(n879), .IN3(n878), .QN(n285) );
  XOR3X1 U893 ( .IN1(n506), .IN2(n539), .IN3(n451), .Q(n312) );
  NAND2X0 U894 ( .IN1(n451), .IN2(n506), .QN(n880) );
  NAND2X0 U895 ( .IN1(n539), .IN2(n506), .QN(n881) );
  NAND2X1 U896 ( .IN1(n539), .IN2(n451), .QN(n882) );
  NAND3X0 U897 ( .IN1(n880), .IN2(n882), .IN3(n881), .QN(n311) );
  OR2X4 U898 ( .IN1(n550), .IN2(n573), .Q(n539) );
  XOR2X1 U899 ( .IN1(n343), .IN2(n328), .Q(n883) );
  XOR2X2 U900 ( .IN1(n883), .IN2(n326), .Q(n322) );
  NAND2X0 U901 ( .IN1(n328), .IN2(n326), .QN(n884) );
  NAND2X0 U902 ( .IN1(n343), .IN2(n326), .QN(n885) );
  NAND2X0 U903 ( .IN1(n343), .IN2(n328), .QN(n886) );
  NAND3X0 U904 ( .IN1(n643), .IN2(n886), .IN3(n648), .QN(n321) );
  XOR2X2 U905 ( .IN1(n349), .IN2(n485), .Q(n887) );
  NAND2X0 U906 ( .IN1(n529), .IN2(n441), .QN(n888) );
  NAND2X0 U907 ( .IN1(n529), .IN2(n518), .QN(n889) );
  NAND2X0 U908 ( .IN1(n441), .IN2(n518), .QN(n890) );
  NAND2X0 U909 ( .IN1(n349), .IN2(n485), .QN(n891) );
  NAND2X0 U910 ( .IN1(n349), .IN2(n332), .QN(n892) );
  NAND2X0 U911 ( .IN1(n485), .IN2(n332), .QN(n893) );
  NAND3X0 U912 ( .IN1(n891), .IN2(n892), .IN3(n893), .QN(n325) );
  OR2X4 U913 ( .IN1(n767), .IN2(n677), .Q(n410) );
  XNOR2X1 U914 ( .IN1(n894), .IN2(n13), .Q(product[13]) );
  AO21X1 U915 ( .IN1(n644), .IN2(n107), .IN3(n108), .Q(n894) );
  XOR3X1 U916 ( .IN1(n671), .IN2(n323), .IN3(n304), .Q(n300) );
  NAND2X0 U917 ( .IN1(n304), .IN2(n321), .QN(n895) );
  NAND2X0 U918 ( .IN1(n323), .IN2(n321), .QN(n896) );
  NAND3X0 U919 ( .IN1(n895), .IN2(n897), .IN3(n896), .QN(n299) );
  XOR3X1 U920 ( .IN1(n238), .IN2(n253), .IN3(n251), .Q(n234) );
  NAND2X0 U921 ( .IN1(n238), .IN2(n253), .QN(n899) );
  NAND2X0 U922 ( .IN1(n238), .IN2(n251), .QN(n900) );
  NAND2X0 U923 ( .IN1(n253), .IN2(n251), .QN(n901) );
  NAND3X0 U924 ( .IN1(n899), .IN2(n900), .IN3(n901), .QN(n233) );
  NAND2X0 U925 ( .IN1(n249), .IN2(n236), .QN(n902) );
  NAND2X0 U926 ( .IN1(n249), .IN2(n234), .QN(n903) );
  NAND2X0 U927 ( .IN1(n236), .IN2(n234), .QN(n904) );
  NAND3X0 U928 ( .IN1(n904), .IN2(n903), .IN3(n902), .QN(n231) );
  NAND2X0 U929 ( .IN1(n480), .IN2(n257), .QN(n905) );
  NAND2X0 U930 ( .IN1(n425), .IN2(n257), .QN(n906) );
  NAND3X0 U931 ( .IN1(n905), .IN2(n907), .IN3(n906), .QN(n237) );
  XOR3X1 U932 ( .IN1(n361), .IN2(n363), .IN3(n348), .Q(n342) );
  NAND2X0 U933 ( .IN1(n361), .IN2(n363), .QN(n908) );
  NAND2X0 U934 ( .IN1(n361), .IN2(n348), .QN(n909) );
  NAND2X1 U935 ( .IN1(n363), .IN2(n348), .QN(n910) );
  NAND3X0 U936 ( .IN1(n908), .IN2(n909), .IN3(n910), .QN(n341) );
  XOR2X2 U937 ( .IN1(n911), .IN2(n341), .Q(n320) );
  NAND2X0 U938 ( .IN1(n324), .IN2(n709), .QN(n912) );
  NAND2X0 U939 ( .IN1(n324), .IN2(n341), .QN(n913) );
  NAND2X0 U940 ( .IN1(n341), .IN2(n709), .QN(n914) );
  NAND3X0 U941 ( .IN1(n912), .IN2(n913), .IN3(n914), .QN(n319) );
  XOR2X2 U942 ( .IN1(n279), .IN2(n264), .Q(n915) );
  XOR2X2 U943 ( .IN1(n915), .IN2(n262), .Q(n260) );
  NAND2X1 U944 ( .IN1(n266), .IN2(n283), .QN(n916) );
  NAND2X0 U945 ( .IN1(n266), .IN2(n281), .QN(n917) );
  NAND2X0 U946 ( .IN1(n283), .IN2(n281), .QN(n918) );
  NAND2X0 U947 ( .IN1(n693), .IN2(n264), .QN(n919) );
  NAND2X0 U948 ( .IN1(n693), .IN2(n262), .QN(n920) );
  NAND2X0 U949 ( .IN1(n264), .IN2(n262), .QN(n921) );
  NAND3X0 U950 ( .IN1(n919), .IN2(n920), .IN3(n921), .QN(n259) );
  OAI21X2 U951 ( .IN1(n100), .IN2(n128), .IN3(n101), .QN(n922) );
  XOR3X1 U952 ( .IN1(n325), .IN2(n308), .IN3(n625), .Q(n302) );
  NAND2X0 U953 ( .IN1(n325), .IN2(n308), .QN(n923) );
  NAND2X0 U954 ( .IN1(n325), .IN2(n306), .QN(n924) );
  NAND2X0 U955 ( .IN1(n308), .IN2(n306), .QN(n925) );
  NAND3X0 U956 ( .IN1(n924), .IN2(n925), .IN3(n923), .QN(n301) );
  NAND2X0 U957 ( .IN1(n284), .IN2(n303), .QN(n927) );
  NAND2X0 U958 ( .IN1(n284), .IN2(n301), .QN(n928) );
  NAND2X0 U959 ( .IN1(n303), .IN2(n301), .QN(n929) );
  NAND3X0 U960 ( .IN1(n929), .IN2(n928), .IN3(n927), .QN(n279) );
  NAND2X0 U961 ( .IN1(n246), .IN2(n683), .QN(n930) );
  NAND2X0 U962 ( .IN1(n248), .IN2(n683), .QN(n931) );
  NAND3X0 U963 ( .IN1(n930), .IN2(n932), .IN3(n931), .QN(n243) );
  XOR2X2 U964 ( .IN1(n959), .IN2(n960), .Q(product[22]) );
  XOR3X1 U965 ( .IN1(n474), .IN2(n452), .IN3(n496), .Q(n330) );
  NAND2X0 U966 ( .IN1(n474), .IN2(n452), .QN(n933) );
  NAND2X0 U967 ( .IN1(n474), .IN2(n496), .QN(n934) );
  NAND2X0 U968 ( .IN1(n452), .IN2(n496), .QN(n935) );
  XOR2X2 U969 ( .IN1(n936), .IN2(n329), .Q(n306) );
  NAND2X0 U970 ( .IN1(n314), .IN2(n331), .QN(n937) );
  NAND2X0 U971 ( .IN1(n314), .IN2(n329), .QN(n938) );
  NAND2X0 U972 ( .IN1(n331), .IN2(n329), .QN(n939) );
  NAND3X0 U973 ( .IN1(n937), .IN2(n938), .IN3(n939), .QN(n305) );
  NAND2X0 U974 ( .IN1(n285), .IN2(n287), .QN(n940) );
  NAND2X0 U975 ( .IN1(n285), .IN2(n268), .QN(n941) );
  NAND2X0 U976 ( .IN1(n287), .IN2(n268), .QN(n942) );
  NAND3X0 U977 ( .IN1(n941), .IN2(n940), .IN3(n942), .QN(n263) );
  NAND2X0 U978 ( .IN1(n619), .IN2(n642), .QN(n944) );
  NAND2X0 U979 ( .IN1(n619), .IN2(n263), .QN(n945) );
  NAND2X0 U980 ( .IN1(n642), .IN2(n263), .QN(n946) );
  NAND2X0 U981 ( .IN1(n184), .IN2(n132), .QN(n947) );
  NAND2X0 U982 ( .IN1(n183), .IN2(n678), .QN(n16) );
  NAND2X0 U983 ( .IN1(n185), .IN2(n135), .QN(n18) );
  XOR2X2 U984 ( .IN1(n955), .IN2(n956), .Q(product[19]) );
  INVX0 U985 ( .INP(n128), .ZN(n127) );
  INVX0 U986 ( .INP(n137), .ZN(n136) );
  NOR2X0 U987 ( .IN1(n116), .IN2(n673), .QN(n107) );
  INVX0 U988 ( .INP(n114), .ZN(n116) );
  XNOR2X1 U989 ( .IN1(n948), .IN2(n19), .Q(product[7]) );
  AO21X1 U990 ( .IN1(n149), .IN2(n951), .IN3(n952), .Q(n948) );
  NAND2X0 U991 ( .IN1(n178), .IN2(n93), .QN(n11) );
  INVX0 U992 ( .INP(n691), .ZN(n178) );
  NAND2X0 U993 ( .IN1(n816), .IN2(n121), .QN(n15) );
  INVX0 U994 ( .INP(n125), .ZN(n183) );
  INVX0 U995 ( .INP(n97), .ZN(n95) );
  NAND2X0 U996 ( .IN1(n181), .IN2(n112), .QN(n14) );
  INVX0 U997 ( .INP(n673), .ZN(n181) );
  INVX0 U998 ( .INP(n650), .ZN(n180) );
  NAND2X0 U999 ( .IN1(n180), .IN2(n105), .QN(n13) );
  INVX0 U1000 ( .INP(n131), .ZN(n184) );
  INVX0 U1001 ( .INP(n143), .ZN(n141) );
  INVX0 U1002 ( .INP(n134), .ZN(n185) );
  NAND2X0 U1003 ( .IN1(n95), .IN2(n674), .QN(n12) );
  NAND2X0 U1004 ( .IN1(n176), .IN2(n77), .QN(n9) );
  INVX0 U1005 ( .INP(n820), .ZN(n176) );
  NAND2X0 U1006 ( .IN1(n175), .IN2(n621), .QN(n8) );
  INVX0 U1007 ( .INP(n65), .ZN(n175) );
  INVX0 U1008 ( .INP(n58), .ZN(n56) );
  INVX0 U1009 ( .INP(n86), .ZN(n88) );
  NAND2X0 U1010 ( .IN1(n352), .IN2(n365), .QN(n135) );
  NAND2X0 U1011 ( .IN1(n259), .IN2(n244), .QN(n98) );
  NOR2X0 U1012 ( .IN1(n352), .IN2(n365), .QN(n134) );
  NOR2X0 U1013 ( .IN1(n336), .IN2(n351), .QN(n131) );
  NAND2X0 U1014 ( .IN1(n336), .IN2(n351), .QN(n132) );
  NAND2X0 U1015 ( .IN1(n278), .IN2(n297), .QN(n112) );
  NOR2X0 U1016 ( .IN1(n388), .IN2(n395), .QN(n153) );
  NAND2X0 U1017 ( .IN1(n177), .IN2(n640), .QN(n10) );
  INVX0 U1018 ( .INP(n81), .ZN(n177) );
  NAND2X0 U1019 ( .IN1(n298), .IN2(n317), .QN(n121) );
  NAND2X0 U1020 ( .IN1(n260), .IN2(n277), .QN(n105) );
  NAND2X0 U1021 ( .IN1(n366), .IN2(n377), .QN(n143) );
  OR2X1 U1022 ( .IN1(n366), .IN2(n377), .Q(n949) );
  OA21X1 U1023 ( .IN1(n950), .IN2(n153), .IN3(n154), .Q(n150) );
  OA21X1 U1024 ( .IN1(n156), .IN2(n158), .IN3(n157), .Q(n950) );
  OA21X1 U1025 ( .IN1(n167), .IN2(n170), .IN3(n168), .Q(n164) );
  OR2X1 U1026 ( .IN1(n378), .IN2(n387), .Q(n951) );
  AND2X1 U1027 ( .IN1(n378), .IN2(n387), .Q(n952) );
  INVX0 U1028 ( .INP(n622), .ZN(n57) );
  OA21X1 U1029 ( .IN1(n161), .IN2(n164), .IN3(n162), .Q(n158) );
  INVX0 U1030 ( .INP(n87), .ZN(n89) );
  NAND2X0 U1031 ( .IN1(n388), .IN2(n395), .QN(n154) );
  NOR2X0 U1032 ( .IN1(n229), .IN2(n218), .QN(n81) );
  NOR2X0 U1033 ( .IN1(n406), .IN2(n537), .QN(n167) );
  NAND2X0 U1034 ( .IN1(n406), .IN2(n537), .QN(n168) );
  NAND2X0 U1035 ( .IN1(n58), .IN2(n25), .QN(n23) );
  AND2X1 U1036 ( .IN1(n961), .IN2(n52), .Q(n954) );
  NAND2X0 U1037 ( .IN1(n207), .IN2(n200), .QN(n68) );
  NOR2X0 U1038 ( .IN1(n402), .IN2(n405), .QN(n161) );
  NAND2X0 U1039 ( .IN1(n402), .IN2(n405), .QN(n162) );
  NOR2X0 U1040 ( .IN1(n396), .IN2(n401), .QN(n156) );
  AO21X1 U1041 ( .IN1(n1), .IN2(n63), .IN3(n64), .Q(n955) );
  AND2X1 U1042 ( .IN1(n680), .IN2(n61), .Q(n956) );
  INVX0 U1043 ( .INP(n37), .ZN(n35) );
  NAND2X0 U1044 ( .IN1(n549), .IN2(n538), .QN(n170) );
  NOR2X0 U1045 ( .IN1(n708), .IN2(n561), .QN(n538) );
  NAND2X0 U1046 ( .IN1(n396), .IN2(n401), .QN(n157) );
  INVX0 U1047 ( .INP(a[1]), .ZN(n572) );
  INVX0 U1048 ( .INP(b[4]), .ZN(n557) );
  INVX0 U1049 ( .INP(a[4]), .ZN(n569) );
  INVX0 U1050 ( .INP(b[1]), .ZN(n560) );
  NOR2X0 U1051 ( .IN1(n672), .IN2(n561), .QN(n514) );
  NOR2X0 U1052 ( .IN1(n699), .IN2(n561), .QN(n526) );
  NAND2X0 U1053 ( .IN1(n194), .IN2(n199), .QN(n61) );
  NOR2X0 U1054 ( .IN1(n199), .IN2(n194), .QN(n60) );
  NAND2X0 U1055 ( .IN1(n193), .IN2(n190), .QN(n52) );
  AO21X1 U1056 ( .IN1(n922), .IN2(n43), .IN3(n44), .Q(n957) );
  AND2X1 U1057 ( .IN1(n962), .IN2(n41), .Q(n958) );
  AO21X1 U1058 ( .IN1(n922), .IN2(n30), .IN3(n31), .Q(n959) );
  AND2X1 U1059 ( .IN1(n171), .IN2(n28), .Q(n960) );
  OR2X1 U1060 ( .IN1(n193), .IN2(n190), .Q(n961) );
  INVX0 U1061 ( .INP(n41), .ZN(n39) );
  INVX0 U1062 ( .INP(a[0]), .ZN(n573) );
  INVX0 U1063 ( .INP(a[3]), .ZN(n570) );
  INVX0 U1064 ( .INP(b[5]), .ZN(n556) );
  INVX0 U1065 ( .INP(a[5]), .ZN(n568) );
  INVX0 U1066 ( .INP(b[3]), .ZN(n558) );
  INVX0 U1067 ( .INP(b[2]), .ZN(n559) );
  OR2X1 U1068 ( .IN1(n189), .IN2(n188), .Q(n962) );
  NAND2X0 U1069 ( .IN1(n189), .IN2(n188), .QN(n41) );
  NAND2X0 U1070 ( .IN1(n187), .IN2(n407), .QN(n28) );
  NOR2X0 U1071 ( .IN1(n187), .IN2(n407), .QN(n27) );
  OR2X1 U1072 ( .IN1(n784), .IN2(n550), .Q(n443) );
  OR2X1 U1073 ( .IN1(n712), .IN2(n550), .Q(n467) );
  NOR2X0 U1074 ( .IN1(n550), .IN2(n677), .QN(n407) );
  OR2X1 U1075 ( .IN1(n695), .IN2(n550), .Q(n431) );
  INVX0 U1076 ( .INP(b[11]), .ZN(n550) );
  INVX0 U1077 ( .INP(a[11]), .ZN(n562) );
  INVX0 U1078 ( .INP(b[10]), .ZN(n551) );
  INVX0 U1079 ( .INP(a[2]), .ZN(n571) );
  INVX0 U1080 ( .INP(b[9]), .ZN(n552) );
  NOR2X0 U1081 ( .IN1(n679), .IN2(n561), .QN(n466) );
  NOR2X0 U1082 ( .IN1(n638), .IN2(n65), .QN(n63) );
  INVX0 U1083 ( .INP(n638), .ZN(n70) );
  NAND2X0 U1084 ( .IN1(n86), .IN2(n641), .QN(n3) );
  NOR2X0 U1085 ( .IN1(n36), .IN2(n27), .QN(n25) );
  INVX0 U1086 ( .INP(n36), .ZN(n34) );
  INVX0 U1087 ( .INP(a[9]), .ZN(n564) );
  NOR2X0 U1088 ( .IN1(n629), .IN2(n573), .QN(n549) );
  NOR2X0 U1089 ( .IN1(n629), .IN2(n708), .QN(n537) );
  NOR2X0 U1090 ( .IN1(n672), .IN2(n629), .QN(n513) );
  NOR2X0 U1091 ( .IN1(n629), .IN2(n699), .QN(n525) );
  NOR2X0 U1092 ( .IN1(n566), .IN2(n560), .QN(n465) );
  NOR2X0 U1093 ( .IN1(n682), .IN2(n573), .QN(n547) );
  NOR2X0 U1094 ( .IN1(n682), .IN2(n706), .QN(n535) );
  NOR2X0 U1095 ( .IN1(n682), .IN2(n571), .QN(n523) );
  NOR2X0 U1096 ( .IN1(n558), .IN2(n570), .QN(n511) );
  NOR2X0 U1097 ( .IN1(n566), .IN2(n558), .QN(n463) );
  NOR2X0 U1098 ( .IN1(n711), .IN2(n561), .QN(n502) );
  NOR2X0 U1099 ( .IN1(n569), .IN2(n560), .QN(n501) );
  NOR2X0 U1100 ( .IN1(n772), .IN2(n561), .QN(n490) );
  NOR2X0 U1101 ( .IN1(n772), .IN2(n560), .QN(n489) );
  NOR2X0 U1102 ( .IN1(n568), .IN2(n682), .QN(n487) );
  INVX0 U1103 ( .INP(b[7]), .ZN(n554) );
  INVX0 U1104 ( .INP(b[6]), .ZN(n555) );
  INVX0 U1105 ( .INP(a[6]), .ZN(n567) );
  INVX0 U1106 ( .INP(a[8]), .ZN(n565) );
  INVX0 U1107 ( .INP(b[8]), .ZN(n553) );
  INVX0 U1108 ( .INP(a[7]), .ZN(n566) );
  NOR2X0 U1109 ( .IN1(n563), .IN2(n558), .QN(n427) );
  NOR2X0 U1110 ( .IN1(n697), .IN2(n637), .QN(n429) );
  INVX0 U1111 ( .INP(a[10]), .ZN(n563) );
  NOR2X0 U1112 ( .IN1(n701), .IN2(n705), .QN(n420) );
  NOR2X0 U1113 ( .IN1(n568), .IN2(n687), .QN(n480) );
  NOR2X0 U1114 ( .IN1(n566), .IN2(n701), .QN(n456) );
  NOR2X0 U1115 ( .IN1(n551), .IN2(n573), .QN(n540) );
  NOR2X0 U1116 ( .IN1(n551), .IN2(n571), .QN(n516) );
  NOR2X0 U1117 ( .IN1(n551), .IN2(n570), .QN(n504) );
  NOR2X0 U1118 ( .IN1(n564), .IN2(n561), .QN(n442) );
  NOR2X0 U1119 ( .IN1(n564), .IN2(n560), .QN(n441) );
  NOR2X0 U1120 ( .IN1(n630), .IN2(n687), .QN(n432) );
  NOR2X0 U1121 ( .IN1(n318), .IN2(n335), .QN(n125) );
  NOR2X0 U1122 ( .IN1(n686), .IN2(n573), .QN(n545) );
  NOR2X0 U1123 ( .IN1(n659), .IN2(n686), .QN(n533) );
  NOR2X0 U1124 ( .IN1(n556), .IN2(n697), .QN(n425) );
  NOR2X0 U1125 ( .IN1(n686), .IN2(n695), .QN(n437) );
  NOR2X0 U1126 ( .IN1(n686), .IN2(n711), .QN(n497) );
  NOR2X0 U1127 ( .IN1(n686), .IN2(n566), .QN(n461) );
  NOR2X0 U1128 ( .IN1(n556), .IN2(n772), .QN(n485) );
  NOR2X0 U1129 ( .IN1(n556), .IN2(n688), .QN(n521) );
  NOR2X0 U1130 ( .IN1(n556), .IN2(n672), .QN(n509) );
  NOR2X0 U1131 ( .IN1(n684), .IN2(n573), .QN(n548) );
  NOR2X0 U1132 ( .IN1(n706), .IN2(n684), .QN(n536) );
  NOR2X0 U1133 ( .IN1(n559), .IN2(n571), .QN(n524) );
  NOR2X0 U1134 ( .IN1(n772), .IN2(n684), .QN(n488) );
  NOR2X0 U1135 ( .IN1(n672), .IN2(n559), .QN(n512) );
  NOR2X0 U1136 ( .IN1(n711), .IN2(n559), .QN(n500) );
  NOR2X0 U1137 ( .IN1(n714), .IN2(n684), .QN(n464) );
  NOR2X0 U1138 ( .IN1(n563), .IN2(n559), .QN(n428) );
  NOR2X0 U1139 ( .IN1(n564), .IN2(n559), .QN(n440) );
  NAND2X0 U1140 ( .IN1(n102), .IN2(n114), .QN(n100) );
  NOR2X0 U1141 ( .IN1(n554), .IN2(n630), .QN(n435) );
  NOR2X0 U1142 ( .IN1(n554), .IN2(n566), .QN(n459) );
  NOR2X0 U1143 ( .IN1(n721), .IN2(n705), .QN(n423) );
  NOR2X0 U1144 ( .IN1(n568), .IN2(n554), .QN(n483) );
  NOR2X0 U1145 ( .IN1(n554), .IN2(n569), .QN(n495) );
  NOR2X0 U1146 ( .IN1(n721), .IN2(n570), .QN(n507) );
  NOR2X0 U1147 ( .IN1(n554), .IN2(n659), .QN(n531) );
  NOR2X0 U1148 ( .IN1(n721), .IN2(n573), .QN(n543) );
  NOR2X0 U1149 ( .IN1(n721), .IN2(n688), .QN(n519) );
  NOR2X0 U1150 ( .IN1(n3), .IN2(n56), .QN(n54) );
  NAND2X0 U1151 ( .IN1(n217), .IN2(n208), .QN(n77) );
  NOR2X0 U1152 ( .IN1(n217), .IN2(n208), .QN(n76) );
  NOR2X0 U1153 ( .IN1(n557), .IN2(n573), .QN(n546) );
  NOR2X0 U1154 ( .IN1(n703), .IN2(n659), .QN(n534) );
  NOR2X0 U1155 ( .IN1(n772), .IN2(n703), .QN(n486) );
  NOR2X0 U1156 ( .IN1(n557), .IN2(n571), .QN(n522) );
  NOR2X0 U1157 ( .IN1(n679), .IN2(n557), .QN(n462) );
  NOR2X0 U1158 ( .IN1(n703), .IN2(n569), .QN(n498) );
  NOR2X0 U1159 ( .IN1(n570), .IN2(n703), .QN(n510) );
  NOR2X0 U1160 ( .IN1(n563), .IN2(n557), .QN(n426) );
  NOR2X0 U1161 ( .IN1(n675), .IN2(n705), .QN(n421) );
  NOR2X0 U1162 ( .IN1(n568), .IN2(n675), .QN(n481) );
  NOR2X0 U1163 ( .IN1(n552), .IN2(n573), .QN(n541) );
  NOR2X0 U1164 ( .IN1(n675), .IN2(n564), .QN(n433) );
  NOR2X0 U1165 ( .IN1(n566), .IN2(n675), .QN(n457) );
  NOR2X0 U1166 ( .IN1(n552), .IN2(n572), .QN(n529) );
  NOR2X0 U1167 ( .IN1(n552), .IN2(n571), .QN(n517) );
  NOR2X0 U1168 ( .IN1(n552), .IN2(n570), .QN(n505) );
  NOR2X0 U1169 ( .IN1(n552), .IN2(n569), .QN(n493) );
  NOR2X0 U1170 ( .IN1(n88), .IN2(n776), .QN(n79) );
  NOR2X0 U1171 ( .IN1(n568), .IN2(n766), .QN(n482) );
  NOR2X0 U1172 ( .IN1(n766), .IN2(n563), .QN(n422) );
  NOR2X0 U1173 ( .IN1(n566), .IN2(n767), .QN(n458) );
  NOR2X0 U1174 ( .IN1(n766), .IN2(n569), .QN(n494) );
  NOR2X0 U1175 ( .IN1(n767), .IN2(n659), .QN(n530) );
  NOR2X0 U1176 ( .IN1(n766), .IN2(n695), .QN(n434) );
  NOR2X0 U1177 ( .IN1(n767), .IN2(n573), .QN(n542) );
  NOR2X0 U1178 ( .IN1(n553), .IN2(n571), .QN(n518) );
  NOR2X0 U1179 ( .IN1(n766), .IN2(n570), .QN(n506) );
  NAND2X0 U1180 ( .IN1(n949), .IN2(n649), .QN(n19) );
  NAND2X0 U1181 ( .IN1(n949), .IN2(n951), .QN(n138) );
  NOR2X0 U1182 ( .IN1(n772), .IN2(n710), .QN(n484) );
  NOR2X0 U1183 ( .IN1(n555), .IN2(n672), .QN(n508) );
  NOR2X0 U1184 ( .IN1(n710), .IN2(n571), .QN(n520) );
  NOR2X0 U1185 ( .IN1(n710), .IN2(n569), .QN(n496) );
  NOR2X0 U1186 ( .IN1(n710), .IN2(n630), .QN(n436) );
  NOR2X0 U1187 ( .IN1(n555), .IN2(n563), .QN(n424) );
  NOR2X0 U1188 ( .IN1(n555), .IN2(n573), .QN(n544) );
  NOR2X0 U1189 ( .IN1(n710), .IN2(n659), .QN(n532) );
  NOR2X0 U1190 ( .IN1(n564), .IN2(n558), .QN(n439) );
  NAND2X0 U1191 ( .IN1(n229), .IN2(n218), .QN(n84) );
  NOR2X0 U1192 ( .IN1(n244), .IN2(n259), .QN(n97) );
  NAND2X0 U1193 ( .IN1(n230), .IN2(n243), .QN(n93) );
  NOR2X0 U1194 ( .IN1(n243), .IN2(n230), .QN(n92) );
  NOR2X0 U1195 ( .IN1(n784), .IN2(n561), .QN(n454) );
  NOR2X0 U1196 ( .IN1(n753), .IN2(n646), .QN(n444) );
  NOR2X0 U1197 ( .IN1(n686), .IN2(n753), .QN(n449) );
  NOR2X0 U1198 ( .IN1(n554), .IN2(n784), .QN(n447) );
  NOR2X0 U1199 ( .IN1(n753), .IN2(n560), .QN(n453) );
  NOR2X0 U1200 ( .IN1(n784), .IN2(n675), .QN(n445) );
  NOR2X0 U1201 ( .IN1(n766), .IN2(n784), .QN(n446) );
  NOR2X0 U1202 ( .IN1(n710), .IN2(n753), .QN(n448) );
  NOR2X0 U1203 ( .IN1(n753), .IN2(n558), .QN(n451) );
  NOR2X0 U1204 ( .IN1(n565), .IN2(n557), .QN(n450) );
  NOR2X0 U1205 ( .IN1(n565), .IN2(n559), .QN(n452) );
  NOR2X0 U1206 ( .IN1(n3), .IN2(n45), .QN(n43) );
  NOR2X0 U1207 ( .IN1(n702), .IN2(n125), .QN(n114) );
  NOR2X0 U1208 ( .IN1(n317), .IN2(n298), .QN(n120) );
  NOR2X0 U1209 ( .IN1(n3), .IN2(n23), .QN(n21) );
  NAND2X0 U1210 ( .IN1(n58), .IN2(n961), .QN(n45) );
  NAND2X0 U1211 ( .IN1(n961), .IN2(n962), .QN(n36) );
  NOR2X0 U1212 ( .IN1(n638), .IN2(n32), .QN(n30) );
  NAND2X0 U1213 ( .IN1(n58), .IN2(n34), .QN(n32) );
  NOR2X0 U1214 ( .IN1(n65), .IN2(n60), .QN(n58) );
  NOR2X0 U1215 ( .IN1(n207), .IN2(n200), .QN(n65) );
  NOR2X0 U1216 ( .IN1(n628), .IN2(n569), .QN(n492) );
  NOR2X0 U1217 ( .IN1(n650), .IN2(n673), .QN(n102) );
  NOR2X0 U1218 ( .IN1(n260), .IN2(n277), .QN(n104) );
  NOR2X0 U1219 ( .IN1(n131), .IN2(n134), .QN(n129) );
  NOR2X0 U1220 ( .IN1(n553), .IN2(n567), .QN(n470) );
  NOR2X0 U1221 ( .IN1(n712), .IN2(n675), .QN(n469) );
  NOR2X0 U1222 ( .IN1(n555), .IN2(n567), .QN(n472) );
  NOR2X0 U1223 ( .IN1(n556), .IN2(n712), .QN(n473) );
  NOR2X0 U1224 ( .IN1(n721), .IN2(n712), .QN(n471) );
  NOR2X0 U1225 ( .IN1(n561), .IN2(n712), .QN(n478) );
  NOR2X0 U1226 ( .IN1(n712), .IN2(n682), .QN(n475) );
  NOR2X0 U1227 ( .IN1(n712), .IN2(n560), .QN(n477) );
  NOR2X0 U1228 ( .IN1(n567), .IN2(n557), .QN(n474) );
  NOR2X0 U1229 ( .IN1(n567), .IN2(n559), .QN(n476) );
  NOR2X0 U1230 ( .IN1(n558), .IN2(n711), .QN(n499) );
  NOR2X0 U1231 ( .IN1(n691), .IN2(n97), .QN(n86) );
  NOR2X0 U1232 ( .IN1(n820), .IN2(n81), .QN(n74) );
  OAI21X2 U1233 ( .IN1(n100), .IN2(n128), .IN3(n101), .QN(n1) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2 ( in_a, in_b, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [11:0] \output ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  wire   [23:7] pre_out;
  wire   [11:0] rnd_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2_DW01_inc_2 add_37_round ( .A({
        n2, pre_out[18:7]}), .SUM({rnd_out, SYNOPSYS_UNCONNECTED__0}) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2_DW_mult_tc_6 mult_35 ( .a(in_a), 
        .b(in_b), .product({pre_out, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7}) );
  INVX0 U2 ( .INP(pre_out[19]), .ZN(n1) );
  INVX0 U3 ( .INP(n1), .ZN(n2) );
  OR3X1 U4 ( .IN1(n11), .IN2(n3), .IN3(n12), .Q(n8) );
  AND2X1 U5 ( .IN1(n19), .IN2(n18), .Q(n9) );
  AND2X1 U6 ( .IN1(n7), .IN2(n18), .Q(n10) );
  INVX0 U7 ( .INP(pre_out[19]), .ZN(n3) );
  NAND2X0 U8 ( .IN1(n19), .IN2(n20), .QN(n4) );
  NAND2X0 U9 ( .IN1(n19), .IN2(n20), .QN(n5) );
  AND2X2 U10 ( .IN1(n7), .IN2(n18), .Q(n6) );
  NAND3X0 U11 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(n7) );
  AO21X1 U12 ( .IN1(rnd_out[10]), .IN2(n4), .IN3(n9), .Q(\output [10]) );
  AO21X1 U13 ( .IN1(rnd_out[7]), .IN2(n21), .IN3(n9), .Q(\output [7]) );
  AO21X1 U14 ( .IN1(rnd_out[6]), .IN2(n21), .IN3(n9), .Q(\output [6]) );
  INVX0 U15 ( .INP(n4), .ZN(n22) );
  AO221X1 U16 ( .IN1(rnd_out[0]), .IN2(n18), .IN3(n17), .IN4(rnd_out[0]), 
        .IN5(n10), .Q(\output [0]) );
  INVX0 U17 ( .INP(pre_out[23]), .ZN(n18) );
  NAND2X0 U18 ( .IN1(pre_out[23]), .IN2(pre_out[20]), .QN(n12) );
  NOR2X0 U19 ( .IN1(n11), .IN2(n12), .QN(n13) );
  AO21X1 U20 ( .IN1(rnd_out[8]), .IN2(n21), .IN3(n6), .Q(\output [8]) );
  NOR2X0 U21 ( .IN1(pre_out[20]), .IN2(pre_out[23]), .QN(n14) );
  AO21X1 U22 ( .IN1(rnd_out[1]), .IN2(n4), .IN3(n6), .Q(\output [1]) );
  AO21X1 U23 ( .IN1(rnd_out[9]), .IN2(n4), .IN3(n6), .Q(\output [9]) );
  INVX0 U24 ( .INP(n8), .ZN(n17) );
  NAND2X0 U25 ( .IN1(n2), .IN2(n13), .QN(n20) );
  AO21X1 U26 ( .IN1(rnd_out[5]), .IN2(n21), .IN3(n6), .Q(\output [5]) );
  INVX0 U27 ( .INP(pre_out[19]), .ZN(n15) );
  NOR2X0 U28 ( .IN1(pre_out[21]), .IN2(pre_out[22]), .QN(n16) );
  NAND2X0 U29 ( .IN1(pre_out[22]), .IN2(pre_out[21]), .QN(n11) );
  NAND2X0 U30 ( .IN1(n19), .IN2(n8), .QN(n21) );
  NAND3X0 U31 ( .IN1(n15), .IN2(n16), .IN3(n14), .QN(n19) );
  AO21X1 U32 ( .IN1(rnd_out[2]), .IN2(n5), .IN3(n10), .Q(\output [2]) );
  AO21X1 U33 ( .IN1(rnd_out[3]), .IN2(n5), .IN3(n9), .Q(\output [3]) );
  AO21X1 U34 ( .IN1(rnd_out[4]), .IN2(n5), .IN3(n6), .Q(\output [4]) );
  MUX21X1 U35 ( .IN1(rnd_out[11]), .IN2(pre_out[23]), .S(n22), .Q(\output [11]) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1_DW01_inc_2 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;
  wire   n2, n5, n6, n7, n8, n10, n11, n12, n14, n15, n18, n19, n20, n21, n22,
         n24, n26, n27, n28, n29, n33, n35, n36, n37, n38, n69, n70, n71, n72,
         n73, n74;
  assign n5 = A[11];
  assign n8 = A[10];
  assign n12 = A[9];
  assign n15 = A[8];
  assign n26 = A[5];
  assign n29 = A[4];
  assign n33 = A[3];
  assign n38 = A[1];

  XNOR2X1 U22 ( .IN1(n21), .IN2(n20), .Q(SUM[7]) );
  XOR2X1 U27 ( .IN1(n70), .IN2(n22), .Q(SUM[6]) );
  XOR2X1 U30 ( .IN1(n27), .IN2(n28), .Q(SUM[5]) );
  AND2X1 U54 ( .IN1(n24), .IN2(n19), .Q(n69) );
  NAND4X0 U55 ( .IN1(n26), .IN2(n29), .IN3(A[2]), .IN4(n73), .QN(n70) );
  AND2X4 U56 ( .IN1(n33), .IN2(n35), .Q(n71) );
  AND2X1 U57 ( .IN1(n38), .IN2(A[0]), .Q(n72) );
  AND4X1 U58 ( .IN1(n26), .IN2(n29), .IN3(A[2]), .IN4(n73), .Q(n24) );
  AND2X1 U59 ( .IN1(n33), .IN2(n72), .Q(n73) );
  AND2X1 U60 ( .IN1(A[2]), .IN2(n72), .Q(n35) );
  AND2X1 U61 ( .IN1(A[6]), .IN2(A[7]), .Q(n19) );
  XOR2X2 U62 ( .IN1(n10), .IN2(n8), .Q(SUM[10]) );
  NAND2X0 U63 ( .IN1(n24), .IN2(n19), .QN(n18) );
  NAND2X0 U64 ( .IN1(n12), .IN2(n15), .QN(n11) );
  XOR2X2 U65 ( .IN1(n7), .IN2(n6), .Q(SUM[11]) );
  AND2X1 U66 ( .IN1(n8), .IN2(n5), .Q(n74) );
  XOR2X1 U67 ( .IN1(n15), .IN2(n69), .Q(SUM[8]) );
  INVX0 U68 ( .INP(n26), .ZN(n27) );
  XOR2X1 U69 ( .IN1(n33), .IN2(n35), .Q(SUM[3]) );
  XOR2X1 U70 ( .IN1(n29), .IN2(n71), .Q(SUM[4]) );
  NOR2X0 U71 ( .IN1(n11), .IN2(n18), .QN(n10) );
  XNOR2X1 U72 ( .IN1(n12), .IN2(n14), .Q(SUM[9]) );
  NAND2X0 U73 ( .IN1(n10), .IN2(n8), .QN(n7) );
  NAND2X0 U74 ( .IN1(n15), .IN2(n69), .QN(n14) );
  INVX0 U75 ( .INP(n5), .ZN(n6) );
  XOR2X1 U76 ( .IN1(n38), .IN2(A[0]), .Q(SUM[1]) );
  XOR2X1 U77 ( .IN1(n36), .IN2(n37), .Q(SUM[2]) );
  XNOR2X1 U78 ( .IN1(n2), .IN2(A[12]), .Q(SUM[12]) );
  NAND2X0 U79 ( .IN1(n38), .IN2(A[0]), .QN(n37) );
  INVX0 U80 ( .INP(A[7]), .ZN(n20) );
  NAND2X0 U81 ( .IN1(n10), .IN2(n74), .QN(n2) );
  INVX0 U82 ( .INP(A[2]), .ZN(n36) );
  NAND2X0 U83 ( .IN1(n71), .IN2(n29), .QN(n28) );
  NOR2X0 U84 ( .IN1(n70), .IN2(n22), .QN(n21) );
  INVX0 U85 ( .INP(A[6]), .ZN(n22) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1_DW_mult_tc_7 ( a, b, 
        product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n4, n5, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50,
         n52, n54, n55, n56, n57, n63, n65, n66, n67, n68, n69, n70, n73, n74,
         n75, n78, n79, n81, n82, n83, n84, n85, n88, n90, n91, n92, n93, n96,
         n97, n99, n101, n102, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n116, n117, n118, n119, n120, n121, n124, n125, n126,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n145, n147, n148, n153, n154, n157, n158,
         n159, n160, n162, n163, n164, n167, n168, n170, n171, n176, n177,
         n178, n180, n181, n182, n183, n184, n185, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n299, n301, n303,
         n305, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n517, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673;
  assign n1 = a[0];
  assign n464 = a[11];
  assign n465 = a[10];
  assign n466 = a[9];
  assign n467 = a[8];
  assign n468 = a[7];
  assign n469 = a[6];
  assign n470 = a[5];
  assign n471 = a[4];
  assign n472 = a[3];
  assign n473 = a[2];
  assign n474 = a[1];
  assign n500 = b[11];
  assign n501 = b[9];
  assign n502 = b[7];
  assign n503 = b[5];
  assign n504 = b[3];
  assign n505 = b[1];

  AOI21X1 U8 ( .IN1(n646), .IN2(n23), .IN3(n24), .QN(product[23]) );
  OAI21X1 U10 ( .IN1(n25), .IN2(n594), .IN3(n26), .QN(n24) );
  AOI21X1 U12 ( .IN1(n46), .IN2(n27), .IN3(n28), .QN(n26) );
  OAI21X1 U14 ( .IN1(n29), .IN2(n39), .IN3(n30), .QN(n28) );
  OAI21X1 U22 ( .IN1(n34), .IN2(n4), .IN3(n35), .QN(n33) );
  AOI21X1 U24 ( .IN1(n46), .IN2(n36), .IN3(n37), .QN(n35) );
  AOI21X1 U32 ( .IN1(n645), .IN2(n41), .IN3(n42), .QN(n40) );
  OAI21X1 U34 ( .IN1(n43), .IN2(n599), .IN3(n44), .QN(n42) );
  OAI21X1 U38 ( .IN1(n47), .IN2(n68), .IN3(n48), .QN(n46) );
  AOI21X1 U40 ( .IN1(n608), .IN2(n666), .IN3(n50), .QN(n48) );
  OAI21X1 U50 ( .IN1(n56), .IN2(n599), .IN3(n57), .QN(n55) );
  AOI21X1 U52 ( .IN1(n70), .IN2(n665), .IN3(n608), .QN(n57) );
  XOR2X1 U61 ( .IN1(n73), .IN2(n10), .Q(product[18]) );
  OAI21X1 U64 ( .IN1(n67), .IN2(n4), .IN3(n68), .QN(n66) );
  XOR2X1 U73 ( .IN1(n82), .IN2(n11), .Q(product[17]) );
  AOI21X1 U74 ( .IN1(n646), .IN2(n74), .IN3(n75), .QN(n73) );
  AOI21X1 U78 ( .IN1(n91), .IN2(n78), .IN3(n79), .QN(n4) );
  OAI21X1 U80 ( .IN1(n605), .IN2(n88), .IN3(n81), .QN(n79) );
  AOI21X1 U86 ( .IN1(n646), .IN2(n83), .IN3(n84), .QN(n82) );
  OAI21X1 U102 ( .IN1(n102), .IN2(n96), .IN3(n97), .QN(n91) );
  XNOR2X1 U107 ( .IN1(n646), .IN2(n14), .Q(product[14]) );
  XOR2X1 U115 ( .IN1(n110), .IN2(n15), .Q(product[13]) );
  AOI21X1 U118 ( .IN1(n119), .IN2(n106), .IN3(n107), .QN(n105) );
  OAI21X1 U120 ( .IN1(n108), .IN2(n116), .IN3(n109), .QN(n107) );
  AOI21X1 U126 ( .IN1(n601), .IN2(n111), .IN3(n112), .QN(n110) );
  OAI21X1 U128 ( .IN1(n629), .IN2(n121), .IN3(n607), .QN(n112) );
  OAI21X1 U142 ( .IN1(n124), .IN2(n130), .IN3(n125), .QN(n119) );
  XNOR2X1 U147 ( .IN1(n601), .IN2(n18), .Q(product[10]) );
  AOI21X1 U148 ( .IN1(n131), .IN2(n183), .IN3(n600), .QN(n126) );
  XNOR2X1 U155 ( .IN1(n137), .IN2(n19), .Q(product[9]) );
  AOI21X1 U157 ( .IN1(n141), .IN2(n133), .IN3(n134), .QN(n132) );
  OAI21X1 U159 ( .IN1(n139), .IN2(n135), .IN3(n136), .QN(n134) );
  OAI21X1 U165 ( .IN1(n138), .IN2(n140), .IN3(n139), .QN(n137) );
  OAI21X1 U172 ( .IN1(n142), .IN2(n154), .IN3(n143), .QN(n141) );
  AOI21X1 U174 ( .IN1(n667), .IN2(n669), .IN3(n145), .QN(n143) );
  AOI21X1 U181 ( .IN1(n153), .IN2(n668), .IN3(n669), .QN(n148) );
  FADDX1 U205 ( .A(n315), .B(n325), .CI(n193), .CO(n189), .S(n190) );
  FADDX1 U206 ( .A(n194), .B(n316), .CI(n197), .CO(n191), .S(n192) );
  FADDX1 U208 ( .A(n198), .B(n317), .CI(n201), .CO(n195), .S(n196) );
  FADDX1 U209 ( .A(n326), .B(n337), .CI(n203), .CO(n197), .S(n198) );
  FADDX1 U210 ( .A(n202), .B(n209), .CI(n207), .CO(n199), .S(n200) );
  FADDX1 U211 ( .A(n204), .B(n327), .CI(n318), .CO(n201), .S(n202) );
  FADDX1 U214 ( .A(n319), .B(n328), .CI(n210), .CO(n207), .S(n208) );
  FADDX1 U215 ( .A(n338), .B(n349), .CI(n217), .CO(n209), .S(n210) );
  FADDX1 U218 ( .A(n339), .B(n218), .CI(n329), .CO(n215), .S(n216) );
  FADDX1 U221 ( .A(n226), .B(n233), .CI(n231), .CO(n221), .S(n222) );
  FADDX1 U222 ( .A(n340), .B(n350), .CI(n330), .CO(n223), .S(n224) );
  FADDX1 U223 ( .A(n235), .B(n361), .CI(n321), .CO(n225), .S(n226) );
  FADDX1 U227 ( .A(n236), .B(n362), .CI(n351), .CO(n233), .S(n234) );
  FADDX1 U231 ( .A(n342), .B(n255), .CI(n246), .CO(n241), .S(n242) );
  FADDX1 U232 ( .A(n602), .B(n363), .CI(n591), .CO(n243) );
  XNOR2X1 U233 ( .IN1(n322), .IN2(n374), .Q(n246) );
  OR2X1 U234 ( .IN1(n322), .IN2(n374), .Q(n245) );
  FADDX1 U238 ( .A(n375), .B(n333), .CI(n364), .CO(n253), .S(n254) );
  HADDX1 U239 ( .A0(n308), .B0(n323), .C1(n255), .SO(n256) );
  FADDX1 U240 ( .A(n267), .B(n262), .CI(n260), .CO(n257), .S(n258) );
  FADDX1 U242 ( .A(n271), .B(n376), .CI(n365), .CO(n261), .S(n262) );
  FADDX1 U243 ( .A(n334), .B(n324), .CI(n344), .CO(n263), .S(n264) );
  FADDX1 U244 ( .A(n275), .B(n270), .CI(n268), .CO(n265), .S(n266) );
  FADDX1 U246 ( .A(n377), .B(n345), .CI(n272), .CO(n269), .S(n270) );
  HADDX1 U247 ( .A0(n309), .B0(n335), .C1(n271), .SO(n272) );
  FADDX1 U248 ( .A(n281), .B(n278), .CI(n276), .CO(n273), .S(n274) );
  FADDX1 U249 ( .A(n283), .B(n378), .CI(n367), .CO(n275), .S(n276) );
  FADDX1 U252 ( .A(n284), .B(n357), .CI(n379), .CO(n281), .S(n282) );
  HADDX1 U253 ( .A0(n310), .B0(n347), .C1(n283), .SO(n284) );
  FADDX1 U254 ( .A(n380), .B(n291), .CI(n288), .CO(n285), .S(n286) );
  FADDX1 U255 ( .A(n358), .B(n348), .CI(n369), .CO(n287), .S(n288) );
  FADDX1 U256 ( .A(n292), .B(n370), .CI(n381), .CO(n289), .S(n290) );
  HADDX1 U257 ( .A0(n311), .B0(n359), .C1(n291), .SO(n292) );
  FADDX1 U258 ( .A(n371), .B(n360), .CI(n382), .CO(n293), .S(n294) );
  HADDX1 U259 ( .A0(n312), .B0(n372), .C1(n295), .SO(n296) );
  OAI22X1 U260 ( .IN1(n494), .IN2(n482), .IN3(n488), .IN4(n398), .QN(n308) );
  AO21X1 U261 ( .IN1(n482), .IN2(n488), .IN3(n386), .Q(n314) );
  OAI22X1 U262 ( .IN1(n482), .IN2(n387), .IN3(n488), .IN4(n386), .QN(n187) );
  OAI22X1 U263 ( .IN1(n488), .IN2(n387), .IN3(n482), .IN4(n388), .QN(n315) );
  OAI22X1 U264 ( .IN1(n488), .IN2(n388), .IN3(n482), .IN4(n389), .QN(n316) );
  OAI22X1 U265 ( .IN1(n488), .IN2(n389), .IN3(n482), .IN4(n390), .QN(n317) );
  OAI22X1 U266 ( .IN1(n482), .IN2(n391), .IN3(n488), .IN4(n390), .QN(n318) );
  OAI22X1 U267 ( .IN1(n488), .IN2(n391), .IN3(n482), .IN4(n392), .QN(n319) );
  OAI22X1 U268 ( .IN1(n482), .IN2(n393), .IN3(n488), .IN4(n392), .QN(n320) );
  OAI22X1 U269 ( .IN1(n488), .IN2(n393), .IN3(n482), .IN4(n394), .QN(n321) );
  OAI22X1 U270 ( .IN1(n482), .IN2(n395), .IN3(n488), .IN4(n394), .QN(n235) );
  OAI22X1 U271 ( .IN1(n488), .IN2(n395), .IN3(n482), .IN4(n396), .QN(n322) );
  OAI22X1 U272 ( .IN1(n482), .IN2(n397), .IN3(n488), .IN4(n396), .QN(n323) );
  XNOR2X1 U283 ( .IN1(n472), .IN2(n500), .Q(n394) );
  XNOR2X1 U286 ( .IN1(n624), .IN2(n500), .Q(n397) );
  OAI22X1 U289 ( .IN1(n495), .IN2(n483), .IN3(n489), .IN4(n411), .QN(n309) );
  AO21X1 U290 ( .IN1(n483), .IN2(n489), .IN3(n399), .Q(n325) );
  OAI22X1 U291 ( .IN1(n483), .IN2(n400), .IN3(n489), .IN4(n399), .QN(n193) );
  OAI22X1 U293 ( .IN1(n489), .IN2(n401), .IN3(n483), .IN4(n402), .QN(n327) );
  OAI22X1 U296 ( .IN1(n489), .IN2(n404), .IN3(n483), .IN4(n405), .QN(n330) );
  OAI22X1 U299 ( .IN1(n483), .IN2(n408), .IN3(n489), .IN4(n407), .QN(n333) );
  OAI22X1 U300 ( .IN1(n489), .IN2(n408), .IN3(n483), .IN4(n409), .QN(n334) );
  OAI22X1 U301 ( .IN1(n483), .IN2(n410), .IN3(n489), .IN4(n409), .QN(n335) );
  XNOR2X1 U312 ( .IN1(n472), .IN2(n501), .Q(n407) );
  XNOR2X1 U315 ( .IN1(n673), .IN2(n501), .Q(n410) );
  OAI22X1 U318 ( .IN1(n496), .IN2(n484), .IN3(n490), .IN4(n424), .QN(n310) );
  AO21X1 U319 ( .IN1(n484), .IN2(n490), .IN3(n412), .Q(n337) );
  OAI22X1 U320 ( .IN1(n484), .IN2(n413), .IN3(n490), .IN4(n412), .QN(n203) );
  OAI22X1 U325 ( .IN1(n490), .IN2(n417), .IN3(n484), .IN4(n418), .QN(n342) );
  OAI22X1 U326 ( .IN1(n484), .IN2(n419), .IN3(n490), .IN4(n418), .QN(n343) );
  OAI22X1 U328 ( .IN1(n484), .IN2(n421), .IN3(n490), .IN4(n420), .QN(n345) );
  OAI22X1 U329 ( .IN1(n490), .IN2(n421), .IN3(n484), .IN4(n422), .QN(n346) );
  OAI22X1 U330 ( .IN1(n484), .IN2(n423), .IN3(n490), .IN4(n422), .QN(n347) );
  XNOR2X1 U341 ( .IN1(n472), .IN2(n502), .Q(n420) );
  XNOR2X1 U344 ( .IN1(n624), .IN2(n502), .Q(n423) );
  OAI22X1 U347 ( .IN1(n497), .IN2(n485), .IN3(n491), .IN4(n437), .QN(n311) );
  AO21X1 U348 ( .IN1(n485), .IN2(n491), .IN3(n425), .Q(n349) );
  OAI22X1 U349 ( .IN1(n485), .IN2(n426), .IN3(n491), .IN4(n425), .QN(n217) );
  OAI22X1 U350 ( .IN1(n491), .IN2(n426), .IN3(n485), .IN4(n427), .QN(n350) );
  OAI22X1 U351 ( .IN1(n491), .IN2(n427), .IN3(n485), .IN4(n428), .QN(n351) );
  OAI22X1 U354 ( .IN1(n491), .IN2(n430), .IN3(n485), .IN4(n431), .QN(n354) );
  OAI22X1 U355 ( .IN1(n485), .IN2(n432), .IN3(n491), .IN4(n431), .QN(n355) );
  OAI22X1 U356 ( .IN1(n491), .IN2(n432), .IN3(n485), .IN4(n433), .QN(n356) );
  OAI22X1 U357 ( .IN1(n485), .IN2(n434), .IN3(n491), .IN4(n433), .QN(n357) );
  OAI22X1 U358 ( .IN1(n491), .IN2(n434), .IN3(n485), .IN4(n435), .QN(n358) );
  OAI22X1 U359 ( .IN1(n485), .IN2(n436), .IN3(n491), .IN4(n435), .QN(n359) );
  XNOR2X1 U370 ( .IN1(n472), .IN2(n672), .Q(n433) );
  XNOR2X1 U373 ( .IN1(n673), .IN2(n672), .Q(n436) );
  OAI22X1 U376 ( .IN1(n498), .IN2(n486), .IN3(n492), .IN4(n450), .QN(n312) );
  AO21X1 U377 ( .IN1(n486), .IN2(n492), .IN3(n438), .Q(n361) );
  OAI22X1 U378 ( .IN1(n486), .IN2(n439), .IN3(n492), .IN4(n438), .QN(n362) );
  OAI22X1 U379 ( .IN1(n492), .IN2(n439), .IN3(n486), .IN4(n440), .QN(n363) );
  OAI22X1 U380 ( .IN1(n492), .IN2(n440), .IN3(n486), .IN4(n441), .QN(n364) );
  OAI22X1 U383 ( .IN1(n492), .IN2(n443), .IN3(n486), .IN4(n444), .QN(n367) );
  OAI22X1 U385 ( .IN1(n492), .IN2(n445), .IN3(n486), .IN4(n446), .QN(n369) );
  OAI22X1 U386 ( .IN1(n486), .IN2(n447), .IN3(n492), .IN4(n446), .QN(n370) );
  OAI22X1 U387 ( .IN1(n492), .IN2(n447), .IN3(n486), .IN4(n448), .QN(n371) );
  OAI22X1 U388 ( .IN1(n486), .IN2(n449), .IN3(n492), .IN4(n448), .QN(n372) );
  XNOR2X1 U399 ( .IN1(n472), .IN2(n670), .Q(n446) );
  OAI22X1 U405 ( .IN1(n499), .IN2(n487), .IN3(n517), .IN4(n463), .QN(n313) );
  AO21X1 U406 ( .IN1(n487), .IN2(n517), .IN3(n451), .Q(n374) );
  OAI22X1 U407 ( .IN1(n487), .IN2(n452), .IN3(n517), .IN4(n451), .QN(n375) );
  OAI22X1 U408 ( .IN1(n517), .IN2(n452), .IN3(n487), .IN4(n453), .QN(n376) );
  OAI22X1 U409 ( .IN1(n517), .IN2(n453), .IN3(n487), .IN4(n454), .QN(n377) );
  OAI22X1 U412 ( .IN1(n517), .IN2(n456), .IN3(n487), .IN4(n457), .QN(n380) );
  OAI22X1 U413 ( .IN1(n487), .IN2(n458), .IN3(n517), .IN4(n457), .QN(n381) );
  OAI22X1 U414 ( .IN1(n517), .IN2(n458), .IN3(n487), .IN4(n459), .QN(n382) );
  OAI22X1 U415 ( .IN1(n487), .IN2(n460), .IN3(n517), .IN4(n459), .QN(n383) );
  OAI22X1 U416 ( .IN1(n517), .IN2(n460), .IN3(n487), .IN4(n461), .QN(n384) );
  OAI22X1 U417 ( .IN1(n487), .IN2(n462), .IN3(n517), .IN4(n461), .QN(n385) );
  XNOR2X1 U426 ( .IN1(n472), .IN2(n505), .Q(n459) );
  XOR2X1 U468 ( .IN1(n500), .IN2(b[10]), .Q(n476) );
  XOR2X1 U471 ( .IN1(n501), .IN2(b[8]), .Q(n477) );
  XOR2X1 U474 ( .IN1(n502), .IN2(b[6]), .Q(n478) );
  XOR2X1 U477 ( .IN1(n671), .IN2(b[4]), .Q(n479) );
  XOR2X1 U480 ( .IN1(n670), .IN2(b[2]), .Q(n480) );
  XOR2X1 U483 ( .IN1(n505), .IN2(b[0]), .Q(n481) );
  XOR3X1 U487 ( .IN1(n254), .IN2(n263), .IN3(n261), .Q(n562) );
  NAND2X0 U488 ( .IN1(n220), .IN2(n227), .QN(n563) );
  NAND2X0 U489 ( .IN1(n254), .IN2(n261), .QN(n618) );
  NAND2X0 U490 ( .IN1(n665), .IN2(n666), .QN(n564) );
  OR2X2 U491 ( .IN1(n195), .IN2(n192), .Q(n665) );
  NBUFFX4 U492 ( .INP(n1), .Z(n624) );
  NBUFFX4 U493 ( .INP(n1), .Z(n673) );
  NOR2X0 U494 ( .IN1(n206), .IN2(n211), .QN(n565) );
  XOR2X2 U495 ( .IN1(n650), .IN2(n251), .Q(n566) );
  XNOR2X2 U496 ( .IN1(n468), .IN2(n670), .Q(n442) );
  XNOR2X2 U497 ( .IN1(n468), .IN2(n502), .Q(n416) );
  XNOR2X2 U498 ( .IN1(n468), .IN2(n505), .Q(n455) );
  XNOR2X2 U499 ( .IN1(n468), .IN2(n500), .Q(n390) );
  XNOR2X2 U500 ( .IN1(n468), .IN2(n501), .Q(n403) );
  INVX0 U501 ( .INP(n471), .ZN(n567) );
  INVX0 U502 ( .INP(n567), .ZN(n568) );
  INVX0 U503 ( .INP(n575), .ZN(n569) );
  XNOR2X2 U504 ( .IN1(n568), .IN2(n505), .Q(n458) );
  XNOR2X2 U505 ( .IN1(n471), .IN2(n670), .Q(n445) );
  XNOR2X2 U506 ( .IN1(n471), .IN2(n502), .Q(n419) );
  XOR2X1 U507 ( .IN1(n368), .IN2(n287), .Q(n570) );
  XOR2X1 U508 ( .IN1(n570), .IN2(n282), .Q(n280) );
  NAND2X0 U509 ( .IN1(n287), .IN2(n282), .QN(n571) );
  NAND2X0 U510 ( .IN1(n368), .IN2(n282), .QN(n572) );
  NAND2X0 U511 ( .IN1(n368), .IN2(n287), .QN(n573) );
  NAND3X0 U512 ( .IN1(n571), .IN2(n573), .IN3(n572), .QN(n279) );
  OAI22X2 U513 ( .IN1(n486), .IN2(n445), .IN3(n492), .IN4(n444), .QN(n368) );
  XOR2X2 U514 ( .IN1(n117), .IN2(n16), .Q(product[12]) );
  OAI22X2 U515 ( .IN1(n487), .IN2(n456), .IN3(n517), .IN4(n455), .QN(n379) );
  OAI22X2 U516 ( .IN1(n517), .IN2(n454), .IN3(n487), .IN4(n455), .QN(n378) );
  OAI22X1 U517 ( .IN1(n491), .IN2(n428), .IN3(n485), .IN4(n429), .QN(n352) );
  NAND2X0 U518 ( .IN1(n211), .IN2(n206), .QN(n574) );
  INVX0 U519 ( .INP(n466), .ZN(n575) );
  INVX0 U520 ( .INP(n575), .ZN(n576) );
  XOR3X1 U521 ( .IN1(n346), .IN2(n336), .IN3(n356), .Q(n278) );
  NAND2X0 U522 ( .IN1(n346), .IN2(n336), .QN(n577) );
  NAND2X0 U523 ( .IN1(n346), .IN2(n356), .QN(n578) );
  NAND2X0 U524 ( .IN1(n336), .IN2(n356), .QN(n579) );
  NAND3X0 U525 ( .IN1(n577), .IN2(n578), .IN3(n579), .QN(n277) );
  XOR2X1 U526 ( .IN1(n355), .IN2(n366), .Q(n580) );
  XOR2X2 U527 ( .IN1(n580), .IN2(n277), .Q(n268) );
  NAND2X0 U528 ( .IN1(n355), .IN2(n366), .QN(n581) );
  NAND2X0 U529 ( .IN1(n355), .IN2(n277), .QN(n582) );
  NAND2X0 U530 ( .IN1(n366), .IN2(n277), .QN(n583) );
  NAND3X0 U531 ( .IN1(n581), .IN2(n582), .IN3(n583), .QN(n267) );
  XNOR2X2 U532 ( .IN1(n471), .IN2(n500), .Q(n393) );
  XOR3X1 U533 ( .IN1(n225), .IN2(n320), .IN3(n216), .Q(n214) );
  NAND2X1 U534 ( .IN1(n225), .IN2(n320), .QN(n584) );
  NAND2X0 U535 ( .IN1(n225), .IN2(n216), .QN(n585) );
  NAND2X0 U536 ( .IN1(n320), .IN2(n216), .QN(n586) );
  NAND3X1 U537 ( .IN1(n584), .IN2(n585), .IN3(n586), .QN(n213) );
  XOR2X2 U538 ( .IN1(n208), .IN2(n215), .Q(n587) );
  XOR2X2 U539 ( .IN1(n587), .IN2(n213), .Q(n206) );
  NAND2X0 U540 ( .IN1(n215), .IN2(n208), .QN(n588) );
  NAND2X0 U541 ( .IN1(n213), .IN2(n208), .QN(n589) );
  NAND2X0 U542 ( .IN1(n215), .IN2(n213), .QN(n590) );
  NAND3X0 U543 ( .IN1(n588), .IN2(n589), .IN3(n590), .QN(n205) );
  NAND3X0 U544 ( .IN1(n617), .IN2(n618), .IN3(n619), .QN(n249) );
  NAND3X0 U545 ( .IN1(n647), .IN2(n648), .IN3(n649), .QN(n251) );
  OAI22X1 U546 ( .IN1(n483), .IN2(n406), .IN3(n489), .IN4(n405), .QN(n331) );
  XOR3X1 U547 ( .IN1(n229), .IN2(n224), .IN3(n222), .Q(n220) );
  XOR2X1 U548 ( .IN1(n148), .IN2(n21), .Q(product[7]) );
  AOI21X1 U549 ( .IN1(n131), .IN2(n118), .IN3(n597), .QN(n117) );
  OAI22X2 U550 ( .IN1(n491), .IN2(n428), .IN3(n485), .IN4(n429), .QN(n591) );
  XNOR2X2 U551 ( .IN1(n471), .IN2(n501), .Q(n406) );
  XNOR2X1 U552 ( .IN1(n592), .IN2(n8), .Q(product[20]) );
  AO21X1 U553 ( .IN1(n54), .IN2(n645), .IN3(n55), .Q(n592) );
  INVX0 U554 ( .INP(n92), .ZN(n593) );
  XOR2X2 U555 ( .IN1(n140), .IN2(n20), .Q(product[8]) );
  INVX0 U556 ( .INP(n75), .ZN(n594) );
  XOR2X1 U557 ( .IN1(n595), .IN2(n596), .Q(product[22]) );
  AO21X1 U558 ( .IN1(n645), .IN2(n32), .IN3(n33), .Q(n595) );
  AND2X2 U559 ( .IN1(n171), .IN2(n30), .Q(n596) );
  OAI22X2 U560 ( .IN1(n489), .IN2(n402), .IN3(n483), .IN4(n403), .QN(n328) );
  OAI21X2 U561 ( .IN1(n628), .IN2(n93), .IN3(n574), .QN(n84) );
  INVX0 U562 ( .INP(n121), .ZN(n597) );
  XOR2X1 U563 ( .IN1(n630), .IN2(n230), .Q(n228) );
  XOR2X2 U564 ( .IN1(n126), .IN2(n17), .Q(product[11]) );
  XNOR3X1 U565 ( .IN1(n598), .IN2(n363), .IN3(n352), .Q(n244) );
  OA22X1 U566 ( .IN1(n489), .IN2(n406), .IN3(n483), .IN4(n407), .Q(n598) );
  AOI21X1 U567 ( .IN1(n78), .IN2(n91), .IN3(n79), .QN(n599) );
  AND2X1 U568 ( .IN1(n258), .IN2(n265), .Q(n600) );
  OAI22X2 U569 ( .IN1(n490), .IN2(n413), .IN3(n484), .IN4(n414), .QN(n338) );
  XOR2X2 U570 ( .IN1(n634), .IN2(n232), .Q(n230) );
  INVX0 U571 ( .INP(n132), .ZN(n601) );
  OAI22X2 U572 ( .IN1(n489), .IN2(n406), .IN3(n483), .IN4(n407), .QN(n602) );
  NAND3X0 U573 ( .IN1(n632), .IN2(n633), .IN3(n631), .QN(n603) );
  XOR3X1 U574 ( .IN1(n221), .IN2(n223), .IN3(n214), .Q(n604) );
  NAND2X0 U575 ( .IN1(n178), .IN2(n97), .QN(n13) );
  NOR2X0 U576 ( .IN1(n205), .IN2(n200), .QN(n605) );
  INVX0 U577 ( .INP(n116), .ZN(n606) );
  INVX0 U578 ( .INP(n606), .ZN(n607) );
  AND2X1 U579 ( .IN1(n195), .IN2(n192), .Q(n608) );
  NOR2X0 U580 ( .IN1(n219), .IN2(n212), .QN(n609) );
  XNOR2X2 U581 ( .IN1(n466), .IN2(n502), .Q(n414) );
  OAI22X2 U582 ( .IN1(n489), .IN2(n400), .IN3(n483), .IN4(n401), .QN(n326) );
  XOR3X1 U583 ( .IN1(n264), .IN2(n354), .IN3(n269), .Q(n260) );
  NAND2X0 U584 ( .IN1(n264), .IN2(n354), .QN(n610) );
  NAND2X0 U585 ( .IN1(n264), .IN2(n269), .QN(n611) );
  NAND2X0 U586 ( .IN1(n354), .IN2(n269), .QN(n612) );
  NAND3X0 U587 ( .IN1(n610), .IN2(n611), .IN3(n612), .QN(n259) );
  XOR2X1 U588 ( .IN1(n252), .IN2(n250), .Q(n613) );
  XOR2X2 U589 ( .IN1(n613), .IN2(n259), .Q(n248) );
  NAND2X0 U590 ( .IN1(n252), .IN2(n562), .QN(n614) );
  NAND2X0 U591 ( .IN1(n252), .IN2(n259), .QN(n615) );
  NAND2X0 U592 ( .IN1(n562), .IN2(n259), .QN(n616) );
  NAND3X0 U593 ( .IN1(n614), .IN2(n615), .IN3(n616), .QN(n247) );
  XNOR2X2 U594 ( .IN1(n474), .IN2(n670), .Q(n448) );
  XNOR2X2 U595 ( .IN1(n474), .IN2(n500), .Q(n396) );
  XNOR2X2 U596 ( .IN1(n474), .IN2(n672), .Q(n435) );
  XNOR2X2 U597 ( .IN1(n474), .IN2(n502), .Q(n422) );
  XNOR2X2 U598 ( .IN1(n474), .IN2(n501), .Q(n409) );
  XOR3X1 U599 ( .IN1(n254), .IN2(n263), .IN3(n261), .Q(n250) );
  NAND2X0 U600 ( .IN1(n254), .IN2(n263), .QN(n617) );
  NAND2X0 U601 ( .IN1(n263), .IN2(n261), .QN(n619) );
  XOR2X1 U602 ( .IN1(n242), .IN2(n240), .Q(n620) );
  XOR2X2 U603 ( .IN1(n620), .IN2(n249), .Q(n238) );
  NAND2X0 U604 ( .IN1(n242), .IN2(n566), .QN(n621) );
  NAND2X0 U605 ( .IN1(n242), .IN2(n249), .QN(n622) );
  NAND2X0 U606 ( .IN1(n566), .IN2(n249), .QN(n623) );
  NAND3X0 U607 ( .IN1(n621), .IN2(n622), .IN3(n623), .QN(n237) );
  XNOR2X2 U608 ( .IN1(n474), .IN2(n505), .Q(n461) );
  OAI22X2 U609 ( .IN1(n420), .IN2(n484), .IN3(n490), .IN4(n419), .QN(n344) );
  NOR2X0 U610 ( .IN1(n266), .IN2(n273), .QN(n625) );
  NAND2X0 U611 ( .IN1(n177), .IN2(n574), .QN(n12) );
  NOR2X0 U612 ( .IN1(n228), .IN2(n237), .QN(n626) );
  NOR2X0 U613 ( .IN1(n248), .IN2(n257), .QN(n627) );
  INVX0 U614 ( .INP(n177), .ZN(n628) );
  INVX0 U615 ( .INP(n565), .ZN(n177) );
  INVX0 U616 ( .INP(n181), .ZN(n629) );
  XOR2X1 U617 ( .IN1(n241), .IN2(n239), .Q(n630) );
  NAND2X0 U618 ( .IN1(n239), .IN2(n230), .QN(n631) );
  NAND2X0 U619 ( .IN1(n241), .IN2(n230), .QN(n632) );
  NAND2X0 U620 ( .IN1(n241), .IN2(n239), .QN(n633) );
  NAND3X0 U621 ( .IN1(n631), .IN2(n632), .IN3(n633), .QN(n227) );
  XOR2X1 U622 ( .IN1(n234), .IN2(n243), .Q(n634) );
  NAND2X0 U623 ( .IN1(n232), .IN2(n243), .QN(n635) );
  NAND2X0 U624 ( .IN1(n234), .IN2(n232), .QN(n636) );
  NAND2X0 U625 ( .IN1(n234), .IN2(n243), .QN(n637) );
  NAND3X0 U626 ( .IN1(n635), .IN2(n637), .IN3(n636), .QN(n229) );
  XOR3X1 U627 ( .IN1(n341), .IN2(n245), .IN3(n331), .Q(n232) );
  NAND2X0 U628 ( .IN1(n331), .IN2(n341), .QN(n638) );
  NAND2X0 U629 ( .IN1(n245), .IN2(n341), .QN(n639) );
  NAND2X1 U630 ( .IN1(n245), .IN2(n331), .QN(n640) );
  NAND3X0 U631 ( .IN1(n638), .IN2(n640), .IN3(n639), .QN(n231) );
  AND2X1 U632 ( .IN1(n220), .IN2(n603), .Q(n641) );
  XOR3X1 U633 ( .IN1(n221), .IN2(n223), .IN3(n214), .Q(n212) );
  NAND2X0 U634 ( .IN1(n221), .IN2(n214), .QN(n642) );
  NAND2X0 U635 ( .IN1(n223), .IN2(n214), .QN(n643) );
  NAND2X0 U636 ( .IN1(n223), .IN2(n221), .QN(n644) );
  NAND3X0 U637 ( .IN1(n642), .IN2(n644), .IN3(n643), .QN(n211) );
  NOR2X0 U638 ( .IN1(n206), .IN2(n211), .QN(n85) );
  OAI22X2 U639 ( .IN1(n483), .IN2(n404), .IN3(n489), .IN4(n403), .QN(n329) );
  OAI22X1 U640 ( .IN1(n490), .IN2(n414), .IN3(n484), .IN4(n415), .QN(n339) );
  XNOR2X2 U641 ( .IN1(n470), .IN2(n505), .Q(n457) );
  XNOR2X2 U642 ( .IN1(n470), .IN2(n670), .Q(n444) );
  OAI21X2 U643 ( .IN1(n104), .IN2(n132), .IN3(n105), .QN(n645) );
  OAI21X2 U644 ( .IN1(n104), .IN2(n132), .IN3(n105), .QN(n646) );
  XOR3X1 U645 ( .IN1(n353), .IN2(n256), .IN3(n343), .Q(n252) );
  NAND2X0 U646 ( .IN1(n353), .IN2(n256), .QN(n647) );
  NAND2X0 U647 ( .IN1(n353), .IN2(n343), .QN(n648) );
  NAND2X1 U648 ( .IN1(n256), .IN2(n343), .QN(n649) );
  XOR2X2 U649 ( .IN1(n244), .IN2(n253), .Q(n650) );
  XOR2X2 U650 ( .IN1(n650), .IN2(n251), .Q(n240) );
  NAND2X0 U651 ( .IN1(n253), .IN2(n244), .QN(n651) );
  NAND2X0 U652 ( .IN1(n251), .IN2(n244), .QN(n652) );
  NAND2X0 U653 ( .IN1(n253), .IN2(n251), .QN(n653) );
  NAND3X0 U654 ( .IN1(n651), .IN2(n652), .IN3(n653), .QN(n239) );
  NAND2X0 U655 ( .IN1(n222), .IN2(n229), .QN(n654) );
  NAND2X0 U656 ( .IN1(n224), .IN2(n229), .QN(n655) );
  NAND2X1 U657 ( .IN1(n224), .IN2(n222), .QN(n656) );
  NAND3X0 U658 ( .IN1(n654), .IN2(n656), .IN3(n655), .QN(n219) );
  OAI22X2 U659 ( .IN1(n490), .IN2(n415), .IN3(n484), .IN4(n416), .QN(n340) );
  OAI22X2 U660 ( .IN1(n485), .IN2(n430), .IN3(n491), .IN4(n429), .QN(n353) );
  INVX0 U661 ( .INP(n609), .ZN(n178) );
  INVX0 U662 ( .INP(n93), .ZN(n657) );
  OAI22X2 U663 ( .IN1(n486), .IN2(n443), .IN3(n492), .IN4(n442), .QN(n366) );
  OAI22X2 U664 ( .IN1(n492), .IN2(n441), .IN3(n486), .IN4(n442), .QN(n365) );
  XOR2X2 U665 ( .IN1(n40), .IN2(n7), .Q(product[21]) );
  XOR2X2 U666 ( .IN1(n658), .IN2(n659), .Q(product[19]) );
  AO21X1 U667 ( .IN1(n645), .IN2(n65), .IN3(n66), .Q(n658) );
  AND2X4 U668 ( .IN1(n665), .IN2(n63), .Q(n659) );
  NOR2X0 U669 ( .IN1(n238), .IN2(n247), .QN(n113) );
  OAI22X2 U670 ( .IN1(n484), .IN2(n417), .IN3(n490), .IN4(n416), .QN(n341) );
  XNOR2X2 U671 ( .IN1(n470), .IN2(n501), .Q(n405) );
  XNOR2X2 U672 ( .IN1(n470), .IN2(n502), .Q(n418) );
  XNOR2X2 U673 ( .IN1(n470), .IN2(n500), .Q(n392) );
  XNOR2X2 U674 ( .IN1(n473), .IN2(n670), .Q(n447) );
  XNOR2X2 U675 ( .IN1(n473), .IN2(n672), .Q(n434) );
  XNOR2X2 U676 ( .IN1(n473), .IN2(n501), .Q(n408) );
  XNOR2X2 U677 ( .IN1(n473), .IN2(n500), .Q(n395) );
  XNOR2X2 U678 ( .IN1(n464), .IN2(n500), .Q(n386) );
  XNOR2X2 U679 ( .IN1(n464), .IN2(n501), .Q(n399) );
  XNOR2X2 U680 ( .IN1(n464), .IN2(n502), .Q(n412) );
  XNOR2X2 U681 ( .IN1(n464), .IN2(n670), .Q(n438) );
  XNOR2X2 U682 ( .IN1(n464), .IN2(n671), .Q(n425) );
  XNOR2X2 U683 ( .IN1(n464), .IN2(n505), .Q(n451) );
  XNOR2X2 U684 ( .IN1(n576), .IN2(n500), .Q(n388) );
  XNOR2X2 U685 ( .IN1(n569), .IN2(n501), .Q(n401) );
  XNOR2X2 U686 ( .IN1(n473), .IN2(n505), .Q(n460) );
  XNOR2X2 U687 ( .IN1(n466), .IN2(n670), .Q(n440) );
  XNOR2X2 U688 ( .IN1(n466), .IN2(n671), .Q(n427) );
  XNOR2X2 U689 ( .IN1(n466), .IN2(n505), .Q(n453) );
  XNOR2X2 U690 ( .IN1(n568), .IN2(n672), .Q(n432) );
  XNOR2X2 U691 ( .IN1(n465), .IN2(n500), .Q(n387) );
  XNOR2X2 U692 ( .IN1(n465), .IN2(n502), .Q(n413) );
  XNOR2X2 U693 ( .IN1(n465), .IN2(n501), .Q(n400) );
  XNOR2X2 U694 ( .IN1(n465), .IN2(n505), .Q(n452) );
  XNOR2X2 U695 ( .IN1(n465), .IN2(n670), .Q(n439) );
  XNOR2X2 U696 ( .IN1(n468), .IN2(n672), .Q(n429) );
  XNOR2X2 U697 ( .IN1(n469), .IN2(n500), .Q(n391) );
  XNOR2X2 U698 ( .IN1(n469), .IN2(n670), .Q(n443) );
  XNOR2X2 U699 ( .IN1(n469), .IN2(n505), .Q(n456) );
  XNOR2X2 U700 ( .IN1(n469), .IN2(n501), .Q(n404) );
  XNOR2X2 U701 ( .IN1(n469), .IN2(n672), .Q(n430) );
  XNOR2X2 U702 ( .IN1(n469), .IN2(n502), .Q(n417) );
  XNOR2X2 U703 ( .IN1(n467), .IN2(n502), .Q(n415) );
  XNOR2X2 U704 ( .IN1(n467), .IN2(n501), .Q(n402) );
  XNOR2X2 U705 ( .IN1(n467), .IN2(n500), .Q(n389) );
  XNOR2X2 U706 ( .IN1(n467), .IN2(n505), .Q(n454) );
  XNOR2X2 U707 ( .IN1(n467), .IN2(n670), .Q(n441) );
  XNOR2X2 U708 ( .IN1(n467), .IN2(n672), .Q(n428) );
  NAND2X0 U709 ( .IN1(n45), .IN2(n36), .QN(n34) );
  NAND2X0 U710 ( .IN1(n176), .IN2(n81), .QN(n11) );
  NAND2X0 U711 ( .IN1(n183), .IN2(n130), .QN(n18) );
  NAND2X0 U712 ( .IN1(n45), .IN2(n27), .QN(n25) );
  NOR2X0 U713 ( .IN1(n67), .IN2(n564), .QN(n45) );
  NAND2X0 U714 ( .IN1(n185), .IN2(n139), .QN(n20) );
  NAND2X0 U715 ( .IN1(n36), .IN2(n39), .QN(n7) );
  NAND2X0 U716 ( .IN1(n69), .IN2(n68), .QN(n10) );
  NOR2X0 U717 ( .IN1(n199), .IN2(n196), .QN(n67) );
  INVX0 U718 ( .INP(n4), .ZN(n75) );
  NOR2X0 U719 ( .IN1(n92), .IN2(n628), .QN(n83) );
  INVX0 U720 ( .INP(n605), .ZN(n176) );
  XNOR2X1 U721 ( .IN1(n660), .IN2(n12), .Q(product[16]) );
  AO21X1 U722 ( .IN1(n646), .IN2(n593), .IN3(n657), .Q(n660) );
  NOR2X0 U723 ( .IN1(n120), .IN2(n629), .QN(n111) );
  INVX0 U724 ( .INP(n118), .ZN(n120) );
  NOR2X0 U725 ( .IN1(n85), .IN2(n605), .QN(n78) );
  NAND2X0 U726 ( .IN1(n182), .IN2(n125), .QN(n17) );
  INVX0 U727 ( .INP(n101), .ZN(n99) );
  INVX0 U728 ( .INP(n45), .ZN(n43) );
  INVX0 U729 ( .INP(n625), .ZN(n184) );
  INVX0 U730 ( .INP(n626), .ZN(n180) );
  INVX0 U731 ( .INP(n132), .ZN(n131) );
  NAND2X0 U732 ( .IN1(n99), .IN2(n563), .QN(n14) );
  INVX0 U733 ( .INP(n141), .ZN(n140) );
  NAND2X0 U734 ( .IN1(n181), .IN2(n607), .QN(n16) );
  INVX0 U735 ( .INP(n113), .ZN(n181) );
  NAND2X0 U736 ( .IN1(n180), .IN2(n109), .QN(n15) );
  XNOR2X1 U737 ( .IN1(n661), .IN2(n13), .Q(product[15]) );
  AO21X1 U738 ( .IN1(n646), .IN2(n99), .IN3(n641), .Q(n661) );
  INVX0 U739 ( .INP(n91), .ZN(n93) );
  INVX0 U740 ( .INP(n119), .ZN(n121) );
  INVX0 U741 ( .INP(n46), .ZN(n44) );
  INVX0 U742 ( .INP(n129), .ZN(n183) );
  INVX0 U743 ( .INP(n5), .ZN(n74) );
  NOR2X0 U744 ( .IN1(n266), .IN2(n273), .QN(n135) );
  NAND2X0 U745 ( .IN1(n220), .IN2(n227), .QN(n102) );
  INVX0 U746 ( .INP(n138), .ZN(n185) );
  INVX0 U747 ( .INP(n154), .ZN(n153) );
  INVX0 U748 ( .INP(n29), .ZN(n171) );
  NAND2X0 U749 ( .IN1(n666), .IN2(n52), .QN(n8) );
  NAND2X0 U750 ( .IN1(n258), .IN2(n265), .QN(n130) );
  NAND2X0 U751 ( .IN1(n205), .IN2(n200), .QN(n81) );
  NOR2X0 U752 ( .IN1(n228), .IN2(n237), .QN(n108) );
  NAND2X0 U753 ( .IN1(n228), .IN2(n237), .QN(n109) );
  NAND2X0 U754 ( .IN1(n266), .IN2(n273), .QN(n136) );
  NOR2X0 U755 ( .IN1(n220), .IN2(n603), .QN(n101) );
  NAND2X0 U756 ( .IN1(n247), .IN2(n238), .QN(n116) );
  INVX0 U757 ( .INP(n67), .ZN(n69) );
  NAND2X0 U758 ( .IN1(n219), .IN2(n212), .QN(n97) );
  NAND2X0 U759 ( .IN1(n257), .IN2(n248), .QN(n125) );
  NAND2X0 U760 ( .IN1(n184), .IN2(n136), .QN(n19) );
  NOR2X0 U761 ( .IN1(n625), .IN2(n138), .QN(n133) );
  OA21X1 U762 ( .IN1(n662), .IN2(n663), .IN3(n664), .Q(n154) );
  OR2X1 U763 ( .IN1(n157), .IN2(n159), .Q(n662) );
  OA21X1 U764 ( .IN1(n162), .IN2(n164), .IN3(n163), .Q(n663) );
  OA21X1 U765 ( .IN1(n160), .IN2(n157), .IN3(n158), .Q(n664) );
  INVX0 U766 ( .INP(n147), .ZN(n145) );
  INVX0 U767 ( .INP(n68), .ZN(n70) );
  INVX0 U768 ( .INP(n39), .ZN(n37) );
  INVX0 U769 ( .INP(n38), .ZN(n36) );
  NOR2X0 U770 ( .IN1(n38), .IN2(n29), .QN(n27) );
  INVX0 U771 ( .INP(n52), .ZN(n50) );
  NOR2X0 U772 ( .IN1(n274), .IN2(n279), .QN(n138) );
  NOR2X0 U773 ( .IN1(n290), .IN2(n293), .QN(n157) );
  NOR2X0 U774 ( .IN1(n294), .IN2(n295), .QN(n159) );
  NAND2X0 U775 ( .IN1(n274), .IN2(n279), .QN(n139) );
  OR2X1 U776 ( .IN1(n191), .IN2(n190), .Q(n666) );
  NAND2X0 U777 ( .IN1(n290), .IN2(n293), .QN(n158) );
  OR2X1 U778 ( .IN1(n280), .IN2(n285), .Q(n667) );
  OR2X1 U779 ( .IN1(n286), .IN2(n289), .Q(n668) );
  AND2X1 U780 ( .IN1(n286), .IN2(n289), .Q(n669) );
  INVX0 U781 ( .INP(n187), .ZN(n188) );
  NAND2X0 U782 ( .IN1(n199), .IN2(n196), .QN(n68) );
  NOR2X0 U783 ( .IN1(n187), .IN2(n314), .QN(n29) );
  NOR2X0 U784 ( .IN1(n189), .IN2(n188), .QN(n38) );
  NAND2X0 U785 ( .IN1(n189), .IN2(n188), .QN(n39) );
  NAND2X0 U786 ( .IN1(n294), .IN2(n295), .QN(n160) );
  NOR2X0 U787 ( .IN1(n296), .IN2(n383), .QN(n162) );
  NOR2X0 U788 ( .IN1(n384), .IN2(n373), .QN(n167) );
  NAND2X0 U789 ( .IN1(n384), .IN2(n373), .QN(n168) );
  NAND2X0 U790 ( .IN1(n296), .IN2(n383), .QN(n163) );
  OA21X1 U791 ( .IN1(n167), .IN2(n170), .IN3(n168), .Q(n164) );
  NAND2X0 U792 ( .IN1(n187), .IN2(n314), .QN(n30) );
  OR2X1 U793 ( .IN1(n624), .IN2(n498), .Q(n450) );
  INVX0 U794 ( .INP(n235), .ZN(n236) );
  AND2X1 U795 ( .IN1(n673), .IN2(n301), .Q(n348) );
  INVX0 U796 ( .INP(n203), .ZN(n204) );
  OR2X1 U797 ( .IN1(n673), .IN2(n494), .Q(n398) );
  OR2X1 U798 ( .IN1(n673), .IN2(n495), .Q(n411) );
  OR2X1 U799 ( .IN1(n624), .IN2(n496), .Q(n424) );
  OR2X1 U800 ( .IN1(n624), .IN2(n497), .Q(n437) );
  AND2X1 U801 ( .IN1(n624), .IN2(n299), .Q(n336) );
  INVX0 U802 ( .INP(n217), .ZN(n218) );
  AND2X1 U803 ( .IN1(n673), .IN2(n297), .Q(n324) );
  AND2X1 U804 ( .IN1(n624), .IN2(n303), .Q(n360) );
  INVX0 U805 ( .INP(n193), .ZN(n194) );
  XNOR2X1 U806 ( .IN1(n673), .IN2(n670), .Q(n449) );
  AND2X1 U807 ( .IN1(n673), .IN2(n305), .Q(n373) );
  INVX0 U808 ( .INP(n492), .ZN(n305) );
  NAND2X0 U809 ( .IN1(n385), .IN2(n313), .QN(n170) );
  OR2X1 U810 ( .IN1(n624), .IN2(n499), .Q(n463) );
  INVX0 U811 ( .INP(n670), .ZN(n498) );
  INVX0 U812 ( .INP(n671), .ZN(n497) );
  INVX0 U813 ( .INP(n490), .ZN(n301) );
  INVX0 U814 ( .INP(n491), .ZN(n303) );
  INVX0 U815 ( .INP(n489), .ZN(n299) );
  INVX0 U816 ( .INP(n488), .ZN(n297) );
  XNOR2X1 U817 ( .IN1(n673), .IN2(n505), .Q(n462) );
  NBUFFX2 U818 ( .INP(n503), .Z(n672) );
  NBUFFX2 U819 ( .INP(n503), .Z(n671) );
  NBUFFX4 U820 ( .INP(n504), .Z(n670) );
  XNOR2X1 U821 ( .IN1(b[6]), .IN2(n671), .Q(n490) );
  XNOR2X1 U822 ( .IN1(n670), .IN2(b[4]), .Q(n491) );
  XNOR2X1 U823 ( .IN1(n505), .IN2(b[2]), .Q(n492) );
  XNOR2X1 U824 ( .IN1(n501), .IN2(b[10]), .Q(n488) );
  XNOR2X1 U825 ( .IN1(n502), .IN2(b[8]), .Q(n489) );
  NAND2X0 U826 ( .IN1(n490), .IN2(n478), .QN(n484) );
  NAND2X0 U827 ( .IN1(n489), .IN2(n477), .QN(n483) );
  NAND2X0 U828 ( .IN1(n491), .IN2(n479), .QN(n485) );
  NAND2X0 U829 ( .IN1(n488), .IN2(n476), .QN(n482) );
  NAND2X1 U830 ( .IN1(n492), .IN2(n480), .QN(n486) );
  INVX0 U831 ( .INP(b[0]), .ZN(n517) );
  NAND2X1 U832 ( .IN1(n481), .IN2(n517), .QN(n487) );
  INVX0 U833 ( .INP(n502), .ZN(n496) );
  INVX0 U834 ( .INP(n501), .ZN(n495) );
  INVX0 U835 ( .INP(n500), .ZN(n494) );
  INVX0 U836 ( .INP(n505), .ZN(n499) );
  NAND2X0 U837 ( .IN1(n665), .IN2(n666), .QN(n47) );
  NAND2X0 U838 ( .IN1(n69), .IN2(n665), .QN(n56) );
  NAND2X0 U839 ( .IN1(n211), .IN2(n206), .QN(n88) );
  NOR2X0 U840 ( .IN1(n627), .IN2(n129), .QN(n118) );
  INVX0 U841 ( .INP(n627), .ZN(n182) );
  NOR2X0 U842 ( .IN1(n258), .IN2(n265), .QN(n129) );
  NAND2X0 U843 ( .IN1(n191), .IN2(n190), .QN(n52) );
  INVX0 U844 ( .INP(n90), .ZN(n92) );
  NAND2X0 U845 ( .IN1(n90), .IN2(n78), .QN(n5) );
  NOR2X0 U846 ( .IN1(n101), .IN2(n609), .QN(n90) );
  NOR2X0 U847 ( .IN1(n248), .IN2(n257), .QN(n124) );
  NAND2X0 U848 ( .IN1(n106), .IN2(n118), .QN(n104) );
  NOR2X0 U849 ( .IN1(n626), .IN2(n113), .QN(n106) );
  NAND2X0 U850 ( .IN1(n195), .IN2(n192), .QN(n63) );
  XNOR2X2 U851 ( .IN1(n470), .IN2(n672), .Q(n431) );
  NOR2X0 U852 ( .IN1(n5), .IN2(n25), .QN(n23) );
  NOR2X0 U853 ( .IN1(n5), .IN2(n34), .QN(n32) );
  NOR2X0 U854 ( .IN1(n5), .IN2(n56), .QN(n54) );
  NOR2X0 U855 ( .IN1(n5), .IN2(n43), .QN(n41) );
  NOR2X0 U856 ( .IN1(n5), .IN2(n67), .QN(n65) );
  NOR2X0 U857 ( .IN1(n219), .IN2(n604), .QN(n96) );
  XNOR2X2 U858 ( .IN1(n465), .IN2(n671), .Q(n426) );
  XNOR2X2 U859 ( .IN1(n473), .IN2(n502), .Q(n421) );
  NAND2X0 U860 ( .IN1(n667), .IN2(n147), .QN(n21) );
  NAND2X0 U861 ( .IN1(n667), .IN2(n668), .QN(n142) );
  NAND2X0 U862 ( .IN1(n280), .IN2(n285), .QN(n147) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1 ( in_a, in_b, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [11:0] \output ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [23:7] pre_out;
  wire   [11:0] rnd_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1_DW01_inc_2 add_37_round ( .A({
        n1, pre_out[18:7]}), .SUM({rnd_out, SYNOPSYS_UNCONNECTED__0}) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1_DW_mult_tc_7 mult_35 ( .a(in_a), 
        .b(in_b), .product({pre_out, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7}) );
  AO21X2 U2 ( .IN1(rnd_out[6]), .IN2(n11), .IN3(n3), .Q(\output [6]) );
  INVX0 U3 ( .INP(pre_out[23]), .ZN(n10) );
  AO21X2 U4 ( .IN1(rnd_out[0]), .IN2(n4), .IN3(n3), .Q(\output [0]) );
  AO21X2 U5 ( .IN1(rnd_out[7]), .IN2(n4), .IN3(n3), .Q(\output [7]) );
  AO22X2 U6 ( .IN1(pre_out[23]), .IN2(n2), .IN3(n4), .IN4(rnd_out[11]), .Q(
        \output [11]) );
  AND2X1 U7 ( .IN1(n12), .IN2(n10), .Q(n5) );
  AO21X2 U8 ( .IN1(rnd_out[1]), .IN2(n11), .IN3(n3), .Q(\output [1]) );
  AND2X1 U9 ( .IN1(n12), .IN2(n10), .Q(n3) );
  AO21X1 U10 ( .IN1(rnd_out[2]), .IN2(n4), .IN3(n5), .Q(\output [2]) );
  AO21X1 U11 ( .IN1(rnd_out[8]), .IN2(n4), .IN3(n5), .Q(\output [8]) );
  DELLN1X2 U12 ( .INP(pre_out[19]), .Z(n1) );
  INVX0 U13 ( .INP(n4), .ZN(n2) );
  INVX0 U14 ( .INP(n12), .ZN(n4) );
  NAND4X0 U15 ( .IN1(pre_out[21]), .IN2(pre_out[20]), .IN3(pre_out[22]), .IN4(
        pre_out[19]), .QN(n8) );
  AO21X1 U16 ( .IN1(rnd_out[10]), .IN2(n11), .IN3(n5), .Q(\output [10]) );
  AO21X1 U17 ( .IN1(rnd_out[9]), .IN2(n11), .IN3(n5), .Q(\output [9]) );
  AO21X1 U18 ( .IN1(rnd_out[3]), .IN2(n11), .IN3(n5), .Q(\output [3]) );
  INVX0 U19 ( .INP(n12), .ZN(n11) );
  NAND2X0 U20 ( .IN1(n7), .IN2(n6), .QN(n9) );
  NOR2X0 U21 ( .IN1(pre_out[20]), .IN2(pre_out[19]), .QN(n6) );
  NOR2X0 U22 ( .IN1(pre_out[21]), .IN2(pre_out[22]), .QN(n7) );
  MUX21X1 U23 ( .IN1(n9), .IN2(n8), .S(pre_out[23]), .Q(n12) );
  AO21X1 U24 ( .IN1(rnd_out[4]), .IN2(n4), .IN3(n5), .Q(\output [4]) );
  AO21X1 U25 ( .IN1(rnd_out[5]), .IN2(n11), .IN3(n3), .Q(\output [5]) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0_DW01_inc_2 ( A, SUM );
  input [12:0] A;
  output [12:0] SUM;
  wire   n1, n2, n5, n7, n8, n10, n11, n12, n13, n14, n15, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n29, n30, n31, n32, n33, n34, n35, n36, n37,
         n38, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79;
  assign n5 = A[11];
  assign n8 = A[10];
  assign n12 = A[9];
  assign n15 = A[8];
  assign n19 = A[7];
  assign n23 = A[6];
  assign n26 = A[5];
  assign n38 = A[1];

  XOR2X1 U1 ( .IN1(n2), .IN2(n1), .Q(SUM[12]) );
  XOR2X1 U13 ( .IN1(n13), .IN2(n14), .Q(SUM[9]) );
  XOR2X1 U27 ( .IN1(n25), .IN2(n24), .Q(SUM[6]) );
  XNOR2X1 U36 ( .IN1(n31), .IN2(n32), .Q(SUM[4]) );
  XOR2X1 U44 ( .IN1(n36), .IN2(n37), .Q(SUM[2]) );
  AND2X4 U54 ( .IN1(A[4]), .IN2(A[3]), .Q(n69) );
  NAND2X0 U55 ( .IN1(n26), .IN2(n23), .QN(n70) );
  NOR2X0 U56 ( .IN1(n74), .IN2(n29), .QN(n71) );
  NAND2X0 U57 ( .IN1(n19), .IN2(n71), .QN(n72) );
  AND2X1 U58 ( .IN1(n71), .IN2(n19), .Q(n77) );
  NOR2X0 U59 ( .IN1(n72), .IN2(n11), .QN(n73) );
  NAND2X0 U60 ( .IN1(n26), .IN2(n23), .QN(n74) );
  NOR2X0 U61 ( .IN1(n70), .IN2(n29), .QN(n75) );
  XOR2X2 U62 ( .IN1(n73), .IN2(n8), .Q(SUM[10]) );
  AND2X4 U63 ( .IN1(n19), .IN2(n15), .Q(n76) );
  AND2X1 U64 ( .IN1(A[4]), .IN2(A[3]), .Q(n30) );
  XNOR2X2 U65 ( .IN1(n75), .IN2(n20), .Q(SUM[7]) );
  AND2X4 U66 ( .IN1(n69), .IN2(n35), .Q(n78) );
  XNOR2X1 U67 ( .IN1(n7), .IN2(n5), .Q(SUM[11]) );
  AND2X1 U68 ( .IN1(n8), .IN2(n5), .Q(n79) );
  XOR2X1 U69 ( .IN1(n33), .IN2(n34), .Q(SUM[3]) );
  XOR2X1 U70 ( .IN1(n26), .IN2(n78), .Q(SUM[5]) );
  INVX0 U71 ( .INP(n19), .ZN(n20) );
  XOR2X1 U72 ( .IN1(n15), .IN2(n77), .Q(SUM[8]) );
  INVX0 U73 ( .INP(n23), .ZN(n24) );
  INVX0 U74 ( .INP(n12), .ZN(n13) );
  XOR2X1 U75 ( .IN1(n38), .IN2(A[0]), .Q(SUM[1]) );
  INVX0 U76 ( .INP(A[2]), .ZN(n36) );
  INVX0 U77 ( .INP(A[12]), .ZN(n1) );
  NOR2X0 U78 ( .IN1(n33), .IN2(n34), .QN(n32) );
  NAND2X0 U79 ( .IN1(n30), .IN2(n35), .QN(n29) );
  INVX0 U80 ( .INP(A[4]), .ZN(n31) );
  NAND2X0 U81 ( .IN1(n26), .IN2(n78), .QN(n25) );
  NAND2X0 U82 ( .IN1(n26), .IN2(n23), .QN(n22) );
  NAND2X0 U83 ( .IN1(n75), .IN2(n76), .QN(n14) );
  NAND2X0 U84 ( .IN1(n38), .IN2(A[0]), .QN(n37) );
  INVX0 U85 ( .INP(n35), .ZN(n34) );
  NOR2X0 U86 ( .IN1(n36), .IN2(n37), .QN(n35) );
  NOR2X0 U87 ( .IN1(n18), .IN2(n11), .QN(n10) );
  NAND2X0 U88 ( .IN1(n19), .IN2(n21), .QN(n18) );
  NAND2X0 U89 ( .IN1(n79), .IN2(n10), .QN(n2) );
  NAND2X0 U90 ( .IN1(n8), .IN2(n10), .QN(n7) );
  NAND2X0 U91 ( .IN1(n12), .IN2(n15), .QN(n11) );
  NOR2X0 U92 ( .IN1(n22), .IN2(n29), .QN(n21) );
  INVX0 U93 ( .INP(A[3]), .ZN(n33) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0_DW_mult_tc_3 ( a, b, 
        product );
  input [11:0] a;
  input [11:0] b;
  output [23:0] product;
  wire   n1, n2, n3, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n21, n22, n23, n24, n26, n28, n30, n31, n32, n33, n34, n35, n36, n37,
         n39, n40, n41, n44, n48, n50, n51, n52, n53, n54, n63, n64, n65, n66,
         n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n81, n82, n83, n84,
         n85, n86, n87, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n101,
         n102, n103, n104, n105, n106, n109, n110, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n126, n127, n128, n132,
         n133, n135, n137, n138, n139, n142, n143, n144, n145, n147, n148,
         n149, n152, n153, n155, n156, n157, n162, n163, n166, n167, n169,
         n170, n171, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n541, n544, n545, n546, n547, n548, n549, n551, n552, n553, n555,
         n557, n558, n559, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847;

  AOI21X1 U6 ( .IN1(n835), .IN2(n21), .IN3(n22), .QN(product[23]) );
  OAI21X1 U8 ( .IN1(n23), .IN2(n2), .IN3(n24), .QN(n22) );
  AOI21X1 U10 ( .IN1(n35), .IN2(n846), .IN3(n26), .QN(n24) );
  OAI21X1 U20 ( .IN1(n32), .IN2(n2), .IN3(n33), .QN(n31) );
  OAI21X1 U24 ( .IN1(n36), .IN2(n44), .IN3(n37), .QN(n35) );
  OAI21X1 U32 ( .IN1(n41), .IN2(n2), .IN3(n44), .QN(n40) );
  OAI21X1 U46 ( .IN1(n52), .IN2(n2), .IN3(n53), .QN(n51) );
  XOR2X1 U55 ( .IN1(n67), .IN2(n8), .Q(product[18]) );
  AOI21X1 U60 ( .IN1(n63), .IN2(n76), .IN3(n64), .QN(n2) );
  OAI21X1 U62 ( .IN1(n65), .IN2(n73), .IN3(n66), .QN(n64) );
  XOR2X1 U67 ( .IN1(n74), .IN2(n9), .Q(product[17]) );
  AOI21X1 U68 ( .IN1(n1), .IN2(n68), .IN3(n69), .QN(n67) );
  OAI21X1 U70 ( .IN1(n711), .IN2(n78), .IN3(n73), .QN(n69) );
  XOR2X1 U77 ( .IN1(n83), .IN2(n10), .Q(product[16]) );
  AOI21X1 U78 ( .IN1(n835), .IN2(n75), .IN3(n715), .QN(n74) );
  OAI21X1 U84 ( .IN1(n87), .IN2(n81), .IN3(n82), .QN(n76) );
  AOI21X1 U90 ( .IN1(n835), .IN2(n84), .IN3(n85), .QN(n83) );
  AOI21X1 U100 ( .IN1(n91), .IN2(n104), .IN3(n92), .QN(n90) );
  OAI21X1 U102 ( .IN1(n101), .IN2(n93), .IN3(n94), .QN(n92) );
  AOI21X1 U108 ( .IN1(n746), .IN2(n96), .IN3(n97), .QN(n95) );
  OAI21X1 U124 ( .IN1(n115), .IN2(n109), .IN3(n110), .QN(n104) );
  XNOR2X1 U137 ( .IN1(n122), .IN2(n16), .Q(product[10]) );
  OAI21X1 U141 ( .IN1(n124), .IN2(n120), .IN3(n121), .QN(n119) );
  XOR2X1 U146 ( .IN1(n698), .IN2(n17), .Q(product[9]) );
  OAI21X1 U147 ( .IN1(n123), .IN2(n698), .IN3(n124), .QN(n122) );
  XOR2X1 U152 ( .IN1(n133), .IN2(n18), .Q(product[8]) );
  OAI21X1 U154 ( .IN1(n127), .IN2(n139), .IN3(n128), .QN(n126) );
  AOI21X1 U156 ( .IN1(n837), .IN2(n135), .IN3(n758), .QN(n128) );
  XNOR2X1 U163 ( .IN1(n138), .IN2(n19), .Q(product[7]) );
  AOI21X1 U164 ( .IN1(n138), .IN2(n838), .IN3(n135), .QN(n133) );
  FADDX1 U191 ( .A(n395), .B(n406), .CI(n178), .CO(n174), .S(n175) );
  FADDX1 U192 ( .A(n179), .B(n184), .CI(n182), .CO(n176), .S(n177) );
  FADDX1 U193 ( .A(n418), .B(n407), .CI(n396), .CO(n178), .S(n179) );
  FADDX1 U195 ( .A(n192), .B(n397), .CI(n185), .CO(n182), .S(n183) );
  FADDX1 U196 ( .A(n419), .B(n408), .CI(n430), .CO(n184), .S(n185) );
  FADDX1 U197 ( .A(n189), .B(n198), .CI(n196), .CO(n186), .S(n187) );
  FADDX1 U198 ( .A(n200), .B(n193), .CI(n191), .CO(n188), .S(n189) );
  FADDX1 U199 ( .A(n398), .B(n442), .CI(n202), .CO(n190), .S(n191) );
  FADDX1 U200 ( .A(n409), .B(n431), .CI(n420), .CO(n192), .S(n193) );
  FADDX1 U201 ( .A(n206), .B(n208), .CI(n197), .CO(n194), .S(n195) );
  FADDX1 U202 ( .A(n210), .B(n201), .CI(n199), .CO(n196), .S(n197) );
  FADDX1 U203 ( .A(n203), .B(n214), .CI(n212), .CO(n198), .S(n199) );
  FADDX1 U204 ( .A(n454), .B(n421), .CI(n399), .CO(n200), .S(n201) );
  FADDX1 U205 ( .A(n432), .B(n443), .CI(n410), .CO(n202), .S(n203) );
  FADDX1 U209 ( .A(n228), .B(n400), .CI(n226), .CO(n210), .S(n211) );
  FADDX1 U210 ( .A(n422), .B(n444), .CI(n466), .CO(n212), .S(n213) );
  FADDX1 U211 ( .A(n433), .B(n455), .CI(n411), .CO(n214), .S(n215) );
  FADDX1 U217 ( .A(n445), .B(n434), .CI(n423), .CO(n226), .S(n227) );
  FADDX1 U218 ( .A(n456), .B(n467), .CI(n608), .CO(n228), .S(n229) );
  FADDX1 U221 ( .A(n254), .B(n256), .CI(n239), .CO(n234), .S(n235) );
  FADDX1 U222 ( .A(n258), .B(n243), .CI(n241), .CO(n236), .S(n237) );
  FADDX1 U224 ( .A(n490), .B(n424), .CI(n402), .CO(n240), .S(n241) );
  FADDX1 U225 ( .A(n468), .B(n457), .CI(n446), .CO(n242), .S(n243) );
  FADDX1 U226 ( .A(n435), .B(n479), .CI(n413), .CO(n244), .S(n245) );
  FADDX1 U230 ( .A(n276), .B(n259), .CI(n257), .CO(n252), .S(n253) );
  FADDX1 U231 ( .A(n263), .B(n278), .CI(n261), .CO(n254), .S(n255) );
  FADDX1 U232 ( .A(n282), .B(n403), .CI(n280), .CO(n256) );
  FADDX1 U234 ( .A(n480), .B(n469), .CI(n447), .CO(n260), .S(n261) );
  FADDX1 U241 ( .A(n300), .B(n302), .CI(n298), .CO(n274), .S(n275) );
  FADDX1 U243 ( .A(n437), .B(n492), .CI(n448), .CO(n278), .S(n279) );
  XNOR2X1 U245 ( .IN1(n459), .IN2(n470), .Q(n283) );
  OR2X1 U246 ( .IN1(n459), .IN2(n470), .Q(n282) );
  FADDX1 U250 ( .A(n301), .B(n314), .CI(n297), .CO(n290), .S(n291) );
  FADDX1 U252 ( .A(n303), .B(n320), .CI(n405), .CO(n294), .S(n295) );
  FADDX1 U253 ( .A(n427), .B(n515), .CI(n526), .CO(n296), .S(n297) );
  FADDX1 U254 ( .A(n504), .B(n482), .CI(n493), .CO(n298), .S(n299) );
  FADDX1 U260 ( .A(n317), .B(n332), .CI(n319), .CO(n310) );
  HADDX1 U265 ( .A0(n483), .B0(n450), .C1(n320), .SO(n321) );
  FADDX1 U266 ( .A(n340), .B(n327), .CI(n325), .CO(n322), .S(n323) );
  FADDX1 U267 ( .A(n342), .B(n344), .CI(n329), .CO(n324), .S(n325) );
  FADDX1 U272 ( .A(n528), .B(n484), .CI(n517), .CO(n334), .S(n335) );
  HADDX1 U273 ( .A0(n451), .B0(n462), .C1(n336), .SO(n337) );
  FADDX1 U277 ( .A(n351), .B(n507), .CI(n362), .CO(n344) );
  FADDX1 U278 ( .A(n474), .B(n485), .CI(n518), .CO(n346), .S(n347) );
  FADDX1 U281 ( .A(n366), .B(n357), .CI(n355), .CO(n352), .S(n353) );
  FADDX1 U282 ( .A(n361), .B(n359), .CI(n368), .CO(n354), .S(n355) );
  FADDX1 U285 ( .A(n530), .B(n497), .CI(n519), .CO(n360), .S(n361) );
  HADDX1 U286 ( .A0(n475), .B0(n453), .C1(n362), .SO(n363) );
  FADDX1 U287 ( .A(n376), .B(n369), .CI(n367), .CO(n364), .S(n365) );
  FADDX1 U288 ( .A(n371), .B(n380), .CI(n378), .CO(n366), .S(n367) );
  FADDX1 U289 ( .A(n498), .B(n520), .CI(n373), .CO(n368), .S(n369) );
  FADDX1 U290 ( .A(n531), .B(n509), .CI(n487), .CO(n370), .S(n371) );
  FADDX1 U292 ( .A(n379), .B(n384), .CI(n377), .CO(n374), .S(n375) );
  FADDX1 U293 ( .A(n381), .B(n532), .CI(n386), .CO(n376), .S(n377) );
  FADDX1 U294 ( .A(n510), .B(n499), .CI(n521), .CO(n378), .S(n379) );
  HADDX1 U295 ( .A0(n488), .B0(n477), .C1(n380), .SO(n381) );
  FADDX1 U296 ( .A(n390), .B(n387), .CI(n385), .CO(n382), .S(n383) );
  FADDX1 U297 ( .A(n511), .B(n533), .CI(n522), .CO(n384), .S(n385) );
  HADDX1 U298 ( .A0(n500), .B0(n489), .C1(n386), .SO(n387) );
  FADDX1 U299 ( .A(n523), .B(n534), .CI(n391), .CO(n388), .S(n389) );
  HADDX1 U300 ( .A0(n512), .B0(n501), .C1(n390), .SO(n391) );
  HADDX1 U301 ( .A0(n535), .B0(n524), .C1(n392), .SO(n393) );
  OR2X1 U303 ( .IN1(n744), .IN2(n732), .Q(n395) );
  OR2X1 U304 ( .IN1(n731), .IN2(n626), .Q(n396) );
  OR2X1 U305 ( .IN1(n732), .IN2(n776), .Q(n397) );
  OR2X1 U306 ( .IN1(n731), .IN2(n722), .Q(n398) );
  OR2X1 U307 ( .IN1(n732), .IN2(n742), .Q(n399) );
  OR2X1 U308 ( .IN1(n731), .IN2(n719), .Q(n400) );
  OR2X1 U309 ( .IN1(n732), .IN2(n759), .Q(n401) );
  OR2X1 U310 ( .IN1(n731), .IN2(n729), .Q(n402) );
  OR2X1 U311 ( .IN1(n549), .IN2(n730), .Q(n403) );
  HADDX2 U471 ( .A0(n476), .B0(n465), .C1(n372), .SO(n373) );
  INVX0 U472 ( .INP(n292), .ZN(n606) );
  INVX0 U473 ( .INP(n606), .ZN(n607) );
  AND2X4 U474 ( .IN1(b[5]), .IN2(a[10]), .Q(n608) );
  XOR2X1 U475 ( .IN1(n699), .IN2(n294), .Q(n271) );
  XOR3X1 U476 ( .IN1(n404), .IN2(n426), .IN3(n514), .Q(n277) );
  NAND2X1 U477 ( .IN1(n514), .IN2(n404), .QN(n609) );
  NAND2X0 U478 ( .IN1(n426), .IN2(n404), .QN(n610) );
  NAND2X0 U479 ( .IN1(n426), .IN2(n514), .QN(n611) );
  NAND3X0 U480 ( .IN1(n609), .IN2(n611), .IN3(n610), .QN(n276) );
  OR2X1 U481 ( .IN1(n756), .IN2(n284), .Q(n612) );
  XOR2X1 U482 ( .IN1(n811), .IN2(n268), .Q(n249) );
  XOR3X1 U483 ( .IN1(n503), .IN2(n481), .IN3(n415), .Q(n281) );
  NAND2X0 U484 ( .IN1(n415), .IN2(n503), .QN(n613) );
  NAND2X0 U485 ( .IN1(n481), .IN2(n503), .QN(n614) );
  NAND2X0 U486 ( .IN1(n481), .IN2(n415), .QN(n615) );
  NAND3X0 U487 ( .IN1(n613), .IN2(n615), .IN3(n614), .QN(n280) );
  XOR3X1 U488 ( .IN1(n324), .IN2(n309), .IN3(n307), .Q(n305) );
  NAND2X0 U489 ( .IN1(n307), .IN2(n324), .QN(n616) );
  NAND2X0 U490 ( .IN1(n309), .IN2(n324), .QN(n617) );
  NAND2X1 U491 ( .IN1(n309), .IN2(n307), .QN(n618) );
  NAND3X0 U492 ( .IN1(n616), .IN2(n618), .IN3(n617), .QN(n304) );
  XOR2X1 U493 ( .IN1(n639), .IN2(n326), .Q(n307) );
  AND2X1 U494 ( .IN1(n285), .IN2(n304), .Q(n743) );
  XOR3X1 U495 ( .IN1(n330), .IN2(n315), .IN3(n313), .Q(n309) );
  NAND2X0 U496 ( .IN1(n330), .IN2(n315), .QN(n619) );
  NAND2X0 U497 ( .IN1(n330), .IN2(n313), .QN(n620) );
  NAND2X0 U498 ( .IN1(n315), .IN2(n313), .QN(n621) );
  NAND3X0 U499 ( .IN1(n619), .IN2(n620), .IN3(n621), .QN(n308) );
  XOR2X2 U500 ( .IN1(n291), .IN2(n293), .Q(n622) );
  XOR2X2 U501 ( .IN1(n622), .IN2(n308), .Q(n287) );
  NAND2X0 U502 ( .IN1(n291), .IN2(n293), .QN(n623) );
  NAND2X0 U503 ( .IN1(n291), .IN2(n308), .QN(n624) );
  NAND2X0 U504 ( .IN1(n293), .IN2(n308), .QN(n625) );
  NAND3X0 U505 ( .IN1(n623), .IN2(n624), .IN3(n625), .QN(n286) );
  XOR2X2 U506 ( .IN1(n781), .IN2(n666), .Q(n753) );
  NAND3X1 U507 ( .IN1(n826), .IN2(n825), .IN3(n824), .QN(n232) );
  OR2X4 U508 ( .IN1(n672), .IN2(n738), .Q(n454) );
  OAI21X1 U509 ( .IN1(n89), .IN2(n117), .IN3(n664), .QN(n835) );
  INVX0 U510 ( .INP(b[9]), .ZN(n626) );
  XOR3X1 U511 ( .IN1(n491), .IN2(n502), .IN3(n425), .Q(n259) );
  NAND2X1 U512 ( .IN1(n425), .IN2(n491), .QN(n627) );
  NAND2X1 U513 ( .IN1(n502), .IN2(n491), .QN(n628) );
  NAND2X1 U514 ( .IN1(n502), .IN2(n425), .QN(n629) );
  NAND3X0 U515 ( .IN1(n627), .IN2(n629), .IN3(n628), .QN(n258) );
  AND2X4 U516 ( .IN1(a[5]), .IN2(b[3]), .Q(n474) );
  NAND3X1 U517 ( .IN1(n812), .IN2(n814), .IN3(n813), .QN(n668) );
  AOI21X2 U518 ( .IN1(n118), .IN2(n126), .IN3(n119), .QN(n117) );
  XNOR3X1 U519 ( .IN1(n630), .IN2(n251), .IN3(n249), .Q(n247) );
  AND3X1 U520 ( .IN1(n784), .IN2(n783), .IN3(n782), .Q(n630) );
  HADDX2 U521 ( .A0(n452), .B0(n463), .C1(n350), .SO(n351) );
  OAI21X1 U522 ( .IN1(n631), .IN2(n632), .IN3(n633), .QN(n839) );
  OA21X1 U523 ( .IN1(n89), .IN2(n117), .IN3(n664), .Q(n631) );
  NAND2X0 U524 ( .IN1(n75), .IN2(n63), .QN(n632) );
  AOI21X1 U525 ( .IN1(n76), .IN2(n714), .IN3(n64), .QN(n633) );
  INVX0 U526 ( .INP(n286), .ZN(n634) );
  INVX0 U527 ( .INP(n634), .ZN(n635) );
  XOR3X1 U528 ( .IN1(n335), .IN2(n333), .IN3(n331), .Q(n327) );
  NAND2X0 U529 ( .IN1(n335), .IN2(n333), .QN(n636) );
  NAND2X0 U530 ( .IN1(n335), .IN2(n331), .QN(n637) );
  NAND2X0 U531 ( .IN1(n333), .IN2(n331), .QN(n638) );
  NAND3X0 U532 ( .IN1(n636), .IN2(n637), .IN3(n638), .QN(n326) );
  XOR2X2 U533 ( .IN1(n311), .IN2(n328), .Q(n639) );
  NAND2X0 U534 ( .IN1(n311), .IN2(n328), .QN(n640) );
  NAND2X0 U535 ( .IN1(n311), .IN2(n326), .QN(n641) );
  NAND2X0 U536 ( .IN1(n328), .IN2(n326), .QN(n642) );
  NAND3X0 U537 ( .IN1(n640), .IN2(n641), .IN3(n642), .QN(n306) );
  XOR2X1 U538 ( .IN1(n429), .IN2(n495), .Q(n643) );
  XOR2X2 U539 ( .IN1(n643), .IN2(n337), .Q(n331) );
  NAND2X0 U540 ( .IN1(n495), .IN2(n337), .QN(n644) );
  NAND2X0 U541 ( .IN1(n429), .IN2(n337), .QN(n645) );
  NAND2X0 U542 ( .IN1(n429), .IN2(n495), .QN(n646) );
  NAND3X0 U543 ( .IN1(n644), .IN2(n646), .IN3(n645), .QN(n330) );
  NAND3X2 U544 ( .IN1(n784), .IN2(n783), .IN3(n782), .QN(n661) );
  XNOR3X1 U545 ( .IN1(n647), .IN2(n235), .IN3(n233), .Q(n231) );
  AND3X1 U546 ( .IN1(n812), .IN2(n813), .IN3(n814), .Q(n647) );
  XOR2X1 U547 ( .IN1(n289), .IN2(n306), .Q(n648) );
  XOR2X2 U548 ( .IN1(n648), .IN2(n287), .Q(n285) );
  NAND2X0 U549 ( .IN1(n306), .IN2(n287), .QN(n649) );
  NAND2X0 U550 ( .IN1(n289), .IN2(n287), .QN(n650) );
  NAND2X0 U551 ( .IN1(n289), .IN2(n306), .QN(n651) );
  NAND3X0 U552 ( .IN1(n649), .IN2(n651), .IN3(n650), .QN(n284) );
  XOR3X2 U553 ( .IN1(n312), .IN2(n295), .IN3(n310), .Q(n289) );
  XOR3X1 U554 ( .IN1(n496), .IN2(n529), .IN3(n441), .Q(n349) );
  NAND2X0 U555 ( .IN1(n496), .IN2(n529), .QN(n652) );
  NAND2X0 U556 ( .IN1(n496), .IN2(n441), .QN(n653) );
  NAND2X1 U557 ( .IN1(n529), .IN2(n441), .QN(n654) );
  NAND3X0 U558 ( .IN1(n652), .IN2(n653), .IN3(n654), .QN(n348) );
  XOR2X1 U559 ( .IN1(n350), .IN2(n346), .Q(n655) );
  XOR2X2 U560 ( .IN1(n655), .IN2(n348), .Q(n329) );
  NAND2X0 U561 ( .IN1(n350), .IN2(n346), .QN(n656) );
  NAND2X0 U562 ( .IN1(n350), .IN2(n348), .QN(n657) );
  NAND2X0 U563 ( .IN1(n346), .IN2(n348), .QN(n658) );
  NAND3X0 U564 ( .IN1(n656), .IN2(n657), .IN3(n658), .QN(n328) );
  OR2X1 U565 ( .IN1(n725), .IN2(n537), .Q(n526) );
  FADDX1 U566 ( .A(n505), .B(n516), .CI(n428), .CO(n314), .S(n315) );
  XOR3X1 U567 ( .IN1(n282), .IN2(n403), .IN3(n280), .Q(n257) );
  NAND3X0 U568 ( .IN1(n687), .IN2(n688), .IN3(n689), .QN(n262) );
  NAND3X0 U569 ( .IN1(n761), .IN2(n762), .IN3(n763), .QN(n358) );
  INVX0 U570 ( .INP(a[6]), .ZN(n659) );
  OAI21X1 U571 ( .IN1(n89), .IN2(n117), .IN3(n664), .QN(n660) );
  XOR2X2 U572 ( .IN1(n839), .IN2(n662), .Q(product[19]) );
  AND2X4 U573 ( .IN1(n54), .IN2(n53), .Q(n662) );
  INVX0 U574 ( .INP(a[5]), .ZN(n663) );
  AOI21X1 U575 ( .IN1(n91), .IN2(n104), .IN3(n92), .QN(n664) );
  INVX0 U576 ( .INP(a[10]), .ZN(n665) );
  NAND3X0 U577 ( .IN1(n780), .IN2(n779), .IN3(n778), .QN(n666) );
  AND2X4 U578 ( .IN1(a[4]), .IN2(b[7]), .Q(n482) );
  INVX0 U579 ( .INP(a[5]), .ZN(n667) );
  INVX0 U580 ( .INP(a[9]), .ZN(n669) );
  INVX0 U581 ( .INP(a[9]), .ZN(n670) );
  INVX0 U582 ( .INP(a[9]), .ZN(n551) );
  INVX0 U583 ( .INP(b[11]), .ZN(n671) );
  INVX0 U584 ( .INP(a[6]), .ZN(n672) );
  XOR3X1 U585 ( .IN1(n242), .IN2(n229), .IN3(n227), .Q(n223) );
  NAND2X0 U586 ( .IN1(n227), .IN2(n242), .QN(n673) );
  NAND2X0 U587 ( .IN1(n229), .IN2(n242), .QN(n674) );
  NAND2X0 U588 ( .IN1(n229), .IN2(n227), .QN(n675) );
  NAND3X0 U589 ( .IN1(n673), .IN2(n675), .IN3(n674), .QN(n222) );
  XOR3X1 U590 ( .IN1(n207), .IN2(n220), .IN3(n218), .Q(n205) );
  NAND2X0 U591 ( .IN1(n218), .IN2(n207), .QN(n676) );
  NAND2X0 U592 ( .IN1(n220), .IN2(n207), .QN(n677) );
  NAND2X1 U593 ( .IN1(n220), .IN2(n218), .QN(n678) );
  NAND3X0 U594 ( .IN1(n676), .IN2(n678), .IN3(n677), .QN(n204) );
  XOR2X1 U595 ( .IN1(n222), .IN2(n211), .Q(n789) );
  AOI21X1 U596 ( .IN1(n116), .IN2(n103), .IN3(n104), .QN(n102) );
  XOR3X1 U597 ( .IN1(n345), .IN2(n347), .IN3(n356), .Q(n341) );
  XOR2X2 U598 ( .IN1(n354), .IN2(n343), .Q(n679) );
  XOR2X2 U599 ( .IN1(n679), .IN2(n341), .Q(n339) );
  NAND2X1 U600 ( .IN1(n345), .IN2(n347), .QN(n680) );
  NAND2X0 U601 ( .IN1(n345), .IN2(n356), .QN(n681) );
  NAND2X0 U602 ( .IN1(n347), .IN2(n356), .QN(n682) );
  NAND3X0 U603 ( .IN1(n680), .IN2(n681), .IN3(n682), .QN(n340) );
  NAND2X0 U604 ( .IN1(n354), .IN2(n343), .QN(n683) );
  NAND2X0 U605 ( .IN1(n354), .IN2(n341), .QN(n684) );
  NAND2X0 U606 ( .IN1(n343), .IN2(n341), .QN(n685) );
  NAND3X0 U607 ( .IN1(n683), .IN2(n684), .IN3(n685), .QN(n338) );
  NAND2X0 U608 ( .IN1(n336), .IN2(n321), .QN(n788) );
  XOR2X2 U609 ( .IN1(n336), .IN2(n321), .Q(n785) );
  INVX0 U610 ( .INP(a[8]), .ZN(n686) );
  XOR3X1 U611 ( .IN1(n436), .IN2(n458), .IN3(n414), .Q(n263) );
  NAND2X0 U612 ( .IN1(n436), .IN2(n458), .QN(n687) );
  NAND2X0 U613 ( .IN1(n436), .IN2(n414), .QN(n688) );
  NAND2X1 U614 ( .IN1(n458), .IN2(n414), .QN(n689) );
  XOR2X1 U615 ( .IN1(n260), .IN2(n245), .Q(n690) );
  XOR2X2 U616 ( .IN1(n690), .IN2(n262), .Q(n239) );
  NAND2X0 U617 ( .IN1(n260), .IN2(n245), .QN(n691) );
  NAND2X0 U618 ( .IN1(n260), .IN2(n262), .QN(n692) );
  NAND2X0 U619 ( .IN1(n245), .IN2(n262), .QN(n693) );
  NAND3X0 U620 ( .IN1(n691), .IN2(n692), .IN3(n693), .QN(n238) );
  OR2X1 U621 ( .IN1(n339), .IN2(n352), .Q(n837) );
  XOR3X1 U622 ( .IN1(n527), .IN2(n494), .IN3(n461), .Q(n317) );
  NAND2X1 U623 ( .IN1(n494), .IN2(n527), .QN(n694) );
  NAND2X0 U624 ( .IN1(n461), .IN2(n527), .QN(n695) );
  NAND2X0 U625 ( .IN1(n461), .IN2(n494), .QN(n696) );
  NAND3X0 U626 ( .IN1(n694), .IN2(n696), .IN3(n695), .QN(n316) );
  AOI21X1 U627 ( .IN1(n837), .IN2(n135), .IN3(n758), .QN(n697) );
  OA21X1 U628 ( .IN1(n127), .IN2(n139), .IN3(n697), .Q(n698) );
  AND2X4 U629 ( .IN1(b[10]), .IN2(a[4]), .Q(n479) );
  XOR2X2 U630 ( .IN1(n785), .IN2(n334), .Q(n313) );
  FADDX1 U631 ( .A(n372), .B(n363), .CI(n370), .CO(n356), .S(n357) );
  XOR2X2 U632 ( .IN1(n102), .IN2(n13), .Q(product[13]) );
  XNOR2X2 U633 ( .IN1(n703), .IN2(n14), .Q(product[12]) );
  NAND3X0 U634 ( .IN1(n824), .IN2(n825), .IN3(n826), .QN(n775) );
  FADDX1 U635 ( .A(n471), .B(n460), .CI(n416), .CO(n300), .S(n301) );
  XOR2X1 U636 ( .IN1(n281), .IN2(n277), .Q(n699) );
  NAND2X0 U637 ( .IN1(n277), .IN2(n294), .QN(n700) );
  NAND2X0 U638 ( .IN1(n281), .IN2(n294), .QN(n701) );
  NAND2X0 U639 ( .IN1(n281), .IN2(n277), .QN(n702) );
  NAND3X0 U640 ( .IN1(n700), .IN2(n702), .IN3(n701), .QN(n270) );
  AO21X1 U641 ( .IN1(n116), .IN2(n169), .IN3(n743), .Q(n703) );
  OR2X1 U642 ( .IN1(n748), .IN2(n671), .Q(n478) );
  XOR2X1 U643 ( .IN1(n478), .IN2(n401), .Q(n704) );
  XOR2X1 U644 ( .IN1(n704), .IN2(n244), .Q(n225) );
  NAND2X0 U645 ( .IN1(n401), .IN2(n244), .QN(n705) );
  NAND2X0 U646 ( .IN1(n478), .IN2(n244), .QN(n706) );
  NAND2X1 U647 ( .IN1(n478), .IN2(n401), .QN(n707) );
  NAND3X0 U648 ( .IN1(n705), .IN2(n707), .IN3(n706), .QN(n224) );
  INVX0 U649 ( .INP(b[5]), .ZN(n708) );
  NAND2X0 U650 ( .IN1(n251), .IN2(n661), .QN(n819) );
  AO21X1 U651 ( .IN1(n30), .IN2(n660), .IN3(n31), .Q(n841) );
  XOR3X1 U652 ( .IN1(n332), .IN2(n317), .IN3(n319), .Q(n311) );
  XOR2X2 U653 ( .IN1(n823), .IN2(n250), .Q(n233) );
  XOR3X1 U654 ( .IN1(n507), .IN2(n351), .IN3(n362), .Q(n345) );
  XOR3X1 U655 ( .IN1(n234), .IN2(n219), .IN3(n232), .Q(n217) );
  AND2X4 U656 ( .IN1(a[4]), .IN2(b[4]), .Q(n485) );
  AND2X4 U657 ( .IN1(a[6]), .IN2(b[9]), .Q(n456) );
  NOR2X0 U658 ( .IN1(n194), .IN2(n187), .QN(n709) );
  NOR2X0 U659 ( .IN1(n194), .IN2(n187), .QN(n710) );
  INVX0 U660 ( .INP(n163), .ZN(n711) );
  INVX0 U661 ( .INP(b[1]), .ZN(n712) );
  INVX0 U662 ( .INP(b[1]), .ZN(n547) );
  INVX0 U663 ( .INP(a[7]), .ZN(n713) );
  OR2X1 U664 ( .IN1(n667), .IN2(n671), .Q(n466) );
  OR2X1 U665 ( .IN1(n735), .IN2(n537), .Q(n514) );
  OR2X1 U666 ( .IN1(n720), .IN2(n537), .Q(n490) );
  AND2X4 U667 ( .IN1(a[0]), .IN2(b[6]), .Q(n531) );
  NOR2X0 U668 ( .IN1(n70), .IN2(n710), .QN(n714) );
  INVX0 U669 ( .INP(n78), .ZN(n715) );
  INVX0 U670 ( .INP(b[9]), .ZN(n716) );
  INVX0 U671 ( .INP(n36), .ZN(n717) );
  NOR2X0 U672 ( .IN1(n52), .IN2(n718), .QN(n34) );
  NAND2X0 U673 ( .IN1(n840), .IN2(n717), .QN(n718) );
  INVX0 U674 ( .INP(b[5]), .ZN(n719) );
  INVX0 U675 ( .INP(a[3]), .ZN(n720) );
  NOR2X0 U676 ( .IN1(n205), .IN2(n216), .QN(n721) );
  INVX0 U677 ( .INP(b[7]), .ZN(n722) );
  INVX0 U678 ( .INP(b[6]), .ZN(n723) );
  INVX0 U679 ( .INP(a[0]), .ZN(n724) );
  INVX0 U680 ( .INP(a[0]), .ZN(n725) );
  INVX0 U681 ( .INP(b[6]), .ZN(n726) );
  INVX0 U682 ( .INP(b[7]), .ZN(n541) );
  INVX0 U683 ( .INP(n743), .ZN(n727) );
  INVX0 U684 ( .INP(b[0]), .ZN(n728) );
  INVX0 U685 ( .INP(b[0]), .ZN(n548) );
  INVX0 U686 ( .INP(b[3]), .ZN(n729) );
  INVX0 U687 ( .INP(b[3]), .ZN(n545) );
  INVX0 U688 ( .INP(b[2]), .ZN(n730) );
  INVX0 U689 ( .INP(b[2]), .ZN(n546) );
  AND2X4 U690 ( .IN1(a[5]), .IN2(b[10]), .Q(n467) );
  INVX0 U691 ( .INP(a[11]), .ZN(n731) );
  INVX0 U692 ( .INP(a[11]), .ZN(n732) );
  INVX0 U693 ( .INP(a[11]), .ZN(n549) );
  INVX0 U694 ( .INP(b[8]), .ZN(n733) );
  INVX0 U695 ( .INP(b[8]), .ZN(n734) );
  INVX0 U696 ( .INP(a[1]), .ZN(n735) );
  INVX0 U697 ( .INP(a[1]), .ZN(n736) );
  INVX0 U698 ( .INP(a[1]), .ZN(n559) );
  INVX0 U699 ( .INP(b[5]), .ZN(n737) );
  INVX0 U700 ( .INP(b[11]), .ZN(n738) );
  INVX0 U701 ( .INP(b[11]), .ZN(n537) );
  INVX0 U702 ( .INP(b[9]), .ZN(n739) );
  INVX0 U703 ( .INP(a[8]), .ZN(n740) );
  INVX0 U704 ( .INP(a[8]), .ZN(n741) );
  INVX0 U705 ( .INP(a[8]), .ZN(n552) );
  AND2X4 U706 ( .IN1(a[4]), .IN2(b[6]), .Q(n483) );
  INVX0 U707 ( .INP(b[6]), .ZN(n742) );
  INVX0 U708 ( .INP(b[10]), .ZN(n744) );
  INVX0 U709 ( .INP(b[10]), .ZN(n538) );
  AND2X4 U710 ( .IN1(a[0]), .IN2(b[8]), .Q(n529) );
  INVX0 U711 ( .INP(a[2]), .ZN(n745) );
  OR2X1 U712 ( .IN1(n549), .IN2(n728), .Q(n405) );
  INVX0 U713 ( .INP(n117), .ZN(n746) );
  XNOR2X2 U714 ( .IN1(n746), .IN2(n15), .Q(product[11]) );
  AND2X4 U715 ( .IN1(a[1]), .IN2(b[9]), .Q(n516) );
  NAND2X0 U716 ( .IN1(b[1]), .IN2(a[11]), .QN(n404) );
  NAND2X0 U717 ( .IN1(n235), .IN2(n233), .QN(n833) );
  INVX0 U718 ( .INP(a[10]), .ZN(n747) );
  INVX0 U719 ( .INP(a[4]), .ZN(n748) );
  INVX0 U720 ( .INP(a[4]), .ZN(n749) );
  INVX0 U721 ( .INP(a[6]), .ZN(n750) );
  XNOR3X1 U722 ( .IN1(n286), .IN2(n269), .IN3(n751), .Q(n265) );
  XNOR2X1 U723 ( .IN1(n781), .IN2(n666), .Q(n751) );
  NOR2X0 U724 ( .IN1(n246), .IN2(n231), .QN(n752) );
  AND2X4 U725 ( .IN1(a[2]), .IN2(b[4]), .Q(n509) );
  INVX0 U726 ( .INP(a[7]), .ZN(n754) );
  INVX0 U727 ( .INP(a[7]), .ZN(n755) );
  INVX0 U728 ( .INP(a[7]), .ZN(n553) );
  AND2X4 U729 ( .IN1(a[8]), .IN2(b[4]), .Q(n437) );
  XOR3X1 U730 ( .IN1(n753), .IN2(n269), .IN3(n635), .Q(n756) );
  HADDX2 U731 ( .A0(n438), .B0(n449), .C1(n302), .SO(n303) );
  AND2X4 U732 ( .IN1(a[6]), .IN2(b[7]), .Q(n458) );
  INVX0 U733 ( .INP(a[0]), .ZN(n757) );
  AND2X4 U734 ( .IN1(n339), .IN2(n352), .Q(n758) );
  INVX0 U735 ( .INP(b[4]), .ZN(n759) );
  INVX0 U736 ( .INP(a[10]), .ZN(n760) );
  AND2X4 U737 ( .IN1(a[4]), .IN2(b[5]), .Q(n484) );
  AND2X1 U738 ( .IN1(a[3]), .IN2(b[5]), .Q(n496) );
  XOR2X2 U739 ( .IN1(n770), .IN2(n771), .Q(product[20]) );
  XOR3X1 U740 ( .IN1(n464), .IN2(n508), .IN3(n486), .Q(n359) );
  NAND2X0 U741 ( .IN1(n464), .IN2(n508), .QN(n761) );
  NAND2X0 U742 ( .IN1(n464), .IN2(n486), .QN(n762) );
  NAND2X1 U743 ( .IN1(n508), .IN2(n486), .QN(n763) );
  XOR2X1 U744 ( .IN1(n360), .IN2(n349), .Q(n764) );
  XOR2X2 U745 ( .IN1(n764), .IN2(n358), .Q(n343) );
  NAND2X0 U746 ( .IN1(n360), .IN2(n349), .QN(n765) );
  NAND2X0 U747 ( .IN1(n360), .IN2(n358), .QN(n766) );
  NAND2X0 U748 ( .IN1(n349), .IN2(n358), .QN(n767) );
  NAND3X0 U749 ( .IN1(n765), .IN2(n766), .IN3(n767), .QN(n342) );
  INVX0 U750 ( .INP(a[3]), .ZN(n557) );
  AND2X4 U751 ( .IN1(a[3]), .IN2(b[9]), .Q(n492) );
  XOR2X2 U752 ( .IN1(n834), .IN2(n768), .Q(product[21]) );
  AND2X4 U753 ( .IN1(n717), .IN2(n37), .Q(n768) );
  NOR2X0 U754 ( .IN1(n756), .IN2(n284), .QN(n769) );
  AND2X4 U755 ( .IN1(a[4]), .IN2(b[8]), .Q(n481) );
  AO21X1 U756 ( .IN1(n1), .IN2(n50), .IN3(n51), .Q(n770) );
  AND2X4 U757 ( .IN1(n840), .IN2(n48), .Q(n771) );
  XOR3X1 U758 ( .IN1(n275), .IN2(n290), .IN3(n607), .Q(n269) );
  NAND2X0 U759 ( .IN1(n290), .IN2(n292), .QN(n772) );
  NAND2X0 U760 ( .IN1(n275), .IN2(n292), .QN(n773) );
  NAND2X0 U761 ( .IN1(n275), .IN2(n290), .QN(n774) );
  NAND3X0 U762 ( .IN1(n772), .IN2(n774), .IN3(n773), .QN(n268) );
  FADDX1 U763 ( .A(n318), .B(n316), .CI(n299), .CO(n292), .S(n293) );
  AND2X4 U764 ( .IN1(a[3]), .IN2(b[4]), .Q(n497) );
  AND2X4 U765 ( .IN1(a[3]), .IN2(b[7]), .Q(n494) );
  OR2X4 U766 ( .IN1(n741), .IN2(n738), .Q(n430) );
  XNOR2X2 U767 ( .IN1(n1), .IN2(n11), .Q(product[15]) );
  INVX0 U768 ( .INP(b[8]), .ZN(n776) );
  FADDX1 U769 ( .A(n417), .B(n472), .CI(n439), .CO(n318), .S(n319) );
  INVX0 U770 ( .INP(a[2]), .ZN(n777) );
  XOR2X2 U771 ( .IN1(n95), .IN2(n12), .Q(product[14]) );
  INVX0 U772 ( .INP(a[2]), .ZN(n558) );
  NAND2X0 U773 ( .IN1(n312), .IN2(n295), .QN(n778) );
  NAND2X0 U774 ( .IN1(n312), .IN2(n310), .QN(n779) );
  NAND2X0 U775 ( .IN1(n295), .IN2(n310), .QN(n780) );
  NAND3X0 U776 ( .IN1(n780), .IN2(n779), .IN3(n778), .QN(n288) );
  XOR2X2 U777 ( .IN1(n271), .IN2(n273), .Q(n781) );
  NAND2X0 U778 ( .IN1(n271), .IN2(n273), .QN(n782) );
  NAND2X0 U779 ( .IN1(n271), .IN2(n288), .QN(n783) );
  NAND2X0 U780 ( .IN1(n273), .IN2(n288), .QN(n784) );
  NAND2X0 U781 ( .IN1(n321), .IN2(n334), .QN(n786) );
  NAND2X0 U782 ( .IN1(n336), .IN2(n334), .QN(n787) );
  NAND3X0 U783 ( .IN1(n786), .IN2(n788), .IN3(n787), .QN(n312) );
  XOR3X1 U784 ( .IN1(n213), .IN2(n215), .IN3(n224), .Q(n209) );
  XOR2X2 U785 ( .IN1(n789), .IN2(n209), .Q(n207) );
  NAND2X0 U786 ( .IN1(n213), .IN2(n215), .QN(n790) );
  NAND2X0 U787 ( .IN1(n213), .IN2(n224), .QN(n791) );
  NAND2X0 U788 ( .IN1(n215), .IN2(n224), .QN(n792) );
  NAND3X0 U789 ( .IN1(n790), .IN2(n791), .IN3(n792), .QN(n208) );
  NAND2X0 U790 ( .IN1(n222), .IN2(n211), .QN(n793) );
  NAND2X0 U791 ( .IN1(n222), .IN2(n209), .QN(n794) );
  NAND2X0 U792 ( .IN1(n211), .IN2(n209), .QN(n795) );
  NAND3X0 U793 ( .IN1(n793), .IN2(n794), .IN3(n795), .QN(n206) );
  NAND2X0 U794 ( .IN1(n286), .IN2(n753), .QN(n796) );
  NAND2X0 U795 ( .IN1(n269), .IN2(n753), .QN(n797) );
  NAND2X0 U796 ( .IN1(n269), .IN2(n286), .QN(n798) );
  NAND3X0 U797 ( .IN1(n796), .IN2(n798), .IN3(n797), .QN(n264) );
  XOR3X1 U798 ( .IN1(n440), .IN2(n473), .IN3(n506), .Q(n333) );
  NAND2X0 U799 ( .IN1(n506), .IN2(n440), .QN(n799) );
  NAND2X0 U800 ( .IN1(n473), .IN2(n440), .QN(n800) );
  NAND2X1 U801 ( .IN1(n473), .IN2(n506), .QN(n801) );
  NAND3X0 U802 ( .IN1(n799), .IN2(n801), .IN3(n800), .QN(n332) );
  XOR3X1 U803 ( .IN1(n236), .IN2(n223), .IN3(n221), .Q(n219) );
  NAND2X1 U804 ( .IN1(n236), .IN2(n223), .QN(n802) );
  NAND2X0 U805 ( .IN1(n236), .IN2(n221), .QN(n803) );
  NAND2X0 U806 ( .IN1(n223), .IN2(n221), .QN(n804) );
  NAND3X0 U807 ( .IN1(n804), .IN2(n803), .IN3(n802), .QN(n218) );
  NAND2X0 U808 ( .IN1(n775), .IN2(n234), .QN(n805) );
  NAND2X0 U809 ( .IN1(n775), .IN2(n219), .QN(n806) );
  NAND2X0 U810 ( .IN1(n234), .IN2(n219), .QN(n807) );
  NAND3X0 U811 ( .IN1(n805), .IN2(n806), .IN3(n807), .QN(n216) );
  XOR3X1 U812 ( .IN1(n225), .IN2(n240), .IN3(n238), .Q(n221) );
  NAND2X0 U813 ( .IN1(n238), .IN2(n225), .QN(n808) );
  NAND2X0 U814 ( .IN1(n240), .IN2(n225), .QN(n809) );
  NAND2X1 U815 ( .IN1(n240), .IN2(n238), .QN(n810) );
  NAND3X0 U816 ( .IN1(n808), .IN2(n810), .IN3(n809), .QN(n220) );
  XOR2X1 U817 ( .IN1(n270), .IN2(n253), .Q(n811) );
  NAND2X0 U818 ( .IN1(n253), .IN2(n268), .QN(n812) );
  NAND2X0 U819 ( .IN1(n270), .IN2(n268), .QN(n813) );
  NAND2X0 U820 ( .IN1(n270), .IN2(n253), .QN(n814) );
  INVX0 U821 ( .INP(n167), .ZN(n815) );
  INVX0 U822 ( .INP(a[5]), .ZN(n816) );
  INVX0 U823 ( .INP(a[5]), .ZN(n555) );
  NAND2X0 U824 ( .IN1(n661), .IN2(n249), .QN(n817) );
  NAND2X0 U825 ( .IN1(n251), .IN2(n249), .QN(n818) );
  NAND3X0 U826 ( .IN1(n817), .IN2(n818), .IN3(n819), .QN(n246) );
  OAI21X2 U827 ( .IN1(n815), .IN2(n106), .IN3(n101), .QN(n97) );
  XOR3X1 U828 ( .IN1(n272), .IN2(n274), .IN3(n255), .Q(n251) );
  NAND2X0 U829 ( .IN1(n272), .IN2(n274), .QN(n820) );
  NAND2X0 U830 ( .IN1(n272), .IN2(n255), .QN(n821) );
  NAND2X0 U831 ( .IN1(n274), .IN2(n255), .QN(n822) );
  NAND3X0 U832 ( .IN1(n822), .IN2(n821), .IN3(n820), .QN(n250) );
  XOR2X2 U833 ( .IN1(n252), .IN2(n237), .Q(n823) );
  NAND2X0 U834 ( .IN1(n252), .IN2(n237), .QN(n824) );
  NAND2X0 U835 ( .IN1(n252), .IN2(n250), .QN(n825) );
  NAND2X0 U836 ( .IN1(n237), .IN2(n250), .QN(n826) );
  XOR3X1 U837 ( .IN1(n279), .IN2(n283), .IN3(n296), .Q(n273) );
  NAND2X0 U838 ( .IN1(n296), .IN2(n279), .QN(n827) );
  NAND2X0 U839 ( .IN1(n283), .IN2(n279), .QN(n828) );
  NAND2X0 U840 ( .IN1(n283), .IN2(n296), .QN(n829) );
  NAND3X0 U841 ( .IN1(n827), .IN2(n829), .IN3(n828), .QN(n272) );
  OR2X1 U842 ( .IN1(n216), .IN2(n205), .Q(n830) );
  NAND2X0 U843 ( .IN1(n233), .IN2(n668), .QN(n831) );
  NAND2X0 U844 ( .IN1(n235), .IN2(n668), .QN(n832) );
  NAND3X0 U845 ( .IN1(n831), .IN2(n833), .IN3(n832), .QN(n230) );
  AO21X1 U846 ( .IN1(n39), .IN2(n1), .IN3(n40), .Q(n834) );
  NAND2X0 U847 ( .IN1(n167), .IN2(n101), .QN(n13) );
  NAND2X0 U848 ( .IN1(n169), .IN2(n727), .QN(n15) );
  NAND2X0 U849 ( .IN1(n837), .IN2(n132), .QN(n18) );
  NAND2X0 U850 ( .IN1(n162), .IN2(n66), .QN(n8) );
  NAND2X0 U851 ( .IN1(n170), .IN2(n121), .QN(n16) );
  NAND2X0 U852 ( .IN1(n171), .IN2(n124), .QN(n17) );
  XOR2X2 U853 ( .IN1(n841), .IN2(n842), .Q(product[22]) );
  NOR2X0 U854 ( .IN1(n180), .IN2(n177), .QN(n836) );
  FADDX1 U855 ( .A(n183), .B(n190), .CI(n188), .CO(n180), .S(n181) );
  INVX0 U856 ( .INP(n103), .ZN(n105) );
  INVX0 U857 ( .INP(n98), .ZN(n167) );
  NAND2X0 U858 ( .IN1(n166), .IN2(n94), .QN(n12) );
  INVX0 U859 ( .INP(n752), .ZN(n166) );
  INVX0 U860 ( .INP(n104), .ZN(n106) );
  INVX0 U861 ( .INP(n86), .ZN(n84) );
  NOR2X0 U862 ( .IN1(n247), .IN2(n264), .QN(n98) );
  INVX0 U863 ( .INP(n75), .ZN(n77) );
  NAND2X0 U864 ( .IN1(n163), .IN2(n73), .QN(n9) );
  INVX0 U865 ( .INP(n70), .ZN(n163) );
  INVX0 U866 ( .INP(n114), .ZN(n169) );
  NAND2X0 U867 ( .IN1(n264), .IN2(n247), .QN(n101) );
  NAND2X0 U868 ( .IN1(n82), .IN2(n830), .QN(n10) );
  INVX0 U869 ( .INP(n709), .ZN(n162) );
  NAND2X0 U870 ( .IN1(n612), .IN2(n110), .QN(n14) );
  INVX0 U871 ( .INP(n120), .ZN(n170) );
  INVX0 U872 ( .INP(n123), .ZN(n171) );
  INVX0 U873 ( .INP(n137), .ZN(n135) );
  INVX0 U874 ( .INP(n76), .ZN(n78) );
  NOR2X0 U875 ( .IN1(n204), .IN2(n195), .QN(n70) );
  NAND2X0 U876 ( .IN1(n323), .IN2(n338), .QN(n124) );
  INVX0 U877 ( .INP(n34), .ZN(n32) );
  NAND2X0 U878 ( .IN1(n304), .IN2(n285), .QN(n115) );
  NAND2X0 U879 ( .IN1(n194), .IN2(n187), .QN(n66) );
  NOR2X0 U880 ( .IN1(n323), .IN2(n338), .QN(n123) );
  NOR2X0 U881 ( .IN1(n305), .IN2(n322), .QN(n120) );
  NAND2X0 U882 ( .IN1(n322), .IN2(n305), .QN(n121) );
  NOR2X0 U883 ( .IN1(n194), .IN2(n187), .QN(n65) );
  NAND2X0 U884 ( .IN1(n339), .IN2(n352), .QN(n132) );
  OR2X1 U885 ( .IN1(n353), .IN2(n364), .Q(n838) );
  NAND2X0 U886 ( .IN1(n353), .IN2(n364), .QN(n137) );
  NAND2X0 U887 ( .IN1(n265), .IN2(n284), .QN(n110) );
  INVX0 U888 ( .INP(n52), .ZN(n54) );
  NAND2X0 U889 ( .IN1(n365), .IN2(n374), .QN(n143) );
  OA21X1 U890 ( .IN1(n53), .IN2(n836), .IN3(n48), .Q(n44) );
  INVX0 U891 ( .INP(n139), .ZN(n138) );
  INVX0 U892 ( .INP(n35), .ZN(n33) );
  OR2X1 U893 ( .IN1(n180), .IN2(n177), .Q(n840) );
  NAND2X0 U894 ( .IN1(n180), .IN2(n177), .QN(n48) );
  NOR2X0 U895 ( .IN1(n375), .IN2(n382), .QN(n144) );
  NOR2X0 U896 ( .IN1(n383), .IN2(n388), .QN(n147) );
  AND2X1 U897 ( .IN1(n846), .IN2(n28), .Q(n842) );
  OA21X1 U898 ( .IN1(n843), .IN2(n844), .IN3(n845), .Q(n139) );
  OR2X1 U899 ( .IN1(n142), .IN2(n144), .Q(n843) );
  OA21X1 U900 ( .IN1(n147), .IN2(n149), .IN3(n148), .Q(n844) );
  OA21X1 U901 ( .IN1(n145), .IN2(n142), .IN3(n143), .Q(n845) );
  NAND2X0 U902 ( .IN1(n34), .IN2(n846), .QN(n23) );
  INVX0 U903 ( .INP(n28), .ZN(n26) );
  NAND2X0 U904 ( .IN1(n375), .IN2(n382), .QN(n145) );
  NAND2X0 U905 ( .IN1(n383), .IN2(n388), .QN(n148) );
  NOR2X0 U906 ( .IN1(n176), .IN2(n175), .QN(n36) );
  OR2X1 U907 ( .IN1(n174), .IN2(n394), .Q(n846) );
  NOR2X0 U908 ( .IN1(n393), .IN2(n513), .QN(n155) );
  NAND2X0 U909 ( .IN1(n174), .IN2(n394), .QN(n28) );
  NAND2X0 U910 ( .IN1(n393), .IN2(n513), .QN(n156) );
  NAND2X0 U911 ( .IN1(n176), .IN2(n175), .QN(n37) );
  NOR2X0 U912 ( .IN1(n389), .IN2(n392), .QN(n152) );
  NAND2X0 U913 ( .IN1(n389), .IN2(n392), .QN(n153) );
  OA21X1 U914 ( .IN1(n152), .IN2(n847), .IN3(n153), .Q(n149) );
  OA21X1 U915 ( .IN1(n157), .IN2(n155), .IN3(n156), .Q(n847) );
  OR2X1 U916 ( .IN1(n745), .IN2(n738), .Q(n502) );
  INVX0 U917 ( .INP(b[4]), .ZN(n544) );
  OR2X1 U918 ( .IN1(n713), .IN2(n671), .Q(n442) );
  OR2X1 U919 ( .IN1(n669), .IN2(n671), .Q(n418) );
  OR2X1 U920 ( .IN1(n747), .IN2(n671), .Q(n406) );
  NOR2X0 U921 ( .IN1(n731), .IN2(n738), .QN(n394) );
  NAND2X0 U922 ( .IN1(n536), .IN2(n525), .QN(n157) );
  NOR2X0 U923 ( .IN1(n285), .IN2(n304), .QN(n114) );
  NOR2X0 U924 ( .IN1(n720), .IN2(n728), .QN(n501) );
  NAND2X0 U925 ( .IN1(n84), .IN2(n87), .QN(n11) );
  INVX0 U926 ( .INP(n87), .ZN(n85) );
  INVX0 U927 ( .INP(n117), .ZN(n116) );
  NOR2X0 U928 ( .IN1(n365), .IN2(n374), .QN(n142) );
  NAND2X0 U929 ( .IN1(n246), .IN2(n231), .QN(n94) );
  NAND2X0 U930 ( .IN1(n838), .IN2(n137), .QN(n19) );
  NAND2X0 U931 ( .IN1(n837), .IN2(n838), .QN(n127) );
  NOR2X0 U932 ( .IN1(n720), .IN2(n744), .QN(n491) );
  NAND2X0 U933 ( .IN1(n54), .IN2(n840), .QN(n41) );
  NOR2X0 U934 ( .IN1(n557), .IN2(n726), .QN(n495) );
  NOR2X0 U935 ( .IN1(n720), .IN2(n733), .QN(n493) );
  NAND2X0 U936 ( .IN1(n230), .IN2(n217), .QN(n87) );
  NOR2X0 U937 ( .IN1(n77), .IN2(n711), .QN(n68) );
  NAND2X0 U938 ( .IN1(n75), .IN2(n714), .QN(n3) );
  NOR2X0 U939 ( .IN1(n557), .IN2(n712), .QN(n500) );
  NOR2X0 U940 ( .IN1(n720), .IN2(n729), .QN(n498) );
  NOR2X0 U941 ( .IN1(n120), .IN2(n123), .QN(n118) );
  NOR2X0 U942 ( .IN1(n713), .IN2(n541), .QN(n446) );
  NOR2X0 U943 ( .IN1(n754), .IN2(n742), .QN(n447) );
  NOR2X0 U944 ( .IN1(n754), .IN2(n544), .QN(n449) );
  NOR2X0 U945 ( .IN1(n626), .IN2(n553), .QN(n444) );
  NOR2X0 U946 ( .IN1(n755), .IN2(n737), .QN(n448) );
  NOR2X0 U947 ( .IN1(n553), .IN2(n776), .QN(n445) );
  NOR2X0 U948 ( .IN1(n755), .IN2(n548), .QN(n453) );
  NOR2X0 U949 ( .IN1(n755), .IN2(n545), .QN(n450) );
  NOR2X0 U950 ( .IN1(n553), .IN2(n547), .QN(n452) );
  NOR2X0 U951 ( .IN1(n713), .IN2(n744), .QN(n443) );
  NOR2X0 U952 ( .IN1(n754), .IN2(n546), .QN(n451) );
  NOR2X0 U953 ( .IN1(n769), .IN2(n114), .QN(n103) );
  NOR2X0 U954 ( .IN1(n284), .IN2(n265), .QN(n109) );
  NOR2X0 U955 ( .IN1(n757), .IN2(n712), .QN(n536) );
  NOR2X0 U956 ( .IN1(n757), .IN2(n730), .QN(n535) );
  NOR2X0 U957 ( .IN1(n725), .IN2(n729), .QN(n534) );
  NOR2X0 U958 ( .IN1(n757), .IN2(n708), .QN(n532) );
  NOR2X0 U959 ( .IN1(n724), .IN2(n759), .QN(n533) );
  NOR2X0 U960 ( .IN1(n757), .IN2(n541), .QN(n530) );
  NOR2X0 U961 ( .IN1(n724), .IN2(n716), .QN(n528) );
  NOR2X0 U962 ( .IN1(n744), .IN2(n725), .QN(n527) );
  NOR2X0 U963 ( .IN1(n672), .IN2(n733), .QN(n457) );
  NOR2X0 U964 ( .IN1(n659), .IN2(n723), .QN(n459) );
  NOR2X0 U965 ( .IN1(n672), .IN2(n538), .QN(n455) );
  NOR2X0 U966 ( .IN1(n659), .IN2(n548), .QN(n465) );
  NOR2X0 U967 ( .IN1(n659), .IN2(n546), .QN(n463) );
  NOR2X0 U968 ( .IN1(n750), .IN2(n737), .QN(n460) );
  NOR2X0 U969 ( .IN1(n659), .IN2(n545), .QN(n462) );
  NOR2X0 U970 ( .IN1(n659), .IN2(n544), .QN(n461) );
  NOR2X0 U971 ( .IN1(n659), .IN2(n547), .QN(n464) );
  NOR2X0 U972 ( .IN1(n557), .IN2(n730), .QN(n499) );
  NOR2X0 U973 ( .IN1(n105), .IN2(n815), .QN(n96) );
  NOR2X0 U974 ( .IN1(n752), .IN2(n98), .QN(n91) );
  NOR2X0 U975 ( .IN1(n559), .IN2(n728), .QN(n525) );
  NOR2X0 U976 ( .IN1(n735), .IN2(n712), .QN(n524) );
  NOR2X0 U977 ( .IN1(n559), .IN2(n730), .QN(n523) );
  NOR2X0 U978 ( .IN1(n735), .IN2(n729), .QN(n522) );
  NOR2X0 U979 ( .IN1(n735), .IN2(n708), .QN(n520) );
  NOR2X0 U980 ( .IN1(n559), .IN2(n759), .QN(n521) );
  NOR2X0 U981 ( .IN1(n736), .IN2(n722), .QN(n518) );
  NOR2X0 U982 ( .IN1(n736), .IN2(n538), .QN(n515) );
  NOR2X0 U983 ( .IN1(n559), .IN2(n726), .QN(n519) );
  NOR2X0 U984 ( .IN1(n736), .IN2(n734), .QN(n517) );
  NOR2X0 U985 ( .IN1(n3), .IN2(n23), .QN(n21) );
  NOR2X0 U986 ( .IN1(n3), .IN2(n32), .QN(n30) );
  NOR2X0 U987 ( .IN1(n3), .IN2(n52), .QN(n50) );
  NOR2X0 U988 ( .IN1(n3), .IN2(n41), .QN(n39) );
  NAND2X0 U989 ( .IN1(n204), .IN2(n195), .QN(n73) );
  NOR2X0 U990 ( .IN1(n749), .IN2(n728), .QN(n489) );
  NOR2X0 U991 ( .IN1(n748), .IN2(n712), .QN(n488) );
  NOR2X0 U992 ( .IN1(n749), .IN2(n546), .QN(n487) );
  NOR2X0 U993 ( .IN1(n749), .IN2(n729), .QN(n486) );
  NOR2X0 U994 ( .IN1(n748), .IN2(n716), .QN(n480) );
  NOR2X0 U995 ( .IN1(n558), .IN2(n728), .QN(n513) );
  NOR2X0 U996 ( .IN1(n745), .IN2(n712), .QN(n512) );
  NOR2X0 U997 ( .IN1(n558), .IN2(n730), .QN(n511) );
  NOR2X0 U998 ( .IN1(n558), .IN2(n723), .QN(n507) );
  NOR2X0 U999 ( .IN1(n777), .IN2(n776), .QN(n505) );
  NOR2X0 U1000 ( .IN1(n558), .IN2(n626), .QN(n504) );
  NOR2X0 U1001 ( .IN1(n777), .IN2(n744), .QN(n503) );
  NOR2X0 U1002 ( .IN1(n558), .IN2(n545), .QN(n510) );
  NOR2X0 U1003 ( .IN1(n745), .IN2(n541), .QN(n506) );
  NOR2X0 U1004 ( .IN1(n745), .IN2(n719), .QN(n508) );
  NAND2X0 U1005 ( .IN1(n91), .IN2(n103), .QN(n89) );
  NOR2X0 U1006 ( .IN1(n552), .IN2(n538), .QN(n431) );
  NOR2X0 U1007 ( .IN1(n686), .IN2(n541), .QN(n434) );
  NOR2X0 U1008 ( .IN1(n741), .IN2(n734), .QN(n433) );
  NOR2X0 U1009 ( .IN1(n552), .IN2(n739), .QN(n432) );
  NOR2X0 U1010 ( .IN1(n686), .IN2(n742), .QN(n435) );
  NOR2X0 U1011 ( .IN1(n740), .IN2(n708), .QN(n436) );
  NOR2X0 U1012 ( .IN1(n740), .IN2(n548), .QN(n441) );
  NOR2X0 U1013 ( .IN1(n686), .IN2(n545), .QN(n438) );
  NOR2X0 U1014 ( .IN1(n552), .IN2(n547), .QN(n440) );
  NOR2X0 U1015 ( .IN1(n741), .IN2(n730), .QN(n439) );
  NAND2X0 U1016 ( .IN1(n181), .IN2(n186), .QN(n53) );
  NOR2X0 U1017 ( .IN1(n186), .IN2(n181), .QN(n52) );
  NOR2X0 U1018 ( .IN1(n555), .IN2(n739), .QN(n468) );
  NOR2X0 U1019 ( .IN1(n816), .IN2(n728), .QN(n477) );
  NOR2X0 U1020 ( .IN1(n555), .IN2(n733), .QN(n469) );
  NOR2X0 U1021 ( .IN1(n667), .IN2(n722), .QN(n470) );
  NOR2X0 U1022 ( .IN1(n667), .IN2(n730), .QN(n475) );
  NOR2X0 U1023 ( .IN1(n555), .IN2(n547), .QN(n476) );
  NOR2X0 U1024 ( .IN1(n667), .IN2(n759), .QN(n473) );
  NOR2X0 U1025 ( .IN1(n816), .IN2(n726), .QN(n471) );
  NOR2X0 U1026 ( .IN1(n663), .IN2(n719), .QN(n472) );
  NOR2X0 U1027 ( .IN1(n86), .IN2(n721), .QN(n75) );
  NOR2X0 U1028 ( .IN1(n217), .IN2(n230), .QN(n86) );
  NOR2X0 U1029 ( .IN1(n70), .IN2(n709), .QN(n63) );
  NAND2X0 U1030 ( .IN1(n205), .IN2(n216), .QN(n82) );
  NOR2X0 U1031 ( .IN1(n205), .IN2(n216), .QN(n81) );
  NOR2X0 U1032 ( .IN1(n670), .IN2(n739), .QN(n420) );
  NOR2X0 U1033 ( .IN1(n551), .IN2(n548), .QN(n429) );
  NOR2X0 U1034 ( .IN1(n670), .IN2(n538), .QN(n419) );
  NOR2X0 U1035 ( .IN1(n669), .IN2(n734), .QN(n421) );
  NOR2X0 U1036 ( .IN1(n669), .IN2(n726), .QN(n423) );
  NOR2X0 U1037 ( .IN1(n670), .IN2(n737), .QN(n424) );
  NOR2X0 U1038 ( .IN1(n670), .IN2(n722), .QN(n422) );
  NOR2X0 U1039 ( .IN1(n670), .IN2(n759), .QN(n425) );
  NOR2X0 U1040 ( .IN1(n669), .IN2(n729), .QN(n426) );
  NOR2X0 U1041 ( .IN1(n551), .IN2(n547), .QN(n428) );
  NOR2X0 U1042 ( .IN1(n551), .IN2(n730), .QN(n427) );
  NOR2X0 U1043 ( .IN1(n231), .IN2(n246), .QN(n93) );
  NOR2X0 U1044 ( .IN1(n747), .IN2(n744), .QN(n407) );
  NOR2X0 U1045 ( .IN1(n665), .IN2(n716), .QN(n408) );
  NOR2X0 U1046 ( .IN1(n747), .IN2(n733), .QN(n409) );
  NOR2X0 U1047 ( .IN1(n747), .IN2(n722), .QN(n410) );
  NOR2X0 U1048 ( .IN1(n747), .IN2(n723), .QN(n411) );
  NOR2X0 U1049 ( .IN1(n747), .IN2(n544), .QN(n413) );
  NOR2X0 U1050 ( .IN1(n665), .IN2(n545), .QN(n414) );
  NOR2X0 U1051 ( .IN1(n665), .IN2(n546), .QN(n415) );
  NOR2X0 U1052 ( .IN1(n665), .IN2(n547), .QN(n416) );
  NOR2X0 U1053 ( .IN1(n760), .IN2(n548), .QN(n417) );
  OAI21X2 U1054 ( .IN1(n117), .IN2(n89), .IN3(n90), .QN(n1) );
endmodule


module multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0 ( in_a, in_b, \output  );
  input [11:0] in_a;
  input [11:0] in_b;
  output [11:0] \output ;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;
  wire   [23:7] pre_out;
  wire   [11:0] rnd_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7;

  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0_DW01_inc_2 add_37_round ( .A(
        pre_out[19:7]), .SUM({rnd_out, SYNOPSYS_UNCONNECTED__0}) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0_DW_mult_tc_3 mult_35 ( .a(in_a), 
        .b(in_b), .product({pre_out, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7}) );
  AND2X1 U2 ( .IN1(n17), .IN2(n16), .Q(n3) );
  AND2X1 U3 ( .IN1(n17), .IN2(n16), .Q(n6) );
  AO21X1 U4 ( .IN1(rnd_out[0]), .IN2(n1), .IN3(n6), .Q(\output [0]) );
  DELLN2X2 U5 ( .INP(n10), .Z(n1) );
  INVX0 U6 ( .INP(n4), .ZN(n2) );
  AND2X1 U7 ( .IN1(n17), .IN2(n16), .Q(n12) );
  INVX0 U8 ( .INP(n19), .ZN(n4) );
  INVX0 U9 ( .INP(n4), .ZN(n5) );
  NOR2X0 U10 ( .IN1(pre_out[20]), .IN2(pre_out[21]), .QN(n7) );
  NOR2X0 U11 ( .IN1(pre_out[22]), .IN2(pre_out[19]), .QN(n8) );
  NAND2X0 U12 ( .IN1(n18), .IN2(n11), .QN(n9) );
  NAND2X0 U13 ( .IN1(n18), .IN2(n11), .QN(n10) );
  NAND3X0 U14 ( .IN1(n7), .IN2(n8), .IN3(n16), .QN(n11) );
  AND2X1 U15 ( .IN1(pre_out[21]), .IN2(pre_out[23]), .Q(n13) );
  NAND2X0 U16 ( .IN1(n11), .IN2(n18), .QN(n19) );
  AO21X1 U17 ( .IN1(rnd_out[4]), .IN2(n19), .IN3(n6), .Q(\output [4]) );
  AO21X1 U18 ( .IN1(rnd_out[1]), .IN2(n10), .IN3(n3), .Q(\output [1]) );
  AO21X1 U19 ( .IN1(rnd_out[9]), .IN2(n19), .IN3(n3), .Q(\output [9]) );
  AO21X1 U20 ( .IN1(rnd_out[5]), .IN2(n9), .IN3(n12), .Q(\output [5]) );
  MUX21X1 U21 ( .IN1(pre_out[23]), .IN2(rnd_out[11]), .S(n5), .Q(\output [11])
         );
  INVX0 U22 ( .INP(pre_out[23]), .ZN(n16) );
  AO21X1 U23 ( .IN1(n2), .IN2(rnd_out[10]), .IN3(n3), .Q(\output [10]) );
  AO21X1 U24 ( .IN1(rnd_out[8]), .IN2(n9), .IN3(n6), .Q(\output [8]) );
  AO21X1 U25 ( .IN1(rnd_out[2]), .IN2(n20), .IN3(n6), .Q(\output [2]) );
  AO21X1 U26 ( .IN1(rnd_out[3]), .IN2(n20), .IN3(n12), .Q(\output [3]) );
  AO21X1 U27 ( .IN1(rnd_out[7]), .IN2(n19), .IN3(n3), .Q(\output [7]) );
  NOR2X0 U28 ( .IN1(pre_out[20]), .IN2(pre_out[21]), .QN(n15) );
  NAND2X0 U29 ( .IN1(n11), .IN2(n18), .QN(n20) );
  NOR2X0 U30 ( .IN1(pre_out[22]), .IN2(pre_out[19]), .QN(n14) );
  NAND4X0 U31 ( .IN1(n13), .IN2(pre_out[22]), .IN3(pre_out[19]), .IN4(
        pre_out[20]), .QN(n18) );
  NAND3X0 U32 ( .IN1(n15), .IN2(n14), .IN3(n16), .QN(n17) );
  AO21X1 U33 ( .IN1(rnd_out[6]), .IN2(n10), .IN3(n6), .Q(\output [6]) );
endmodule



    module inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_DW01_sub_4 ( 
        A, B, CI, DIFF, CO );
  input [11:0] A;
  input [11:0] B;
  output [11:0] DIFF;
  input CI;
  output CO;
  wire   n6, n7, n8, n9, n10, n11, n22, n23, n24, n25, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n38, n39, n40, n43, n44, n45, n46, n47, n51, n52,
         n53, n55, n56, n57, n59, n60, n61, n62, n63, n65, n66, n68, n69, n70,
         n71, n73, n74, n75, n76, n77, n79, n80, n81, n82, n84, n88, n90, n92,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174;

  OAI21X1 U17 ( .IN1(n30), .IN2(n24), .IN3(n25), .QN(n23) );
  AOI21X1 U33 ( .IN1(n46), .IN2(n33), .IN3(n34), .QN(n32) );
  OAI21X1 U35 ( .IN1(n43), .IN2(n35), .IN3(n36), .QN(n34) );
  OAI21X1 U57 ( .IN1(n57), .IN2(n51), .IN3(n52), .QN(n46) );
  XNOR2X1 U62 ( .IN1(n171), .IN2(n8), .Q(DIFF[4]) );
  AOI21X1 U63 ( .IN1(n171), .IN2(n139), .IN3(n55), .QN(n53) );
  AOI21X1 U72 ( .IN1(n68), .IN2(n151), .IN3(n61), .QN(n59) );
  OAI21X1 U74 ( .IN1(n66), .IN2(n62), .IN3(n63), .QN(n61) );
  XOR2X2 U108 ( .IN1(n92), .IN2(n135), .Q(DIFF[0]) );
  INVX32 U109 ( .INP(A[0]), .ZN(n135) );
  XOR2X2 U110 ( .IN1(n11), .IN2(n71), .Q(DIFF[1]) );
  XOR2X1 U111 ( .IN1(n136), .IN2(n10), .Q(DIFF[2]) );
  OA21X1 U112 ( .IN1(n71), .IN2(n69), .IN3(n70), .Q(n136) );
  XOR2X2 U113 ( .IN1(n53), .IN2(n7), .Q(DIFF[5]) );
  XOR2X2 U114 ( .IN1(n44), .IN2(n6), .Q(DIFF[6]) );
  XOR2X2 U115 ( .IN1(n137), .IN2(n138), .Q(DIFF[7]) );
  AO21X1 U116 ( .IN1(n171), .IN2(n38), .IN3(n39), .Q(n137) );
  AND2X4 U117 ( .IN1(n75), .IN2(n36), .Q(n138) );
  OR2X1 U118 ( .IN1(B[4]), .IN2(n149), .Q(n57) );
  OR2X1 U119 ( .IN1(n88), .IN2(A[4]), .Q(n139) );
  XOR2X2 U120 ( .IN1(n144), .IN2(n140), .Q(DIFF[8]) );
  AND2X4 U121 ( .IN1(n74), .IN2(n30), .Q(n140) );
  OA21X1 U122 ( .IN1(n57), .IN2(n51), .IN3(n52), .Q(n141) );
  AOI21X1 U123 ( .IN1(n171), .IN2(n45), .IN3(n46), .QN(n44) );
  OAI21X2 U124 ( .IN1(n168), .IN2(n31), .IN3(n32), .QN(n144) );
  OAI21X1 U125 ( .IN1(n71), .IN2(n69), .IN3(n70), .QN(n68) );
  INVX0 U126 ( .INP(A[0]), .ZN(n165) );
  INVX0 U127 ( .INP(A[1]), .ZN(n163) );
  INVX0 U128 ( .INP(A[5]), .ZN(n164) );
  INVX0 U129 ( .INP(A[6]), .ZN(n153) );
  AO21X1 U130 ( .IN1(n68), .IN2(n151), .IN3(n160), .Q(n171) );
  XOR2X2 U131 ( .IN1(n142), .IN2(n9), .Q(DIFF[3]) );
  OA21X1 U132 ( .IN1(n136), .IN2(n150), .IN3(n152), .Q(n142) );
  AND2X1 U133 ( .IN1(n82), .IN2(A[10]), .Q(n143) );
  OR2X1 U134 ( .IN1(B[9]), .IN2(n162), .Q(n25) );
  INVX0 U135 ( .INP(B[2]), .ZN(n145) );
  INVX0 U136 ( .INP(A[7]), .ZN(n146) );
  OR2X1 U137 ( .IN1(B[7]), .IN2(n146), .Q(n36) );
  OAI21X1 U138 ( .IN1(n152), .IN2(n62), .IN3(n63), .QN(n160) );
  XOR2X1 U139 ( .IN1(n147), .IN2(n148), .Q(DIFF[9]) );
  AND2X4 U140 ( .IN1(n73), .IN2(n25), .Q(n147) );
  AO21X1 U141 ( .IN1(n167), .IN2(n74), .IN3(n28), .Q(n148) );
  INVX0 U142 ( .INP(A[9]), .ZN(n162) );
  INVX0 U143 ( .INP(A[4]), .ZN(n149) );
  AND2X1 U144 ( .IN1(B[3]), .IN2(n173), .Q(n62) );
  INVX0 U145 ( .INP(A[3]), .ZN(n173) );
  OR2X1 U146 ( .IN1(B[3]), .IN2(n173), .Q(n63) );
  INVX0 U147 ( .INP(n80), .ZN(n150) );
  NOR2X0 U148 ( .IN1(n65), .IN2(n62), .QN(n151) );
  OR2X1 U149 ( .IN1(B[6]), .IN2(n153), .Q(n43) );
  NAND2X0 U150 ( .IN1(A[2]), .IN2(n145), .QN(n152) );
  AND2X1 U151 ( .IN1(B[6]), .IN2(n153), .Q(n40) );
  XOR2X2 U152 ( .IN1(n154), .IN2(A[11]), .Q(DIFF[11]) );
  OA21X1 U153 ( .IN1(n157), .IN2(n156), .IN3(n158), .Q(n154) );
  XOR2X2 U154 ( .IN1(n169), .IN2(n170), .Q(DIFF[10]) );
  INVX0 U155 ( .INP(B[2]), .ZN(n155) );
  OA21X1 U156 ( .IN1(n31), .IN2(n59), .IN3(n32), .Q(n156) );
  NAND2X0 U157 ( .IN1(n22), .IN2(n174), .QN(n157) );
  AOI21X1 U158 ( .IN1(n23), .IN2(n174), .IN3(n143), .QN(n158) );
  INVX0 U159 ( .INP(n143), .ZN(n159) );
  NAND2X0 U160 ( .IN1(A[4]), .IN2(n88), .QN(n161) );
  OR2X1 U161 ( .IN1(B[1]), .IN2(n163), .Q(n70) );
  AND2X1 U162 ( .IN1(B[9]), .IN2(n162), .Q(n24) );
  OR2X1 U163 ( .IN1(B[5]), .IN2(n164), .Q(n52) );
  AND2X1 U164 ( .IN1(B[1]), .IN2(n163), .Q(n69) );
  AND2X1 U165 ( .IN1(B[5]), .IN2(n164), .Q(n51) );
  AND2X1 U166 ( .IN1(B[0]), .IN2(n165), .Q(n71) );
  AOI21X1 U167 ( .IN1(n68), .IN2(n60), .IN3(n61), .QN(n166) );
  OAI21X1 U168 ( .IN1(n31), .IN2(n166), .IN3(n32), .QN(n167) );
  AOI21X1 U169 ( .IN1(n68), .IN2(n60), .IN3(n160), .QN(n168) );
  AO21X1 U170 ( .IN1(n172), .IN2(n22), .IN3(n23), .Q(n169) );
  AND2X4 U171 ( .IN1(n174), .IN2(n159), .Q(n170) );
  AND2X1 U172 ( .IN1(B[7]), .IN2(n146), .Q(n35) );
  OAI21X1 U173 ( .IN1(n31), .IN2(n168), .IN3(n32), .QN(n172) );
  INVX0 U174 ( .INP(B[0]), .ZN(n92) );
  INVX0 U175 ( .INP(B[8]), .ZN(n84) );
  INVX0 U176 ( .INP(B[4]), .ZN(n88) );
  INVX0 U177 ( .INP(n40), .ZN(n76) );
  INVX0 U178 ( .INP(n51), .ZN(n77) );
  INVX0 U179 ( .INP(n62), .ZN(n79) );
  INVX0 U180 ( .INP(n65), .ZN(n80) );
  INVX0 U181 ( .INP(n69), .ZN(n81) );
  INVX0 U182 ( .INP(n161), .ZN(n55) );
  OAI21X1 U183 ( .IN1(n40), .IN2(n141), .IN3(n43), .QN(n39) );
  INVX0 U184 ( .INP(n45), .ZN(n47) );
  INVX0 U185 ( .INP(n35), .ZN(n75) );
  INVX0 U186 ( .INP(n29), .ZN(n74) );
  INVX0 U187 ( .INP(n24), .ZN(n73) );
  INVX0 U188 ( .INP(n30), .ZN(n28) );
  OR2X1 U189 ( .IN1(n82), .IN2(A[10]), .Q(n174) );
  NAND2X0 U190 ( .IN1(n66), .IN2(n80), .QN(n10) );
  NAND2X0 U191 ( .IN1(n139), .IN2(n161), .QN(n8) );
  NAND2X0 U192 ( .IN1(n79), .IN2(n63), .QN(n9) );
  NAND2X0 U193 ( .IN1(n70), .IN2(n81), .QN(n11) );
  NAND2X0 U194 ( .IN1(n77), .IN2(n52), .QN(n7) );
  NAND2X0 U195 ( .IN1(n76), .IN2(n43), .QN(n6) );
  NOR2X0 U196 ( .IN1(n84), .IN2(A[8]), .QN(n29) );
  NAND2X0 U197 ( .IN1(n84), .IN2(A[8]), .QN(n30) );
  NOR2X0 U198 ( .IN1(n65), .IN2(n62), .QN(n60) );
  INVX0 U199 ( .INP(B[2]), .ZN(n90) );
  NOR2X0 U200 ( .IN1(n56), .IN2(n51), .QN(n45) );
  NOR2X0 U201 ( .IN1(n88), .IN2(A[4]), .QN(n56) );
  INVX0 U202 ( .INP(B[10]), .ZN(n82) );
  NAND2X0 U203 ( .IN1(A[2]), .IN2(n155), .QN(n66) );
  NOR2X0 U204 ( .IN1(n90), .IN2(A[2]), .QN(n65) );
  NOR2X0 U205 ( .IN1(n47), .IN2(n40), .QN(n38) );
  NAND2X0 U206 ( .IN1(n45), .IN2(n33), .QN(n31) );
  NOR2X0 U207 ( .IN1(n40), .IN2(n35), .QN(n33) );
  NOR2X0 U208 ( .IN1(n29), .IN2(n24), .QN(n22) );
endmodule



    module inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16 ( 
        \input , \output , clk, rst, start, done );
  input [11:0] \input ;
  output [11:0] \output ;
  input clk, rst, start;
  output done;
  wire   state, out_reg_enable, N46, N47, N48, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, n82, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n132, n133, n134, n135, n136, n137, n138, N255, N254, N253, N252,
         N251, N250, N249, N248, N247, N246, N245, N244, N220, N228, n1, n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n131, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333;
  wire   [11:0] input_2;
  wire   [3:0] shift_amount;
  wire   [7:1] input_shifted;
  wire   [11:0] sel_poly;
  wire   [3:0] out_shift_amount;
  wire   [11:0] pre_output;
  wire   [11:0] mult1_out;
  wire   [11:0] mult2_out;
  wire   [11:1] mult3_out;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5;

  DFFARX1 state_reg ( .D(n138), .CLK(clk), .RSTB(n129), .Q(state), .QN(n130)
         );
  DFFARX1 \counter_reg[0]  ( .D(n130), .CLK(clk), .RSTB(n129), .QN(n93) );
  DFFARX1 \counter_reg[1]  ( .D(N46), .CLK(clk), .RSTB(n129), .QN(n94) );
  DFFARX1 \counter_reg[2]  ( .D(N47), .CLK(clk), .RSTB(n129), .QN(n95) );
  DFFARX1 \counter_reg[3]  ( .D(N48), .CLK(clk), .RSTB(n129), .QN(n96) );
  DFFARX1 out_reg_enable_reg ( .D(n137), .CLK(clk), .RSTB(n129), .Q(
        out_reg_enable), .QN(n152) );
  DFFARX1 done_reg ( .D(n136), .CLK(clk), .RSTB(n129), .Q(done) );
  DFFX1 \input_reg_reg[10]  ( .D(n127), .CLK(clk), .Q(input_2[10]), .QN(n103)
         );
  DFFX1 \input_reg_reg[3]  ( .D(n120), .CLK(clk), .Q(input_2[3]), .QN(n99) );
  DFFX1 \input_reg_reg[2]  ( .D(n119), .CLK(clk), .Q(input_2[2]), .QN(n98) );
  DFFX1 \output_reg_reg[11]  ( .D(n116), .CLK(clk), .Q(\output [11]), .QN(n17)
         );
  DFFX1 \output_reg_reg[10]  ( .D(n115), .CLK(clk), .Q(\output [10]) );
  DFFX1 \output_reg_reg[9]  ( .D(n114), .CLK(clk), .Q(\output [9]) );
  DFFX1 \output_reg_reg[8]  ( .D(n113), .CLK(clk), .Q(\output [8]) );
  DFFX1 \output_reg_reg[7]  ( .D(n112), .CLK(clk), .Q(\output [7]) );
  DFFX1 \output_reg_reg[6]  ( .D(n111), .CLK(clk), .Q(\output [6]) );
  DFFX1 \output_reg_reg[5]  ( .D(n110), .CLK(clk), .Q(\output [5]) );
  DFFX1 \output_reg_reg[4]  ( .D(n109), .CLK(clk), .Q(\output [4]) );
  DFFX1 \output_reg_reg[3]  ( .D(n108), .CLK(clk), .Q(\output [3]) );
  DFFX1 \output_reg_reg[2]  ( .D(n107), .CLK(clk), .Q(\output [2]) );
  DFFX1 \output_reg_reg[1]  ( .D(n106), .CLK(clk), .Q(\output [1]) );
  DFFX1 \output_reg_reg[0]  ( .D(n105), .CLK(clk), .Q(\output [0]) );
  AO22X1 U86 ( .IN1(n333), .IN2(done), .IN3(state), .IN4(n82), .Q(n136) );
  AO21X1 U88 ( .IN1(start), .IN2(n130), .IN3(n333), .Q(n138) );
  shifter_WORD_WIDTH12_LOG_WORD_WIDTH4_SMALLER_POW2_WW16_MAX_LEFT8_MAX_RIGHT3 in_shift ( 
        .\input ({input_2[11:3], n158, input_2[1], n159}), .\output ({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, input_shifted[7:6], 
        N220, input_shifted[4], N228, input_shifted[2:1], 
        SYNOPSYS_UNCONNECTED__4}), .direction(n11), .amount({n144, 
        shift_amount[2:1], n79}) );
  shifter_WORD_WIDTH12_LOG_WORD_WIDTH4_SMALLER_POW2_WW16_MAX_LEFT4_MAX_RIGHT2 out_shift ( 
        .\input ({1'b0, 1'b0, 1'b0, n332, sel_poly[7:0]}), .\output (
        pre_output), .direction(n11), .amount({1'b0, n144, 
        out_shift_amount[1:0]}) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_2 mult1 ( .in_a(pre_output), 
        .in_b(pre_output), .\output (mult1_out) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_1 mult2 ( .in_a({n6, 
        pre_output[10], n68, pre_output[8], n70, n8, pre_output[5], n67, 
        pre_output[3:0]}), .in_b({input_2[11:3], n88, input_2[1], n80}), 
        .\output (mult2_out) );
  multiplier_WORD_WIDTH12_INT_BITS4_USE_SAT1_0 mult3 ( .in_a(mult1_out), 
        .in_b(mult2_out), .\output ({mult3_out, SYNOPSYS_UNCONNECTED__5}) );
  inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16_DW01_sub_4 sub_0_root_sub_0_root_sub_287 ( 
        .A({N255, N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, 
        N244}), .B({1'b0, mult3_out}), .CI(1'b0), .DIFF({N267, N266, N265, 
        N264, N263, N262, N261, N260, N259, N258, N257, N256}) );
  DFFX2 \input_reg_reg[7]  ( .D(n124), .CLK(clk), .Q(input_2[7]), .QN(n100) );
  DFFX2 \input_reg_reg[1]  ( .D(n118), .CLK(clk), .Q(input_2[1]), .QN(n135) );
  DFFX1 \input_reg_reg[0]  ( .D(n117), .CLK(clk), .Q(input_2[0]), .QN(n97) );
  DFFX1 \input_reg_reg[6]  ( .D(n123), .CLK(clk), .Q(input_2[6]), .QN(n132) );
  DFFX2 \input_reg_reg[9]  ( .D(n126), .CLK(clk), .Q(input_2[9]), .QN(n102) );
  DFFX2 \input_reg_reg[5]  ( .D(n122), .CLK(clk), .Q(input_2[5]), .QN(n133) );
  DFFX1 \input_reg_reg[8]  ( .D(n125), .CLK(clk), .Q(input_2[8]), .QN(n101) );
  DFFX1 \input_reg_reg[4]  ( .D(n121), .CLK(clk), .Q(input_2[4]), .QN(n134) );
  DFFX1 \input_reg_reg[11]  ( .D(n128), .CLK(clk), .Q(input_2[11]), .QN(n104)
         );
  XNOR2X2 U3 ( .IN1(N228), .IN2(input_shifted[6]), .Q(n196) );
  AND2X2 U4 ( .IN1(input_shifted[6]), .IN2(n217), .Q(n71) );
  XOR2X2 U5 ( .IN1(pre_output[0]), .IN2(n45), .Q(N244) );
  INVX0 U6 ( .INP(shift_amount[1]), .ZN(n1) );
  INVX0 U7 ( .INP(n1), .ZN(n2) );
  DELLN1X2 U8 ( .INP(n57), .Z(n3) );
  INVX0 U9 ( .INP(input_2[10]), .ZN(n4) );
  OAI21X2 U10 ( .IN1(n92), .IN2(n176), .IN3(n175), .QN(n177) );
  DELLN2X2 U11 ( .INP(pre_output[10]), .Z(n5) );
  XOR2X1 U12 ( .IN1(n10), .IN2(n249), .Q(n252) );
  NBUFFX4 U13 ( .INP(pre_output[11]), .Z(n6) );
  AND2X4 U14 ( .IN1(n11), .IN2(n79), .Q(n7) );
  INVX0 U15 ( .INP(n265), .ZN(n8) );
  NAND2X0 U16 ( .IN1(n307), .IN2(n305), .QN(n274) );
  OR2X1 U17 ( .IN1(n145), .IN2(n259), .Q(n232) );
  INVX0 U18 ( .INP(pre_output[9]), .ZN(n9) );
  NOR2X0 U19 ( .IN1(n248), .IN2(n247), .QN(n10) );
  MUX21X1 U20 ( .IN1(n210), .IN2(n209), .S(n251), .Q(sel_poly[3]) );
  MUX21X1 U21 ( .IN1(n198), .IN2(n197), .S(n251), .Q(sel_poly[2]) );
  NOR2X0 U22 ( .IN1(n152), .IN2(n309), .QN(n150) );
  INVX0 U23 ( .INP(n250), .ZN(n251) );
  AOI21X1 U24 ( .IN1(n177), .IN2(n25), .IN3(n3), .QN(n11) );
  AND2X1 U25 ( .IN1(n89), .IN2(n85), .Q(n12) );
  AND2X4 U26 ( .IN1(n61), .IN2(n43), .Q(n13) );
  AND2X4 U27 ( .IN1(n153), .IN2(n163), .Q(n14) );
  AND2X1 U28 ( .IN1(n74), .IN2(n75), .Q(n15) );
  AND2X4 U29 ( .IN1(n327), .IN2(n150), .Q(n16) );
  DELLN2X2 U30 ( .INP(pre_output[4]), .Z(n18) );
  MUX21X1 U31 ( .IN1(n226), .IN2(n225), .S(n251), .Q(sel_poly[4]) );
  AND2X1 U32 ( .IN1(n52), .IN2(n246), .Q(n19) );
  INVX0 U33 ( .INP(n234), .ZN(n20) );
  INVX0 U34 ( .INP(n20), .ZN(n21) );
  INVX0 U35 ( .INP(pre_output[4]), .ZN(n22) );
  MUX21X2 U36 ( .IN1(n176), .IN2(\input [11]), .S(start), .Q(n128) );
  NAND2X0 U37 ( .IN1(n61), .IN2(n43), .QN(n23) );
  AND4X1 U38 ( .IN1(n55), .IN2(n164), .IN3(n165), .IN4(n133), .Q(n24) );
  XOR2X1 U39 ( .IN1(n63), .IN2(n237), .Q(n238) );
  AND2X2 U40 ( .IN1(n14), .IN2(n147), .Q(n144) );
  NAND2X0 U41 ( .IN1(n262), .IN2(n307), .QN(n273) );
  NAND2X0 U42 ( .IN1(n262), .IN2(n263), .QN(n278) );
  NAND3X0 U43 ( .IN1(n41), .IN2(n100), .IN3(n132), .QN(n166) );
  OAI221X1 U44 ( .IN1(n149), .IN2(n171), .IN3(n170), .IN4(n169), .IN5(n168), 
        .QN(n25) );
  AO22X1 U45 ( .IN1(n229), .IN2(n228), .IN3(n76), .IN4(n242), .Q(n239) );
  OR3X1 U46 ( .IN1(n40), .IN2(n84), .IN3(n131), .Q(n170) );
  INVX0 U47 ( .INP(N220), .ZN(n26) );
  XNOR2X1 U48 ( .IN1(n235), .IN2(n28), .Q(n259) );
  INVX0 U49 ( .INP(n26), .ZN(n27) );
  OR2X1 U50 ( .IN1(input_shifted[6]), .IN2(N228), .Q(n214) );
  INVX0 U51 ( .INP(input_shifted[4]), .ZN(n28) );
  INVX0 U52 ( .INP(n35), .ZN(n29) );
  INVX0 U53 ( .INP(n298), .ZN(n30) );
  OAI21X1 U54 ( .IN1(n59), .IN2(n215), .IN3(n218), .QN(n201) );
  XOR2X1 U55 ( .IN1(n28), .IN2(input_shifted[1]), .Q(n186) );
  INVX0 U56 ( .INP(n227), .ZN(n31) );
  INVX0 U57 ( .INP(input_shifted[7]), .ZN(n32) );
  DELLN2X2 U58 ( .INP(shift_amount[2]), .Z(n33) );
  AND2X1 U59 ( .IN1(n102), .IN2(n104), .Q(n83) );
  INVX0 U60 ( .INP(n266), .ZN(n34) );
  INVX0 U61 ( .INP(input_shifted[4]), .ZN(n35) );
  OR3X2 U62 ( .IN1(N228), .IN2(input_shifted[4]), .IN3(N220), .Q(n246) );
  NAND2X0 U63 ( .IN1(n143), .IN2(n231), .QN(n222) );
  NAND3X1 U64 ( .IN1(n51), .IN2(n52), .IN3(n246), .QN(n261) );
  XOR2X2 U65 ( .IN1(n213), .IN2(n43), .Q(n255) );
  NOR2X0 U66 ( .IN1(n23), .IN2(n32), .QN(n36) );
  INVX0 U67 ( .INP(n53), .ZN(n37) );
  INVX0 U68 ( .INP(n37), .ZN(n38) );
  MUX21X2 U69 ( .IN1(n287), .IN2(n286), .S(n285), .Q(N250) );
  AO21X1 U70 ( .IN1(n183), .IN2(n7), .IN3(n33), .Q(out_shift_amount[1]) );
  NAND2X0 U71 ( .IN1(n134), .IN2(n133), .QN(n39) );
  AND3X1 U72 ( .IN1(n132), .IN2(n101), .IN3(n99), .Q(n86) );
  AND2X1 U73 ( .IN1(n102), .IN2(n101), .Q(n149) );
  AND2X1 U74 ( .IN1(n100), .IN2(n102), .Q(n164) );
  AND4X1 U75 ( .IN1(n86), .IN2(n100), .IN3(n134), .IN4(n133), .Q(n163) );
  NAND4X0 U76 ( .IN1(n55), .IN2(n39), .IN3(n85), .IN4(n155), .QN(n168) );
  INVX0 U77 ( .INP(n100), .ZN(n40) );
  AND2X1 U78 ( .IN1(n134), .IN2(n133), .Q(n41) );
  MUX21X2 U79 ( .IN1(n297), .IN2(n296), .S(n295), .Q(N245) );
  INVX0 U80 ( .INP(N220), .ZN(n42) );
  INVX0 U81 ( .INP(n42), .ZN(n43) );
  INVX0 U82 ( .INP(pre_output[1]), .ZN(n44) );
  INVX0 U83 ( .INP(n44), .ZN(n45) );
  NAND2X0 U84 ( .IN1(n141), .IN2(n241), .QN(n46) );
  XOR2X2 U85 ( .IN1(n7), .IN2(n2), .Q(out_shift_amount[0]) );
  DELLN2X2 U87 ( .INP(pre_output[7]), .Z(n47) );
  INVX0 U89 ( .INP(n18), .ZN(n48) );
  INVX0 U90 ( .INP(input_shifted[6]), .ZN(n49) );
  INVX0 U91 ( .INP(input_shifted[7]), .ZN(n50) );
  INVX0 U92 ( .INP(n50), .ZN(n51) );
  INVX0 U93 ( .INP(n49), .ZN(n52) );
  NAND2X0 U94 ( .IN1(n203), .IN2(n202), .QN(n53) );
  INVX0 U95 ( .INP(n235), .ZN(n54) );
  AND2X1 U96 ( .IN1(n104), .IN2(n103), .Q(n55) );
  DELLN1X2 U97 ( .INP(input_2[9]), .Z(n56) );
  AO21X1 U98 ( .IN1(n60), .IN2(n166), .IN3(n148), .Q(n57) );
  MUX21X2 U99 ( .IN1(n56), .IN2(\input [9]), .S(start), .Q(n126) );
  INVX0 U100 ( .INP(input_shifted[1]), .ZN(n58) );
  AND2X1 U101 ( .IN1(n52), .IN2(n246), .Q(n146) );
  MUX21X2 U102 ( .IN1(input_2[6]), .IN2(\input [6]), .S(start), .Q(n123) );
  INVX0 U103 ( .INP(n79), .ZN(n250) );
  AND3X1 U104 ( .IN1(n139), .IN2(n184), .IN3(n180), .Q(n79) );
  OA221X1 U105 ( .IN1(n261), .IN2(n142), .IN3(n260), .IN4(n261), .IN5(n251), 
        .Q(n332) );
  INVX0 U106 ( .INP(N220), .ZN(n59) );
  AND2X1 U107 ( .IN1(n149), .IN2(n55), .Q(n60) );
  INVX0 U108 ( .INP(n49), .ZN(n61) );
  INVX0 U109 ( .INP(n61), .ZN(n62) );
  INVX0 U110 ( .INP(n245), .ZN(n63) );
  INVX0 U111 ( .INP(n305), .ZN(n64) );
  OAI221X1 U112 ( .IN1(n149), .IN2(n171), .IN3(n170), .IN4(n169), .IN5(n168), 
        .QN(n182) );
  NAND2X0 U113 ( .IN1(n298), .IN2(n48), .QN(n302) );
  NAND2X0 U114 ( .IN1(n48), .IN2(n300), .QN(n268) );
  DELLN2X2 U115 ( .INP(pre_output[8]), .Z(n65) );
  INVX0 U116 ( .INP(n300), .ZN(n66) );
  INVX0 U117 ( .INP(n22), .ZN(n67) );
  INVX0 U118 ( .INP(n9), .ZN(n68) );
  NAND2X0 U119 ( .IN1(n223), .IN2(n222), .QN(n258) );
  NAND2X0 U120 ( .IN1(n222), .IN2(n221), .QN(n207) );
  NAND2X0 U121 ( .IN1(n141), .IN2(n53), .QN(n69) );
  NBUFFX4 U122 ( .INP(pre_output[7]), .Z(n70) );
  MUX21X2 U123 ( .IN1(n162), .IN2(\input [4]), .S(start), .Q(n121) );
  AND2X1 U124 ( .IN1(n160), .IN2(n83), .Q(n154) );
  MUX21X1 U125 ( .IN1(n191), .IN2(n190), .S(n251), .Q(sel_poly[1]) );
  NAND2X0 U126 ( .IN1(n16), .IN2(N267), .QN(n328) );
  NAND3X0 U127 ( .IN1(n178), .IN2(n12), .IN3(n24), .QN(n179) );
  AND2X1 U128 ( .IN1(n218), .IN2(n227), .Q(n72) );
  AND3X1 U129 ( .IN1(n220), .IN2(n219), .IN3(n72), .Q(n145) );
  AND2X1 U130 ( .IN1(n218), .IN2(n205), .Q(n143) );
  INVX0 U131 ( .INP(n307), .ZN(n73) );
  MUX21X2 U132 ( .IN1(n156), .IN2(\input [3]), .S(start), .Q(n120) );
  NAND2X0 U133 ( .IN1(n15), .IN2(n328), .QN(n116) );
  OR2X4 U134 ( .IN1(n330), .IN2(n329), .Q(n75) );
  OR2X1 U135 ( .IN1(out_reg_enable), .IN2(n17), .Q(n74) );
  NAND2X0 U136 ( .IN1(out_reg_enable), .IN2(n309), .QN(n330) );
  NAND2X0 U137 ( .IN1(n64), .IN2(n327), .QN(n329) );
  MUX21X1 U138 ( .IN1(n238), .IN2(n239), .S(n250), .Q(sel_poly[5]) );
  NOR2X0 U139 ( .IN1(n69), .IN2(n211), .QN(n76) );
  NAND2X0 U140 ( .IN1(n201), .IN2(n221), .QN(n192) );
  NAND3X1 U141 ( .IN1(n200), .IN2(n201), .IN3(n221), .QN(n199) );
  INVX0 U142 ( .INP(n265), .ZN(n77) );
  MUX21X2 U143 ( .IN1(n158), .IN2(\input [2]), .S(start), .Q(n119) );
  INVX0 U144 ( .INP(n262), .ZN(n78) );
  MUX21X2 U145 ( .IN1(input_2[8]), .IN2(\input [8]), .S(start), .Q(n125) );
  INVX0 U146 ( .INP(n97), .ZN(n80) );
  AND3X1 U147 ( .IN1(n81), .IN2(n103), .IN3(n98), .Q(n147) );
  NAND2X0 U148 ( .IN1(n135), .IN2(n97), .QN(n81) );
  INVX0 U149 ( .INP(n132), .ZN(n84) );
  INVX0 U150 ( .INP(n84), .ZN(n85) );
  INVX0 U151 ( .INP(input_2[2]), .ZN(n87) );
  INVX0 U152 ( .INP(n87), .ZN(n88) );
  INVX0 U153 ( .INP(input_2[8]), .ZN(n89) );
  INVX0 U154 ( .INP(n100), .ZN(n90) );
  INVX0 U155 ( .INP(n131), .ZN(n91) );
  INVX0 U156 ( .INP(input_2[10]), .ZN(n92) );
  NAND2X0 U157 ( .IN1(n147), .IN2(n99), .QN(n169) );
  INVX0 U158 ( .INP(n104), .ZN(n131) );
  OA21X1 U159 ( .IN1(n92), .IN2(n176), .IN3(n175), .Q(n139) );
  OR2X1 U160 ( .IN1(n46), .IN2(n211), .Q(n229) );
  NAND2X0 U161 ( .IN1(n233), .IN2(n232), .QN(n140) );
  NAND2X0 U162 ( .IN1(n255), .IN2(n140), .QN(n237) );
  NAND2X0 U163 ( .IN1(n233), .IN2(n232), .QN(n256) );
  MUX21X2 U164 ( .IN1(input_2[1]), .IN2(\input [1]), .S(start), .Q(n118) );
  XOR2X2 U165 ( .IN1(n65), .IN2(n78), .Q(n281) );
  NAND2X0 U166 ( .IN1(n49), .IN2(n235), .QN(n221) );
  NAND2X0 U167 ( .IN1(n71), .IN2(n216), .QN(n219) );
  MUX21X2 U168 ( .IN1(n189), .IN2(n186), .S(n251), .Q(sel_poly[0]) );
  NAND2X0 U169 ( .IN1(n266), .IN2(n300), .QN(n267) );
  INVX0 U170 ( .INP(n283), .ZN(n304) );
  INVX0 U171 ( .INP(n289), .ZN(n269) );
  INVX0 U172 ( .INP(n228), .ZN(n242) );
  INVX0 U173 ( .INP(n211), .ZN(n240) );
  INVX0 U174 ( .INP(pre_output[3]), .ZN(n300) );
  INVX0 U175 ( .INP(pre_output[5]), .ZN(n298) );
  XOR2X1 U176 ( .IN1(n77), .IN2(n47), .Q(n287) );
  NAND2X0 U177 ( .IN1(n284), .IN2(n283), .QN(n286) );
  INVX0 U178 ( .INP(pre_output[2]), .ZN(n266) );
  NAND2X0 U179 ( .IN1(n289), .IN2(n302), .QN(n291) );
  INVX0 U180 ( .INP(n301), .ZN(n297) );
  NAND2X0 U181 ( .IN1(n244), .IN2(n243), .QN(n254) );
  INVX0 U182 ( .INP(n201), .ZN(n203) );
  INVX0 U183 ( .INP(n188), .ZN(n185) );
  AND2X1 U184 ( .IN1(n200), .IN2(n59), .Q(n141) );
  XNOR2X1 U185 ( .IN1(n189), .IN2(n193), .Q(n190) );
  INVX0 U186 ( .INP(n230), .ZN(n223) );
  AND2X1 U187 ( .IN1(n245), .IN2(n255), .Q(n142) );
  INVX0 U188 ( .INP(input_shifted[1]), .ZN(n217) );
  INVX0 U189 ( .INP(n261), .ZN(n247) );
  INVX0 U190 ( .INP(n196), .ZN(n187) );
  INVX0 U191 ( .INP(n308), .ZN(n272) );
  NAND3X1 U192 ( .IN1(n43), .IN2(n202), .IN3(n199), .QN(n204) );
  NAND3X0 U193 ( .IN1(n214), .IN2(n215), .IN3(n27), .QN(n220) );
  INVX0 U194 ( .INP(n25), .ZN(n183) );
  NAND2X0 U195 ( .IN1(n278), .IN2(n308), .QN(n280) );
  INVX0 U196 ( .INP(n330), .ZN(n325) );
  INVX0 U197 ( .INP(pre_output[11]), .ZN(n305) );
  INVX0 U198 ( .INP(n82), .ZN(n333) );
  AND4X1 U199 ( .IN1(n55), .IN2(n165), .IN3(n133), .IN4(n164), .Q(n148) );
  INVX0 U200 ( .INP(n134), .ZN(n162) );
  MUX21X1 U201 ( .IN1(input_2[7]), .IN2(\input [7]), .S(start), .Q(n124) );
  INVX0 U202 ( .INP(n99), .ZN(n156) );
  MUX21X1 U203 ( .IN1(n159), .IN2(\input [0]), .S(start), .Q(n117) );
  NOR2X0 U204 ( .IN1(input_2[5]), .IN2(input_2[6]), .QN(n310) );
  NOR2X0 U205 ( .IN1(n327), .IN2(n152), .QN(n151) );
  NOR2X0 U206 ( .IN1(input_2[11]), .IN2(input_2[10]), .QN(n312) );
  INVX0 U207 ( .INP(out_reg_enable), .ZN(n324) );
  NAND2X1 U208 ( .IN1(state), .IN2(n96), .QN(n82) );
  NOR2X0 U209 ( .IN1(n95), .IN2(n130), .QN(N48) );
  NOR2X0 U210 ( .IN1(n94), .IN2(n130), .QN(N47) );
  NOR2X0 U211 ( .IN1(n93), .IN2(n130), .QN(N46) );
  INVX0 U212 ( .INP(rst), .ZN(n129) );
  INVX0 U213 ( .INP(n5), .ZN(n307) );
  INVX0 U214 ( .INP(n206), .ZN(n194) );
  NAND3X0 U215 ( .IN1(n206), .IN2(n58), .IN3(n29), .QN(n231) );
  NAND2X0 U216 ( .IN1(n254), .IN2(n253), .QN(sel_poly[6]) );
  INVX0 U217 ( .INP(pre_output[9]), .ZN(n262) );
  NAND2X0 U218 ( .IN1(input_shifted[2]), .IN2(n42), .QN(n216) );
  NAND2X0 U219 ( .IN1(input_shifted[2]), .IN2(n59), .QN(n206) );
  INVX0 U220 ( .INP(n47), .ZN(n264) );
  INVX0 U221 ( .INP(pre_output[6]), .ZN(n265) );
  INVX0 U222 ( .INP(n65), .ZN(n263) );
  NAND2X0 U223 ( .IN1(n141), .IN2(n241), .QN(n212) );
  NAND2X0 U224 ( .IN1(n203), .IN2(n202), .QN(n241) );
  NAND2X0 U225 ( .IN1(n18), .IN2(n30), .QN(n289) );
  NAND2X0 U226 ( .IN1(n251), .IN2(n257), .QN(sel_poly[7]) );
  NOR2X0 U227 ( .IN1(n251), .IN2(n36), .QN(n244) );
  NOR2X0 U228 ( .IN1(input_2[6]), .IN2(n90), .QN(n157) );
  NAND2X0 U229 ( .IN1(n132), .IN2(n101), .QN(n173) );
  INVX0 U230 ( .INP(n133), .ZN(n161) );
  AND2X1 U231 ( .IN1(n160), .IN2(n83), .Q(n153) );
  NAND4X0 U232 ( .IN1(n99), .IN2(n135), .IN3(n97), .IN4(n98), .QN(n165) );
  NAND2X0 U233 ( .IN1(n149), .IN2(n55), .QN(n181) );
  INVX0 U234 ( .INP(n40), .ZN(n155) );
  NAND2X0 U235 ( .IN1(n153), .IN2(n163), .QN(n184) );
  INVX0 U236 ( .INP(input_shifted[7]), .ZN(n227) );
  XOR2X2 U237 ( .IN1(n172), .IN2(n182), .Q(shift_amount[1]) );
  INVX0 U238 ( .INP(n246), .ZN(n236) );
  INVX0 U239 ( .INP(input_shifted[2]), .ZN(n215) );
  NAND2X0 U240 ( .IN1(n251), .IN2(n252), .QN(n253) );
  NAND2X0 U241 ( .IN1(n258), .IN2(n232), .QN(n224) );
  NAND2X0 U242 ( .IN1(n259), .IN2(n258), .QN(n260) );
  INVX0 U243 ( .INP(n98), .ZN(n158) );
  NAND2X0 U244 ( .IN1(n142), .IN2(n256), .QN(n249) );
  INVX0 U245 ( .INP(n91), .ZN(n176) );
  INVX0 U246 ( .INP(input_shifted[4]), .ZN(n234) );
  NAND2X0 U247 ( .IN1(pre_output[1]), .IN2(pre_output[2]), .QN(n301) );
  NAND2X0 U248 ( .IN1(n91), .IN2(n4), .QN(n171) );
  INVX0 U249 ( .INP(N228), .ZN(n235) );
  INVX0 U250 ( .INP(n97), .ZN(n159) );
  NAND2X0 U251 ( .IN1(pre_output[0]), .IN2(n34), .QN(n299) );
  NAND2X0 U252 ( .IN1(pre_output[0]), .IN2(pre_output[1]), .QN(n295) );
  OAI21X2 U253 ( .IN1(n181), .IN2(n180), .IN3(n179), .QN(shift_amount[2]) );
  NAND2X0 U254 ( .IN1(input_shifted[6]), .IN2(N228), .QN(n218) );
  NAND2X0 U255 ( .IN1(n174), .IN2(n173), .QN(n167) );
  NAND2X0 U256 ( .IN1(n204), .IN2(n212), .QN(n210) );
  NAND2X0 U257 ( .IN1(n51), .IN2(n221), .QN(n230) );
  NAND2X0 U258 ( .IN1(n65), .IN2(n78), .QN(n308) );
  NAND2X0 U259 ( .IN1(input_shifted[4]), .IN2(n58), .QN(n193) );
  NAND2X0 U260 ( .IN1(n51), .IN2(n29), .QN(n202) );
  NAND2X0 U261 ( .IN1(n234), .IN2(n227), .QN(n200) );
  NAND2X0 U262 ( .IN1(n234), .IN2(n235), .QN(n213) );
  NOR2X0 U263 ( .IN1(n19), .IN2(n51), .QN(n248) );
  NAND2X0 U264 ( .IN1(n101), .IN2(n40), .QN(n174) );
  NAND2X0 U265 ( .IN1(n77), .IN2(n47), .QN(n283) );
  NAND2X0 U266 ( .IN1(input_shifted[2]), .IN2(N220), .QN(n188) );
  NAND2X0 U267 ( .IN1(n215), .IN2(N220), .QN(n205) );
  MUX21X1 U268 ( .IN1(n161), .IN2(\input [5]), .S(start), .Q(n122) );
  MUX21X1 U269 ( .IN1(input_2[10]), .IN2(\input [10]), .S(start), .Q(n127) );
  NAND4X0 U270 ( .IN1(n157), .IN2(n83), .IN3(n133), .IN4(n162), .QN(n180) );
  AO21X1 U271 ( .IN1(input_2[0]), .IN2(n135), .IN3(input_2[2]), .Q(n160) );
  NAND4X0 U272 ( .IN1(n57), .IN2(n167), .IN3(n184), .IN4(n180), .QN(n172) );
  NAND4X0 U273 ( .IN1(n102), .IN2(n173), .IN3(n91), .IN4(n174), .QN(n175) );
  NAND3X0 U274 ( .IN1(n154), .IN2(n147), .IN3(n86), .QN(n178) );
  AO21X1 U276 ( .IN1(n59), .IN2(n215), .IN3(n185), .Q(n189) );
  XOR2X1 U277 ( .IN1(n188), .IN2(n187), .Q(n191) );
  XOR3X1 U278 ( .IN1(n51), .IN2(n29), .IN3(n192), .Q(n198) );
  OA21X1 U279 ( .IN1(n194), .IN2(n193), .IN3(n205), .Q(n195) );
  XOR2X1 U280 ( .IN1(n196), .IN2(n195), .Q(n197) );
  XOR3X1 U281 ( .IN1(n31), .IN2(n54), .IN3(n21), .Q(n208) );
  XOR2X1 U282 ( .IN1(n208), .IN2(n207), .Q(n209) );
  AO21X1 U283 ( .IN1(n59), .IN2(n62), .IN3(n13), .Q(n211) );
  AO21X1 U284 ( .IN1(n212), .IN2(n211), .IN3(n76), .Q(n226) );
  XOR2X1 U285 ( .IN1(n255), .IN2(n224), .Q(n225) );
  AO21X1 U286 ( .IN1(n23), .IN2(n32), .IN3(n36), .Q(n228) );
  AO21X1 U287 ( .IN1(n143), .IN2(n231), .IN3(n230), .Q(n233) );
  AO21X1 U288 ( .IN1(n236), .IN2(n62), .IN3(n146), .Q(n245) );
  NAND4X0 U289 ( .IN1(n242), .IN2(n141), .IN3(n38), .IN4(n240), .QN(n243) );
  AO21X1 U290 ( .IN1(n255), .IN2(n140), .IN3(n261), .Q(n257) );
  MUX21X1 U292 ( .IN1(out_reg_enable), .IN2(state), .S(n82), .Q(n137) );
  NAND2X1 U293 ( .IN1(n263), .IN2(n264), .QN(n271) );
  NAND2X1 U294 ( .IN1(n264), .IN2(n265), .QN(n284) );
  NAND2X1 U295 ( .IN1(n265), .IN2(n298), .QN(n270) );
  NAND2X1 U296 ( .IN1(n295), .IN2(n301), .QN(n294) );
  AO22X1 U297 ( .IN1(n66), .IN2(n34), .IN3(n267), .IN4(n294), .Q(n293) );
  AO22X1 U298 ( .IN1(n66), .IN2(n18), .IN3(n268), .IN4(n293), .Q(n290) );
  AO21X1 U299 ( .IN1(n290), .IN2(n302), .IN3(n269), .Q(n288) );
  AO22X1 U300 ( .IN1(n30), .IN2(n77), .IN3(n270), .IN4(n288), .Q(n285) );
  AO21X1 U301 ( .IN1(n284), .IN2(n285), .IN3(n304), .Q(n282) );
  AO22X1 U302 ( .IN1(n47), .IN2(n65), .IN3(n271), .IN4(n282), .Q(n279) );
  AO21X1 U303 ( .IN1(n278), .IN2(n279), .IN3(n272), .Q(n277) );
  AO22X1 U304 ( .IN1(n73), .IN2(n78), .IN3(n273), .IN4(n277), .Q(n276) );
  AO22X1 U305 ( .IN1(n73), .IN2(n64), .IN3(n274), .IN4(n276), .Q(n275) );
  XOR2X1 U306 ( .IN1(n275), .IN2(n64), .Q(N255) );
  XOR3X1 U307 ( .IN1(n64), .IN2(n73), .IN3(n276), .Q(N254) );
  XOR3X1 U308 ( .IN1(n73), .IN2(n78), .IN3(n277), .Q(N253) );
  MUX21X1 U309 ( .IN1(n281), .IN2(n280), .S(n279), .Q(N252) );
  XOR3X1 U310 ( .IN1(n47), .IN2(n65), .IN3(n282), .Q(N251) );
  XOR3X1 U311 ( .IN1(n30), .IN2(n77), .IN3(n288), .Q(N249) );
  XOR2X1 U312 ( .IN1(n18), .IN2(n30), .Q(n292) );
  MUX21X1 U313 ( .IN1(n292), .IN2(n291), .S(n290), .Q(N248) );
  XOR3X1 U314 ( .IN1(n66), .IN2(n18), .IN3(n293), .Q(N247) );
  XOR3X1 U315 ( .IN1(n66), .IN2(n34), .IN3(n294), .Q(N246) );
  XOR2X1 U316 ( .IN1(n45), .IN2(n34), .Q(n296) );
  NAND4X0 U317 ( .IN1(n301), .IN2(n300), .IN3(n299), .IN4(n298), .QN(n303) );
  NAND4X0 U318 ( .IN1(n304), .IN2(n78), .IN3(n303), .IN4(n302), .QN(n306) );
  NAND4X0 U319 ( .IN1(n308), .IN2(n307), .IN3(n306), .IN4(n305), .QN(n309) );
  NOR3X0 U320 ( .IN1(input_2[9]), .IN2(input_2[8]), .IN3(input_2[7]), .QN(n313) );
  NOR3X0 U321 ( .IN1(input_2[4]), .IN2(n88), .IN3(input_2[3]), .QN(n311) );
  NAND4X0 U322 ( .IN1(n313), .IN2(n312), .IN3(n311), .IN4(n310), .QN(n327) );
  AO21X1 U323 ( .IN1(n325), .IN2(pre_output[0]), .IN3(n151), .Q(n314) );
  AO221X1 U324 ( .IN1(N256), .IN2(n150), .IN3(\output [0]), .IN4(n324), .IN5(
        n314), .Q(n105) );
  AO21X1 U325 ( .IN1(n325), .IN2(n45), .IN3(n151), .Q(n315) );
  AO221X1 U326 ( .IN1(N257), .IN2(n150), .IN3(\output [1]), .IN4(n324), .IN5(
        n315), .Q(n106) );
  AO21X1 U327 ( .IN1(n325), .IN2(n34), .IN3(n151), .Q(n316) );
  AO221X1 U328 ( .IN1(N258), .IN2(n150), .IN3(\output [2]), .IN4(n324), .IN5(
        n316), .Q(n107) );
  AO21X1 U329 ( .IN1(n66), .IN2(n325), .IN3(n151), .Q(n317) );
  AO221X1 U330 ( .IN1(N259), .IN2(n150), .IN3(\output [3]), .IN4(n324), .IN5(
        n317), .Q(n108) );
  AO21X1 U331 ( .IN1(n18), .IN2(n325), .IN3(n151), .Q(n318) );
  AO221X1 U332 ( .IN1(N260), .IN2(n150), .IN3(\output [4]), .IN4(n324), .IN5(
        n318), .Q(n109) );
  AO21X1 U333 ( .IN1(n30), .IN2(n325), .IN3(n151), .Q(n319) );
  AO221X1 U334 ( .IN1(N261), .IN2(n150), .IN3(\output [5]), .IN4(n324), .IN5(
        n319), .Q(n110) );
  AO21X1 U335 ( .IN1(n325), .IN2(n77), .IN3(n151), .Q(n320) );
  AO221X1 U336 ( .IN1(N262), .IN2(n150), .IN3(\output [6]), .IN4(n324), .IN5(
        n320), .Q(n111) );
  AO21X1 U337 ( .IN1(n325), .IN2(n47), .IN3(n151), .Q(n321) );
  AO221X1 U338 ( .IN1(N263), .IN2(n150), .IN3(\output [7]), .IN4(n324), .IN5(
        n321), .Q(n112) );
  AO21X1 U339 ( .IN1(n325), .IN2(n65), .IN3(n151), .Q(n322) );
  AO221X1 U340 ( .IN1(N264), .IN2(n150), .IN3(\output [8]), .IN4(n324), .IN5(
        n322), .Q(n113) );
  AO221X1 U341 ( .IN1(n325), .IN2(n78), .IN3(\output [9]), .IN4(n324), .IN5(
        n151), .Q(n323) );
  AO21X1 U342 ( .IN1(N265), .IN2(n150), .IN3(n323), .Q(n114) );
  AO221X1 U343 ( .IN1(n73), .IN2(n325), .IN3(\output [10]), .IN4(n324), .IN5(
        n151), .Q(n326) );
  AO21X1 U344 ( .IN1(n150), .IN2(N266), .IN3(n326), .Q(n115) );
endmodule


module qr_decomp_ctl_mux_1 ( .in_A_r({\in_A_r[0][11] , \in_A_r[0][10] , 
        \in_A_r[0][9] , \in_A_r[0][8] , \in_A_r[0][7] , \in_A_r[0][6] , 
        \in_A_r[0][5] , \in_A_r[0][4] , \in_A_r[0][3] , \in_A_r[0][2] , 
        \in_A_r[0][1] , \in_A_r[0][0] , \in_A_r[1][11] , \in_A_r[1][10] , 
        \in_A_r[1][9] , \in_A_r[1][8] , \in_A_r[1][7] , \in_A_r[1][6] , 
        \in_A_r[1][5] , \in_A_r[1][4] , \in_A_r[1][3] , \in_A_r[1][2] , 
        \in_A_r[1][1] , \in_A_r[1][0] , \in_A_r[2][11] , \in_A_r[2][10] , 
        \in_A_r[2][9] , \in_A_r[2][8] , \in_A_r[2][7] , \in_A_r[2][6] , 
        \in_A_r[2][5] , \in_A_r[2][4] , \in_A_r[2][3] , \in_A_r[2][2] , 
        \in_A_r[2][1] , \in_A_r[2][0] , \in_A_r[3][11] , \in_A_r[3][10] , 
        \in_A_r[3][9] , \in_A_r[3][8] , \in_A_r[3][7] , \in_A_r[3][6] , 
        \in_A_r[3][5] , \in_A_r[3][4] , \in_A_r[3][3] , \in_A_r[3][2] , 
        \in_A_r[3][1] , \in_A_r[3][0] }), .out_r_vec_mult({
        \out_r_vec_mult[0][11] , \out_r_vec_mult[0][10] , 
        \out_r_vec_mult[0][9] , \out_r_vec_mult[0][8] , \out_r_vec_mult[0][7] , 
        \out_r_vec_mult[0][6] , \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] , 
        \out_r_vec_mult[0][3] , \out_r_vec_mult[0][2] , \out_r_vec_mult[0][1] , 
        \out_r_vec_mult[0][0] , \out_r_vec_mult[1][11] , 
        \out_r_vec_mult[1][10] , \out_r_vec_mult[1][9] , 
        \out_r_vec_mult[1][8] , \out_r_vec_mult[1][7] , \out_r_vec_mult[1][6] , 
        \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] , \out_r_vec_mult[1][3] , 
        \out_r_vec_mult[1][2] , \out_r_vec_mult[1][1] , \out_r_vec_mult[1][0] , 
        \out_r_vec_mult[2][11] , \out_r_vec_mult[2][10] , 
        \out_r_vec_mult[2][9] , \out_r_vec_mult[2][8] , \out_r_vec_mult[2][7] , 
        \out_r_vec_mult[2][6] , \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] , 
        \out_r_vec_mult[2][3] , \out_r_vec_mult[2][2] , \out_r_vec_mult[2][1] , 
        \out_r_vec_mult[2][0] , \out_r_vec_mult[3][11] , 
        \out_r_vec_mult[3][10] , \out_r_vec_mult[3][9] , 
        \out_r_vec_mult[3][8] , \out_r_vec_mult[3][7] , \out_r_vec_mult[3][6] , 
        \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] , \out_r_vec_mult[3][3] , 
        \out_r_vec_mult[3][2] , \out_r_vec_mult[3][1] , \out_r_vec_mult[3][0] 
        }), .out_r_vec_sub({\out_r_vec_sub[0][11] , \out_r_vec_sub[0][10] , 
        \out_r_vec_sub[0][9] , \out_r_vec_sub[0][8] , \out_r_vec_sub[0][7] , 
        \out_r_vec_sub[0][6] , \out_r_vec_sub[0][5] , \out_r_vec_sub[0][4] , 
        \out_r_vec_sub[0][3] , \out_r_vec_sub[0][2] , \out_r_vec_sub[0][1] , 
        \out_r_vec_sub[0][0] , \out_r_vec_sub[1][11] , \out_r_vec_sub[1][10] , 
        \out_r_vec_sub[1][9] , \out_r_vec_sub[1][8] , \out_r_vec_sub[1][7] , 
        \out_r_vec_sub[1][6] , \out_r_vec_sub[1][5] , \out_r_vec_sub[1][4] , 
        \out_r_vec_sub[1][3] , \out_r_vec_sub[1][2] , \out_r_vec_sub[1][1] , 
        \out_r_vec_sub[1][0] , \out_r_vec_sub[2][11] , \out_r_vec_sub[2][10] , 
        \out_r_vec_sub[2][9] , \out_r_vec_sub[2][8] , \out_r_vec_sub[2][7] , 
        \out_r_vec_sub[2][6] , \out_r_vec_sub[2][5] , \out_r_vec_sub[2][4] , 
        \out_r_vec_sub[2][3] , \out_r_vec_sub[2][2] , \out_r_vec_sub[2][1] , 
        \out_r_vec_sub[2][0] , \out_r_vec_sub[3][11] , \out_r_vec_sub[3][10] , 
        \out_r_vec_sub[3][9] , \out_r_vec_sub[3][8] , \out_r_vec_sub[3][7] , 
        \out_r_vec_sub[3][6] , \out_r_vec_sub[3][5] , \out_r_vec_sub[3][4] , 
        \out_r_vec_sub[3][3] , \out_r_vec_sub[3][2] , \out_r_vec_sub[3][1] , 
        \out_r_vec_sub[3][0] }), .vec_in_r_AQ_mux({\vec_in_r_AQ_mux[0][11] , 
        \vec_in_r_AQ_mux[0][10] , \vec_in_r_AQ_mux[0][9] , 
        \vec_in_r_AQ_mux[0][8] , \vec_in_r_AQ_mux[0][7] , 
        \vec_in_r_AQ_mux[0][6] , \vec_in_r_AQ_mux[0][5] , 
        \vec_in_r_AQ_mux[0][4] , \vec_in_r_AQ_mux[0][3] , 
        \vec_in_r_AQ_mux[0][2] , \vec_in_r_AQ_mux[0][1] , 
        \vec_in_r_AQ_mux[0][0] , \vec_in_r_AQ_mux[1][11] , 
        \vec_in_r_AQ_mux[1][10] , \vec_in_r_AQ_mux[1][9] , 
        \vec_in_r_AQ_mux[1][8] , \vec_in_r_AQ_mux[1][7] , 
        \vec_in_r_AQ_mux[1][6] , \vec_in_r_AQ_mux[1][5] , 
        \vec_in_r_AQ_mux[1][4] , \vec_in_r_AQ_mux[1][3] , 
        \vec_in_r_AQ_mux[1][2] , \vec_in_r_AQ_mux[1][1] , 
        \vec_in_r_AQ_mux[1][0] , \vec_in_r_AQ_mux[2][11] , 
        \vec_in_r_AQ_mux[2][10] , \vec_in_r_AQ_mux[2][9] , 
        \vec_in_r_AQ_mux[2][8] , \vec_in_r_AQ_mux[2][7] , 
        \vec_in_r_AQ_mux[2][6] , \vec_in_r_AQ_mux[2][5] , 
        \vec_in_r_AQ_mux[2][4] , \vec_in_r_AQ_mux[2][3] , 
        \vec_in_r_AQ_mux[2][2] , \vec_in_r_AQ_mux[2][1] , 
        \vec_in_r_AQ_mux[2][0] , \vec_in_r_AQ_mux[3][11] , 
        \vec_in_r_AQ_mux[3][10] , \vec_in_r_AQ_mux[3][9] , 
        \vec_in_r_AQ_mux[3][8] , \vec_in_r_AQ_mux[3][7] , 
        \vec_in_r_AQ_mux[3][6] , \vec_in_r_AQ_mux[3][5] , 
        \vec_in_r_AQ_mux[3][4] , \vec_in_r_AQ_mux[3][3] , 
        \vec_in_r_AQ_mux[3][2] , \vec_in_r_AQ_mux[3][1] , 
        \vec_in_r_AQ_mux[3][0] }), .in_A_i({\in_A_i[0][11] , \in_A_i[0][10] , 
        \in_A_i[0][9] , \in_A_i[0][8] , \in_A_i[0][7] , \in_A_i[0][6] , 
        \in_A_i[0][5] , \in_A_i[0][4] , \in_A_i[0][3] , \in_A_i[0][2] , 
        \in_A_i[0][1] , \in_A_i[0][0] , \in_A_i[1][11] , \in_A_i[1][10] , 
        \in_A_i[1][9] , \in_A_i[1][8] , \in_A_i[1][7] , \in_A_i[1][6] , 
        \in_A_i[1][5] , \in_A_i[1][4] , \in_A_i[1][3] , \in_A_i[1][2] , 
        \in_A_i[1][1] , \in_A_i[1][0] , \in_A_i[2][11] , \in_A_i[2][10] , 
        \in_A_i[2][9] , \in_A_i[2][8] , \in_A_i[2][7] , \in_A_i[2][6] , 
        \in_A_i[2][5] , \in_A_i[2][4] , \in_A_i[2][3] , \in_A_i[2][2] , 
        \in_A_i[2][1] , \in_A_i[2][0] , \in_A_i[3][11] , \in_A_i[3][10] , 
        \in_A_i[3][9] , \in_A_i[3][8] , \in_A_i[3][7] , \in_A_i[3][6] , 
        \in_A_i[3][5] , \in_A_i[3][4] , \in_A_i[3][3] , \in_A_i[3][2] , 
        \in_A_i[3][1] , \in_A_i[3][0] }), .out_i_vec_mult({
        \out_i_vec_mult[0][11] , \out_i_vec_mult[0][10] , 
        \out_i_vec_mult[0][9] , \out_i_vec_mult[0][8] , \out_i_vec_mult[0][7] , 
        \out_i_vec_mult[0][6] , \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] , 
        \out_i_vec_mult[0][3] , \out_i_vec_mult[0][2] , \out_i_vec_mult[0][1] , 
        \out_i_vec_mult[0][0] , \out_i_vec_mult[1][11] , 
        \out_i_vec_mult[1][10] , \out_i_vec_mult[1][9] , 
        \out_i_vec_mult[1][8] , \out_i_vec_mult[1][7] , \out_i_vec_mult[1][6] , 
        \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] , \out_i_vec_mult[1][3] , 
        \out_i_vec_mult[1][2] , \out_i_vec_mult[1][1] , \out_i_vec_mult[1][0] , 
        \out_i_vec_mult[2][11] , \out_i_vec_mult[2][10] , 
        \out_i_vec_mult[2][9] , \out_i_vec_mult[2][8] , \out_i_vec_mult[2][7] , 
        \out_i_vec_mult[2][6] , \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] , 
        \out_i_vec_mult[2][3] , \out_i_vec_mult[2][2] , \out_i_vec_mult[2][1] , 
        \out_i_vec_mult[2][0] , \out_i_vec_mult[3][11] , 
        \out_i_vec_mult[3][10] , \out_i_vec_mult[3][9] , 
        \out_i_vec_mult[3][8] , \out_i_vec_mult[3][7] , \out_i_vec_mult[3][6] , 
        \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] , \out_i_vec_mult[3][3] , 
        \out_i_vec_mult[3][2] , \out_i_vec_mult[3][1] , \out_i_vec_mult[3][0] 
        }), .out_i_vec_sub({\out_i_vec_sub[0][11] , \out_i_vec_sub[0][10] , 
        \out_i_vec_sub[0][9] , \out_i_vec_sub[0][8] , \out_i_vec_sub[0][7] , 
        \out_i_vec_sub[0][6] , \out_i_vec_sub[0][5] , \out_i_vec_sub[0][4] , 
        \out_i_vec_sub[0][3] , \out_i_vec_sub[0][2] , \out_i_vec_sub[0][1] , 
        \out_i_vec_sub[0][0] , \out_i_vec_sub[1][11] , \out_i_vec_sub[1][10] , 
        \out_i_vec_sub[1][9] , \out_i_vec_sub[1][8] , \out_i_vec_sub[1][7] , 
        \out_i_vec_sub[1][6] , \out_i_vec_sub[1][5] , \out_i_vec_sub[1][4] , 
        \out_i_vec_sub[1][3] , \out_i_vec_sub[1][2] , \out_i_vec_sub[1][1] , 
        \out_i_vec_sub[1][0] , \out_i_vec_sub[2][11] , \out_i_vec_sub[2][10] , 
        \out_i_vec_sub[2][9] , \out_i_vec_sub[2][8] , \out_i_vec_sub[2][7] , 
        \out_i_vec_sub[2][6] , \out_i_vec_sub[2][5] , \out_i_vec_sub[2][4] , 
        \out_i_vec_sub[2][3] , \out_i_vec_sub[2][2] , \out_i_vec_sub[2][1] , 
        \out_i_vec_sub[2][0] , \out_i_vec_sub[3][11] , \out_i_vec_sub[3][10] , 
        \out_i_vec_sub[3][9] , \out_i_vec_sub[3][8] , \out_i_vec_sub[3][7] , 
        \out_i_vec_sub[3][6] , \out_i_vec_sub[3][5] , \out_i_vec_sub[3][4] , 
        \out_i_vec_sub[3][3] , \out_i_vec_sub[3][2] , \out_i_vec_sub[3][1] , 
        \out_i_vec_sub[3][0] }), .vec_in_i_AQ_mux({\vec_in_i_AQ_mux[0][11] , 
        \vec_in_i_AQ_mux[0][10] , \vec_in_i_AQ_mux[0][9] , 
        \vec_in_i_AQ_mux[0][8] , \vec_in_i_AQ_mux[0][7] , 
        \vec_in_i_AQ_mux[0][6] , \vec_in_i_AQ_mux[0][5] , 
        \vec_in_i_AQ_mux[0][4] , \vec_in_i_AQ_mux[0][3] , 
        \vec_in_i_AQ_mux[0][2] , \vec_in_i_AQ_mux[0][1] , 
        \vec_in_i_AQ_mux[0][0] , \vec_in_i_AQ_mux[1][11] , 
        \vec_in_i_AQ_mux[1][10] , \vec_in_i_AQ_mux[1][9] , 
        \vec_in_i_AQ_mux[1][8] , \vec_in_i_AQ_mux[1][7] , 
        \vec_in_i_AQ_mux[1][6] , \vec_in_i_AQ_mux[1][5] , 
        \vec_in_i_AQ_mux[1][4] , \vec_in_i_AQ_mux[1][3] , 
        \vec_in_i_AQ_mux[1][2] , \vec_in_i_AQ_mux[1][1] , 
        \vec_in_i_AQ_mux[1][0] , \vec_in_i_AQ_mux[2][11] , 
        \vec_in_i_AQ_mux[2][10] , \vec_in_i_AQ_mux[2][9] , 
        \vec_in_i_AQ_mux[2][8] , \vec_in_i_AQ_mux[2][7] , 
        \vec_in_i_AQ_mux[2][6] , \vec_in_i_AQ_mux[2][5] , 
        \vec_in_i_AQ_mux[2][4] , \vec_in_i_AQ_mux[2][3] , 
        \vec_in_i_AQ_mux[2][2] , \vec_in_i_AQ_mux[2][1] , 
        \vec_in_i_AQ_mux[2][0] , \vec_in_i_AQ_mux[3][11] , 
        \vec_in_i_AQ_mux[3][10] , \vec_in_i_AQ_mux[3][9] , 
        \vec_in_i_AQ_mux[3][8] , \vec_in_i_AQ_mux[3][7] , 
        \vec_in_i_AQ_mux[3][6] , \vec_in_i_AQ_mux[3][5] , 
        \vec_in_i_AQ_mux[3][4] , \vec_in_i_AQ_mux[3][3] , 
        \vec_in_i_AQ_mux[3][2] , \vec_in_i_AQ_mux[3][1] , 
        \vec_in_i_AQ_mux[3][0] }), vec_in_AQ_sel, col_sel_AQ, col_sel_AQ2_int, 
        col_sel_AQ2_mux, col_sel_AQ2_sel, wr_A, wr_en_AQ_int, wr_en_AQ_mux, 
        wr_en_AQ_sel, out_mult, out_inner_prod_r, single_in_r_R_mux, 
        out_inner_prod_i, single_in_i_R_mux, single_in_R_sel, col_sel_R, 
        col_sel_R_int, col_sel_R_mux, col_sel_R_sel, out_inv_sqrt, 
        in_b_r_vec_mult_mux, in_b_i_vec_mult_mux, in_b_vec_mult_sel, 
        w_col_sel_AQ_int, w_col_sel_AQ_mux, w_col_sel_AQ_sel, 
        vec_in_r_AQ_mux_0, single_out_r_AQ, vec_in_i_AQ_mux_0, single_out_i_AQ, 
        in_a_r_inner_prod_mux, in_a_i_inner_prod_mux, in_a_inner_prod_sel, 
        out_r_vec_sub_0, single_out_r_AQ2, out_i_vec_sub_0, single_out_i_AQ2, 
        in_b_r_inner_prod_mux, in_b_i_inner_prod_mux, in_b_inner_prod_sel );
  input [1:0] vec_in_AQ_sel;
  input [1:0] col_sel_AQ;
  input [1:0] col_sel_AQ2_int;
  output [1:0] col_sel_AQ2_mux;
  input [11:0] out_mult;
  input [11:0] out_inner_prod_r;
  output [11:0] single_in_r_R_mux;
  input [11:0] out_inner_prod_i;
  output [11:0] single_in_i_R_mux;
  input [1:0] col_sel_R;
  input [1:0] col_sel_R_int;
  output [1:0] col_sel_R_mux;
  input [11:0] out_inv_sqrt;
  output [11:0] in_b_r_vec_mult_mux;
  output [11:0] in_b_i_vec_mult_mux;
  input [1:0] w_col_sel_AQ_int;
  output [1:0] w_col_sel_AQ_mux;
  input [11:0] vec_in_r_AQ_mux_0;
  input [11:0] single_out_r_AQ;
  input [11:0] vec_in_i_AQ_mux_0;
  input [11:0] single_out_i_AQ;
  output [11:0] in_a_r_inner_prod_mux;
  output [11:0] in_a_i_inner_prod_mux;
  input [11:0] out_r_vec_sub_0;
  input [11:0] single_out_r_AQ2;
  input [11:0] out_i_vec_sub_0;
  input [11:0] single_out_i_AQ2;
  output [11:0] in_b_r_inner_prod_mux;
  output [11:0] in_b_i_inner_prod_mux;
  input \in_A_r[0][11] , \in_A_r[0][10] , \in_A_r[0][9] , \in_A_r[0][8] ,
         \in_A_r[0][7] , \in_A_r[0][6] , \in_A_r[0][5] , \in_A_r[0][4] ,
         \in_A_r[0][3] , \in_A_r[0][2] , \in_A_r[0][1] , \in_A_r[0][0] ,
         \in_A_r[1][11] , \in_A_r[1][10] , \in_A_r[1][9] , \in_A_r[1][8] ,
         \in_A_r[1][7] , \in_A_r[1][6] , \in_A_r[1][5] , \in_A_r[1][4] ,
         \in_A_r[1][3] , \in_A_r[1][2] , \in_A_r[1][1] , \in_A_r[1][0] ,
         \in_A_r[2][11] , \in_A_r[2][10] , \in_A_r[2][9] , \in_A_r[2][8] ,
         \in_A_r[2][7] , \in_A_r[2][6] , \in_A_r[2][5] , \in_A_r[2][4] ,
         \in_A_r[2][3] , \in_A_r[2][2] , \in_A_r[2][1] , \in_A_r[2][0] ,
         \in_A_r[3][11] , \in_A_r[3][10] , \in_A_r[3][9] , \in_A_r[3][8] ,
         \in_A_r[3][7] , \in_A_r[3][6] , \in_A_r[3][5] , \in_A_r[3][4] ,
         \in_A_r[3][3] , \in_A_r[3][2] , \in_A_r[3][1] , \in_A_r[3][0] ,
         \out_r_vec_mult[0][11] , \out_r_vec_mult[0][10] ,
         \out_r_vec_mult[0][9] , \out_r_vec_mult[0][8] ,
         \out_r_vec_mult[0][7] , \out_r_vec_mult[0][6] ,
         \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] ,
         \out_r_vec_mult[0][3] , \out_r_vec_mult[0][2] ,
         \out_r_vec_mult[0][1] , \out_r_vec_mult[0][0] ,
         \out_r_vec_mult[1][11] , \out_r_vec_mult[1][10] ,
         \out_r_vec_mult[1][9] , \out_r_vec_mult[1][8] ,
         \out_r_vec_mult[1][7] , \out_r_vec_mult[1][6] ,
         \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] ,
         \out_r_vec_mult[1][3] , \out_r_vec_mult[1][2] ,
         \out_r_vec_mult[1][1] , \out_r_vec_mult[1][0] ,
         \out_r_vec_mult[2][11] , \out_r_vec_mult[2][10] ,
         \out_r_vec_mult[2][9] , \out_r_vec_mult[2][8] ,
         \out_r_vec_mult[2][7] , \out_r_vec_mult[2][6] ,
         \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] ,
         \out_r_vec_mult[2][3] , \out_r_vec_mult[2][2] ,
         \out_r_vec_mult[2][1] , \out_r_vec_mult[2][0] ,
         \out_r_vec_mult[3][11] , \out_r_vec_mult[3][10] ,
         \out_r_vec_mult[3][9] , \out_r_vec_mult[3][8] ,
         \out_r_vec_mult[3][7] , \out_r_vec_mult[3][6] ,
         \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] ,
         \out_r_vec_mult[3][3] , \out_r_vec_mult[3][2] ,
         \out_r_vec_mult[3][1] , \out_r_vec_mult[3][0] ,
         \out_r_vec_sub[0][11] , \out_r_vec_sub[0][10] , \out_r_vec_sub[0][9] ,
         \out_r_vec_sub[0][8] , \out_r_vec_sub[0][7] , \out_r_vec_sub[0][6] ,
         \out_r_vec_sub[0][5] , \out_r_vec_sub[0][4] , \out_r_vec_sub[0][3] ,
         \out_r_vec_sub[0][2] , \out_r_vec_sub[0][1] , \out_r_vec_sub[0][0] ,
         \out_r_vec_sub[1][11] , \out_r_vec_sub[1][10] , \out_r_vec_sub[1][9] ,
         \out_r_vec_sub[1][8] , \out_r_vec_sub[1][7] , \out_r_vec_sub[1][6] ,
         \out_r_vec_sub[1][5] , \out_r_vec_sub[1][4] , \out_r_vec_sub[1][3] ,
         \out_r_vec_sub[1][2] , \out_r_vec_sub[1][1] , \out_r_vec_sub[1][0] ,
         \out_r_vec_sub[2][11] , \out_r_vec_sub[2][10] , \out_r_vec_sub[2][9] ,
         \out_r_vec_sub[2][8] , \out_r_vec_sub[2][7] , \out_r_vec_sub[2][6] ,
         \out_r_vec_sub[2][5] , \out_r_vec_sub[2][4] , \out_r_vec_sub[2][3] ,
         \out_r_vec_sub[2][2] , \out_r_vec_sub[2][1] , \out_r_vec_sub[2][0] ,
         \out_r_vec_sub[3][11] , \out_r_vec_sub[3][10] , \out_r_vec_sub[3][9] ,
         \out_r_vec_sub[3][8] , \out_r_vec_sub[3][7] , \out_r_vec_sub[3][6] ,
         \out_r_vec_sub[3][5] , \out_r_vec_sub[3][4] , \out_r_vec_sub[3][3] ,
         \out_r_vec_sub[3][2] , \out_r_vec_sub[3][1] , \out_r_vec_sub[3][0] ,
         \in_A_i[0][11] , \in_A_i[0][10] , \in_A_i[0][9] , \in_A_i[0][8] ,
         \in_A_i[0][7] , \in_A_i[0][6] , \in_A_i[0][5] , \in_A_i[0][4] ,
         \in_A_i[0][3] , \in_A_i[0][2] , \in_A_i[0][1] , \in_A_i[0][0] ,
         \in_A_i[1][11] , \in_A_i[1][10] , \in_A_i[1][9] , \in_A_i[1][8] ,
         \in_A_i[1][7] , \in_A_i[1][6] , \in_A_i[1][5] , \in_A_i[1][4] ,
         \in_A_i[1][3] , \in_A_i[1][2] , \in_A_i[1][1] , \in_A_i[1][0] ,
         \in_A_i[2][11] , \in_A_i[2][10] , \in_A_i[2][9] , \in_A_i[2][8] ,
         \in_A_i[2][7] , \in_A_i[2][6] , \in_A_i[2][5] , \in_A_i[2][4] ,
         \in_A_i[2][3] , \in_A_i[2][2] , \in_A_i[2][1] , \in_A_i[2][0] ,
         \in_A_i[3][11] , \in_A_i[3][10] , \in_A_i[3][9] , \in_A_i[3][8] ,
         \in_A_i[3][7] , \in_A_i[3][6] , \in_A_i[3][5] , \in_A_i[3][4] ,
         \in_A_i[3][3] , \in_A_i[3][2] , \in_A_i[3][1] , \in_A_i[3][0] ,
         \out_i_vec_mult[0][11] , \out_i_vec_mult[0][10] ,
         \out_i_vec_mult[0][9] , \out_i_vec_mult[0][8] ,
         \out_i_vec_mult[0][7] , \out_i_vec_mult[0][6] ,
         \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] ,
         \out_i_vec_mult[0][3] , \out_i_vec_mult[0][2] ,
         \out_i_vec_mult[0][1] , \out_i_vec_mult[0][0] ,
         \out_i_vec_mult[1][11] , \out_i_vec_mult[1][10] ,
         \out_i_vec_mult[1][9] , \out_i_vec_mult[1][8] ,
         \out_i_vec_mult[1][7] , \out_i_vec_mult[1][6] ,
         \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] ,
         \out_i_vec_mult[1][3] , \out_i_vec_mult[1][2] ,
         \out_i_vec_mult[1][1] , \out_i_vec_mult[1][0] ,
         \out_i_vec_mult[2][11] , \out_i_vec_mult[2][10] ,
         \out_i_vec_mult[2][9] , \out_i_vec_mult[2][8] ,
         \out_i_vec_mult[2][7] , \out_i_vec_mult[2][6] ,
         \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] ,
         \out_i_vec_mult[2][3] , \out_i_vec_mult[2][2] ,
         \out_i_vec_mult[2][1] , \out_i_vec_mult[2][0] ,
         \out_i_vec_mult[3][11] , \out_i_vec_mult[3][10] ,
         \out_i_vec_mult[3][9] , \out_i_vec_mult[3][8] ,
         \out_i_vec_mult[3][7] , \out_i_vec_mult[3][6] ,
         \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] ,
         \out_i_vec_mult[3][3] , \out_i_vec_mult[3][2] ,
         \out_i_vec_mult[3][1] , \out_i_vec_mult[3][0] ,
         \out_i_vec_sub[0][11] , \out_i_vec_sub[0][10] , \out_i_vec_sub[0][9] ,
         \out_i_vec_sub[0][8] , \out_i_vec_sub[0][7] , \out_i_vec_sub[0][6] ,
         \out_i_vec_sub[0][5] , \out_i_vec_sub[0][4] , \out_i_vec_sub[0][3] ,
         \out_i_vec_sub[0][2] , \out_i_vec_sub[0][1] , \out_i_vec_sub[0][0] ,
         \out_i_vec_sub[1][11] , \out_i_vec_sub[1][10] , \out_i_vec_sub[1][9] ,
         \out_i_vec_sub[1][8] , \out_i_vec_sub[1][7] , \out_i_vec_sub[1][6] ,
         \out_i_vec_sub[1][5] , \out_i_vec_sub[1][4] , \out_i_vec_sub[1][3] ,
         \out_i_vec_sub[1][2] , \out_i_vec_sub[1][1] , \out_i_vec_sub[1][0] ,
         \out_i_vec_sub[2][11] , \out_i_vec_sub[2][10] , \out_i_vec_sub[2][9] ,
         \out_i_vec_sub[2][8] , \out_i_vec_sub[2][7] , \out_i_vec_sub[2][6] ,
         \out_i_vec_sub[2][5] , \out_i_vec_sub[2][4] , \out_i_vec_sub[2][3] ,
         \out_i_vec_sub[2][2] , \out_i_vec_sub[2][1] , \out_i_vec_sub[2][0] ,
         \out_i_vec_sub[3][11] , \out_i_vec_sub[3][10] , \out_i_vec_sub[3][9] ,
         \out_i_vec_sub[3][8] , \out_i_vec_sub[3][7] , \out_i_vec_sub[3][6] ,
         \out_i_vec_sub[3][5] , \out_i_vec_sub[3][4] , \out_i_vec_sub[3][3] ,
         \out_i_vec_sub[3][2] , \out_i_vec_sub[3][1] , \out_i_vec_sub[3][0] ,
         col_sel_AQ2_sel, wr_A, wr_en_AQ_int, wr_en_AQ_sel, single_in_R_sel,
         col_sel_R_sel, in_b_vec_mult_sel, w_col_sel_AQ_sel,
         in_a_inner_prod_sel, in_b_inner_prod_sel;
  output \vec_in_r_AQ_mux[0][11] , \vec_in_r_AQ_mux[0][10] ,
         \vec_in_r_AQ_mux[0][9] , \vec_in_r_AQ_mux[0][8] ,
         \vec_in_r_AQ_mux[0][7] , \vec_in_r_AQ_mux[0][6] ,
         \vec_in_r_AQ_mux[0][5] , \vec_in_r_AQ_mux[0][4] ,
         \vec_in_r_AQ_mux[0][3] , \vec_in_r_AQ_mux[0][2] ,
         \vec_in_r_AQ_mux[0][1] , \vec_in_r_AQ_mux[0][0] ,
         \vec_in_r_AQ_mux[1][11] , \vec_in_r_AQ_mux[1][10] ,
         \vec_in_r_AQ_mux[1][9] , \vec_in_r_AQ_mux[1][8] ,
         \vec_in_r_AQ_mux[1][7] , \vec_in_r_AQ_mux[1][6] ,
         \vec_in_r_AQ_mux[1][5] , \vec_in_r_AQ_mux[1][4] ,
         \vec_in_r_AQ_mux[1][3] , \vec_in_r_AQ_mux[1][2] ,
         \vec_in_r_AQ_mux[1][1] , \vec_in_r_AQ_mux[1][0] ,
         \vec_in_r_AQ_mux[2][11] , \vec_in_r_AQ_mux[2][10] ,
         \vec_in_r_AQ_mux[2][9] , \vec_in_r_AQ_mux[2][8] ,
         \vec_in_r_AQ_mux[2][7] , \vec_in_r_AQ_mux[2][6] ,
         \vec_in_r_AQ_mux[2][5] , \vec_in_r_AQ_mux[2][4] ,
         \vec_in_r_AQ_mux[2][3] , \vec_in_r_AQ_mux[2][2] ,
         \vec_in_r_AQ_mux[2][1] , \vec_in_r_AQ_mux[2][0] ,
         \vec_in_r_AQ_mux[3][11] , \vec_in_r_AQ_mux[3][10] ,
         \vec_in_r_AQ_mux[3][9] , \vec_in_r_AQ_mux[3][8] ,
         \vec_in_r_AQ_mux[3][7] , \vec_in_r_AQ_mux[3][6] ,
         \vec_in_r_AQ_mux[3][5] , \vec_in_r_AQ_mux[3][4] ,
         \vec_in_r_AQ_mux[3][3] , \vec_in_r_AQ_mux[3][2] ,
         \vec_in_r_AQ_mux[3][1] , \vec_in_r_AQ_mux[3][0] ,
         \vec_in_i_AQ_mux[0][11] , \vec_in_i_AQ_mux[0][10] ,
         \vec_in_i_AQ_mux[0][9] , \vec_in_i_AQ_mux[0][8] ,
         \vec_in_i_AQ_mux[0][7] , \vec_in_i_AQ_mux[0][6] ,
         \vec_in_i_AQ_mux[0][5] , \vec_in_i_AQ_mux[0][4] ,
         \vec_in_i_AQ_mux[0][3] , \vec_in_i_AQ_mux[0][2] ,
         \vec_in_i_AQ_mux[0][1] , \vec_in_i_AQ_mux[0][0] ,
         \vec_in_i_AQ_mux[1][11] , \vec_in_i_AQ_mux[1][10] ,
         \vec_in_i_AQ_mux[1][9] , \vec_in_i_AQ_mux[1][8] ,
         \vec_in_i_AQ_mux[1][7] , \vec_in_i_AQ_mux[1][6] ,
         \vec_in_i_AQ_mux[1][5] , \vec_in_i_AQ_mux[1][4] ,
         \vec_in_i_AQ_mux[1][3] , \vec_in_i_AQ_mux[1][2] ,
         \vec_in_i_AQ_mux[1][1] , \vec_in_i_AQ_mux[1][0] ,
         \vec_in_i_AQ_mux[2][11] , \vec_in_i_AQ_mux[2][10] ,
         \vec_in_i_AQ_mux[2][9] , \vec_in_i_AQ_mux[2][8] ,
         \vec_in_i_AQ_mux[2][7] , \vec_in_i_AQ_mux[2][6] ,
         \vec_in_i_AQ_mux[2][5] , \vec_in_i_AQ_mux[2][4] ,
         \vec_in_i_AQ_mux[2][3] , \vec_in_i_AQ_mux[2][2] ,
         \vec_in_i_AQ_mux[2][1] , \vec_in_i_AQ_mux[2][0] ,
         \vec_in_i_AQ_mux[3][11] , \vec_in_i_AQ_mux[3][10] ,
         \vec_in_i_AQ_mux[3][9] , \vec_in_i_AQ_mux[3][8] ,
         \vec_in_i_AQ_mux[3][7] , \vec_in_i_AQ_mux[3][6] ,
         \vec_in_i_AQ_mux[3][5] , \vec_in_i_AQ_mux[3][4] ,
         \vec_in_i_AQ_mux[3][3] , \vec_in_i_AQ_mux[3][2] ,
         \vec_in_i_AQ_mux[3][1] , \vec_in_i_AQ_mux[3][0] , wr_en_AQ_mux;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;

  AO22X1 U50 ( .IN1(wr_en_AQ_sel), .IN2(wr_en_AQ_int), .IN3(wr_A), .IN4(n45), 
        .Q(wr_en_AQ_mux) );
  AO22X1 U51 ( .IN1(w_col_sel_AQ_sel), .IN2(w_col_sel_AQ_int[1]), .IN3(
        col_sel_AQ[1]), .IN4(n44), .Q(w_col_sel_AQ_mux[1]) );
  AO22X1 U52 ( .IN1(w_col_sel_AQ_int[0]), .IN2(w_col_sel_AQ_sel), .IN3(
        col_sel_AQ[0]), .IN4(n44), .Q(w_col_sel_AQ_mux[0]) );
  AO22X1 U149 ( .IN1(out_mult[9]), .IN2(n26), .IN3(single_in_R_sel), .IN4(
        out_inner_prod_r[9]), .Q(single_in_r_R_mux[9]) );
  AO22X1 U150 ( .IN1(out_mult[8]), .IN2(n27), .IN3(out_inner_prod_r[8]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[8]) );
  AO22X1 U151 ( .IN1(out_mult[7]), .IN2(n27), .IN3(out_inner_prod_r[7]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[7]) );
  AO22X1 U152 ( .IN1(out_mult[6]), .IN2(n27), .IN3(out_inner_prod_r[6]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[6]) );
  AO22X1 U153 ( .IN1(out_mult[5]), .IN2(n27), .IN3(out_inner_prod_r[5]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[5]) );
  AO22X1 U158 ( .IN1(out_mult[11]), .IN2(n27), .IN3(out_inner_prod_r[11]), 
        .IN4(single_in_R_sel), .Q(single_in_r_R_mux[11]) );
  AO22X1 U159 ( .IN1(out_mult[10]), .IN2(n27), .IN3(out_inner_prod_r[10]), 
        .IN4(single_in_R_sel), .Q(single_in_r_R_mux[10]) );
  AO22X1 U160 ( .IN1(out_mult[0]), .IN2(n27), .IN3(out_inner_prod_r[0]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[0]) );
  AO22X1 U163 ( .IN1(out_inv_sqrt[7]), .IN2(n33), .IN3(out_inner_prod_r[7]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[7]) );
  AO22X1 U165 ( .IN1(out_inv_sqrt[5]), .IN2(n33), .IN3(out_inner_prod_r[5]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[5]) );
  AO22X1 U221 ( .IN1(col_sel_R_sel), .IN2(col_sel_R_int[1]), .IN3(col_sel_R[1]), .IN4(n42), .Q(col_sel_R_mux[1]) );
  AO22X1 U222 ( .IN1(col_sel_R_int[0]), .IN2(col_sel_R_sel), .IN3(col_sel_R[0]), .IN4(n42), .Q(col_sel_R_mux[0]) );
  AO22X1 U223 ( .IN1(col_sel_AQ[1]), .IN2(n41), .IN3(col_sel_AQ2_sel), .IN4(
        col_sel_AQ2_int[1]), .Q(col_sel_AQ2_mux[1]) );
  AO22X1 U224 ( .IN1(col_sel_AQ[0]), .IN2(n41), .IN3(col_sel_AQ2_int[0]), 
        .IN4(col_sel_AQ2_sel), .Q(col_sel_AQ2_mux[0]) );
  AO22X1 U2 ( .IN1(out_inv_sqrt[1]), .IN2(n33), .IN3(out_inner_prod_r[1]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[1]) );
  AO22X2 U3 ( .IN1(out_inv_sqrt[8]), .IN2(n33), .IN3(out_inner_prod_r[8]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[8]) );
  AO22X2 U4 ( .IN1(out_inv_sqrt[4]), .IN2(n33), .IN3(out_inner_prod_r[4]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[4]) );
  AO22X2 U5 ( .IN1(out_mult[4]), .IN2(n27), .IN3(out_inner_prod_r[4]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[4]) );
  AO22X2 U6 ( .IN1(out_inv_sqrt[3]), .IN2(n33), .IN3(out_inner_prod_r[3]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[3]) );
  AO22X2 U7 ( .IN1(out_mult[3]), .IN2(n27), .IN3(out_inner_prod_r[3]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[3]) );
  AO22X2 U8 ( .IN1(out_inv_sqrt[2]), .IN2(n33), .IN3(out_inner_prod_r[2]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[2]) );
  AO22X2 U9 ( .IN1(out_mult[2]), .IN2(n27), .IN3(out_inner_prod_r[2]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[2]) );
  AO22X2 U10 ( .IN1(out_mult[1]), .IN2(n27), .IN3(out_inner_prod_r[1]), .IN4(
        single_in_R_sel), .Q(single_in_r_R_mux[1]) );
  NBUFFX2 U11 ( .INP(n1), .Z(n10) );
  NBUFFX2 U12 ( .INP(n1), .Z(n11) );
  NBUFFX2 U13 ( .INP(n39), .Z(n2) );
  NBUFFX2 U14 ( .INP(n39), .Z(n3) );
  NBUFFX2 U15 ( .INP(n40), .Z(n18) );
  NBUFFX2 U16 ( .INP(n40), .Z(n19) );
  NBUFFX2 U17 ( .INP(n1), .Z(n14) );
  NBUFFX2 U18 ( .INP(n1), .Z(n13) );
  NBUFFX2 U19 ( .INP(n1), .Z(n12) );
  NBUFFX2 U20 ( .INP(n1), .Z(n17) );
  NBUFFX2 U21 ( .INP(n1), .Z(n16) );
  NBUFFX2 U22 ( .INP(n1), .Z(n15) );
  NBUFFX2 U23 ( .INP(n39), .Z(n6) );
  NBUFFX2 U24 ( .INP(n40), .Z(n22) );
  NBUFFX2 U25 ( .INP(n40), .Z(n21) );
  NBUFFX2 U26 ( .INP(n40), .Z(n20) );
  NBUFFX2 U27 ( .INP(n40), .Z(n25) );
  NBUFFX2 U28 ( .INP(n40), .Z(n24) );
  NBUFFX2 U29 ( .INP(n40), .Z(n23) );
  NBUFFX2 U30 ( .INP(n39), .Z(n5) );
  NBUFFX2 U31 ( .INP(n39), .Z(n4) );
  NBUFFX2 U32 ( .INP(n39), .Z(n9) );
  NBUFFX2 U33 ( .INP(n39), .Z(n8) );
  NBUFFX2 U34 ( .INP(n39), .Z(n7) );
  NBUFFX2 U35 ( .INP(n43), .Z(n26) );
  NBUFFX2 U36 ( .INP(n43), .Z(n27) );
  NOR2X0 U37 ( .IN1(n26), .IN2(n46), .QN(single_in_i_R_mux[0]) );
  NOR2X0 U38 ( .IN1(n26), .IN2(n47), .QN(single_in_i_R_mux[1]) );
  NOR2X0 U39 ( .IN1(n26), .IN2(n48), .QN(single_in_i_R_mux[2]) );
  NOR2X0 U40 ( .IN1(n26), .IN2(n49), .QN(single_in_i_R_mux[3]) );
  NOR2X0 U41 ( .IN1(n26), .IN2(n50), .QN(single_in_i_R_mux[4]) );
  NOR2X0 U42 ( .IN1(n26), .IN2(n51), .QN(single_in_i_R_mux[5]) );
  NOR2X0 U43 ( .IN1(n26), .IN2(n56), .QN(single_in_i_R_mux[10]) );
  NOR2X0 U44 ( .IN1(n26), .IN2(n57), .QN(single_in_i_R_mux[11]) );
  NOR2X0 U45 ( .IN1(n27), .IN2(n52), .QN(single_in_i_R_mux[6]) );
  NOR2X0 U46 ( .IN1(n27), .IN2(n53), .QN(single_in_i_R_mux[7]) );
  NOR2X0 U47 ( .IN1(n27), .IN2(n54), .QN(single_in_i_R_mux[8]) );
  NOR2X0 U48 ( .IN1(n27), .IN2(n55), .QN(single_in_i_R_mux[9]) );
  INVX0 U49 ( .INP(n38), .ZN(n39) );
  INVX0 U53 ( .INP(n37), .ZN(n40) );
  AND2X1 U54 ( .IN1(n37), .IN2(n38), .Q(n1) );
  INVX0 U55 ( .INP(n34), .ZN(n32) );
  NOR2X0 U56 ( .IN1(n32), .IN2(n46), .QN(in_b_i_vec_mult_mux[0]) );
  INVX0 U57 ( .INP(single_in_R_sel), .ZN(n43) );
  INVX0 U58 ( .INP(col_sel_R_sel), .ZN(n42) );
  INVX0 U59 ( .INP(col_sel_AQ2_sel), .ZN(n41) );
  INVX0 U60 ( .INP(vec_in_AQ_sel[0]), .ZN(n35) );
  INVX0 U61 ( .INP(vec_in_AQ_sel[1]), .ZN(n36) );
  INVX0 U62 ( .INP(w_col_sel_AQ_sel), .ZN(n44) );
  INVX0 U63 ( .INP(wr_en_AQ_sel), .ZN(n45) );
  NBUFFX2 U64 ( .INP(in_a_inner_prod_sel), .Z(n30) );
  NBUFFX2 U65 ( .INP(in_a_inner_prod_sel), .Z(n31) );
  NBUFFX2 U66 ( .INP(in_b_inner_prod_sel), .Z(n29) );
  NBUFFX2 U67 ( .INP(in_b_inner_prod_sel), .Z(n28) );
  INVX0 U68 ( .INP(out_inner_prod_i[0]), .ZN(n46) );
  INVX0 U69 ( .INP(out_inner_prod_i[11]), .ZN(n57) );
  INVX0 U70 ( .INP(out_inner_prod_i[7]), .ZN(n53) );
  INVX0 U71 ( .INP(out_inner_prod_i[6]), .ZN(n52) );
  INVX0 U72 ( .INP(out_inner_prod_i[8]), .ZN(n54) );
  INVX0 U73 ( .INP(out_inner_prod_i[9]), .ZN(n55) );
  INVX0 U74 ( .INP(out_inner_prod_i[1]), .ZN(n47) );
  INVX0 U75 ( .INP(out_inner_prod_i[2]), .ZN(n48) );
  INVX0 U76 ( .INP(out_inner_prod_i[3]), .ZN(n49) );
  INVX0 U77 ( .INP(out_inner_prod_i[4]), .ZN(n50) );
  INVX0 U78 ( .INP(out_inner_prod_i[5]), .ZN(n51) );
  INVX0 U79 ( .INP(out_inner_prod_i[10]), .ZN(n56) );
  AO22X1 U80 ( .IN1(out_inv_sqrt[0]), .IN2(n33), .IN3(out_inner_prod_r[0]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[0]) );
  AO22X1 U81 ( .IN1(out_inv_sqrt[6]), .IN2(n33), .IN3(out_inner_prod_r[6]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[6]) );
  AO22X1 U82 ( .IN1(out_inv_sqrt[11]), .IN2(n33), .IN3(out_inner_prod_r[11]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[11]) );
  AO22X1 U83 ( .IN1(out_inv_sqrt[9]), .IN2(n33), .IN3(out_inner_prod_r[9]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[9]) );
  AO22X1 U84 ( .IN1(out_inv_sqrt[10]), .IN2(n33), .IN3(out_inner_prod_r[10]), 
        .IN4(n34), .Q(in_b_r_vec_mult_mux[10]) );
  NOR2X0 U85 ( .IN1(n32), .IN2(n57), .QN(in_b_i_vec_mult_mux[11]) );
  NOR2X0 U86 ( .IN1(n32), .IN2(n52), .QN(in_b_i_vec_mult_mux[6]) );
  NOR2X0 U87 ( .IN1(n32), .IN2(n53), .QN(in_b_i_vec_mult_mux[7]) );
  NOR2X0 U88 ( .IN1(n32), .IN2(n56), .QN(in_b_i_vec_mult_mux[10]) );
  NOR2X0 U89 ( .IN1(n32), .IN2(n54), .QN(in_b_i_vec_mult_mux[8]) );
  NOR2X0 U90 ( .IN1(n32), .IN2(n55), .QN(in_b_i_vec_mult_mux[9]) );
  NOR2X0 U91 ( .IN1(n32), .IN2(n51), .QN(in_b_i_vec_mult_mux[5]) );
  NOR2X0 U92 ( .IN1(n32), .IN2(n50), .QN(in_b_i_vec_mult_mux[4]) );
  NOR2X0 U93 ( .IN1(n32), .IN2(n49), .QN(in_b_i_vec_mult_mux[3]) );
  NOR2X0 U94 ( .IN1(n32), .IN2(n47), .QN(in_b_i_vec_mult_mux[1]) );
  NOR2X0 U95 ( .IN1(n32), .IN2(n48), .QN(in_b_i_vec_mult_mux[2]) );
  INVX0 U96 ( .INP(n34), .ZN(n33) );
  INVX0 U97 ( .INP(in_b_vec_mult_sel), .ZN(n34) );
  MUX21X1 U98 ( .IN1(out_i_vec_sub_0[0]), .IN2(single_out_i_AQ2[0]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[0]) );
  MUX21X1 U99 ( .IN1(out_i_vec_sub_0[1]), .IN2(single_out_i_AQ2[1]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[1]) );
  MUX21X1 U100 ( .IN1(out_i_vec_sub_0[2]), .IN2(single_out_i_AQ2[2]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[2]) );
  MUX21X1 U101 ( .IN1(out_i_vec_sub_0[3]), .IN2(single_out_i_AQ2[3]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[3]) );
  MUX21X1 U102 ( .IN1(out_i_vec_sub_0[4]), .IN2(single_out_i_AQ2[4]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[4]) );
  MUX21X1 U103 ( .IN1(out_i_vec_sub_0[5]), .IN2(single_out_i_AQ2[5]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[5]) );
  MUX21X1 U104 ( .IN1(out_i_vec_sub_0[6]), .IN2(single_out_i_AQ2[6]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[6]) );
  MUX21X1 U105 ( .IN1(out_i_vec_sub_0[7]), .IN2(single_out_i_AQ2[7]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[7]) );
  MUX21X1 U106 ( .IN1(out_i_vec_sub_0[8]), .IN2(single_out_i_AQ2[8]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[8]) );
  MUX21X1 U107 ( .IN1(out_i_vec_sub_0[9]), .IN2(single_out_i_AQ2[9]), .S(n28), 
        .Q(in_b_i_inner_prod_mux[9]) );
  MUX21X1 U108 ( .IN1(out_i_vec_sub_0[10]), .IN2(single_out_i_AQ2[10]), .S(n28), .Q(in_b_i_inner_prod_mux[10]) );
  MUX21X1 U109 ( .IN1(out_i_vec_sub_0[11]), .IN2(single_out_i_AQ2[11]), .S(n28), .Q(in_b_i_inner_prod_mux[11]) );
  MUX21X1 U110 ( .IN1(out_r_vec_sub_0[0]), .IN2(single_out_r_AQ2[0]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[0]) );
  MUX21X1 U111 ( .IN1(out_r_vec_sub_0[1]), .IN2(single_out_r_AQ2[1]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[1]) );
  MUX21X1 U112 ( .IN1(out_r_vec_sub_0[2]), .IN2(single_out_r_AQ2[2]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[2]) );
  MUX21X1 U113 ( .IN1(out_r_vec_sub_0[3]), .IN2(single_out_r_AQ2[3]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[3]) );
  MUX21X1 U114 ( .IN1(out_r_vec_sub_0[4]), .IN2(single_out_r_AQ2[4]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[4]) );
  MUX21X1 U115 ( .IN1(out_r_vec_sub_0[5]), .IN2(single_out_r_AQ2[5]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[5]) );
  MUX21X1 U116 ( .IN1(out_r_vec_sub_0[6]), .IN2(single_out_r_AQ2[6]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[6]) );
  MUX21X1 U117 ( .IN1(out_r_vec_sub_0[7]), .IN2(single_out_r_AQ2[7]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[7]) );
  MUX21X1 U118 ( .IN1(out_r_vec_sub_0[8]), .IN2(single_out_r_AQ2[8]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[8]) );
  MUX21X1 U119 ( .IN1(out_r_vec_sub_0[9]), .IN2(single_out_r_AQ2[9]), .S(n29), 
        .Q(in_b_r_inner_prod_mux[9]) );
  MUX21X1 U120 ( .IN1(out_r_vec_sub_0[10]), .IN2(single_out_r_AQ2[10]), .S(n29), .Q(in_b_r_inner_prod_mux[10]) );
  MUX21X1 U121 ( .IN1(out_r_vec_sub_0[11]), .IN2(single_out_r_AQ2[11]), .S(n29), .Q(in_b_r_inner_prod_mux[11]) );
  MUX21X1 U122 ( .IN1(vec_in_i_AQ_mux_0[0]), .IN2(single_out_i_AQ[0]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[0]) );
  MUX21X1 U123 ( .IN1(vec_in_i_AQ_mux_0[1]), .IN2(single_out_i_AQ[1]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[1]) );
  MUX21X1 U124 ( .IN1(vec_in_i_AQ_mux_0[2]), .IN2(single_out_i_AQ[2]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[2]) );
  MUX21X1 U125 ( .IN1(vec_in_i_AQ_mux_0[3]), .IN2(single_out_i_AQ[3]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[3]) );
  MUX21X1 U126 ( .IN1(vec_in_i_AQ_mux_0[4]), .IN2(single_out_i_AQ[4]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[4]) );
  MUX21X1 U127 ( .IN1(vec_in_i_AQ_mux_0[5]), .IN2(single_out_i_AQ[5]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[5]) );
  MUX21X1 U128 ( .IN1(vec_in_i_AQ_mux_0[6]), .IN2(single_out_i_AQ[6]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[6]) );
  MUX21X1 U129 ( .IN1(vec_in_i_AQ_mux_0[7]), .IN2(single_out_i_AQ[7]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[7]) );
  MUX21X1 U130 ( .IN1(vec_in_i_AQ_mux_0[8]), .IN2(single_out_i_AQ[8]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[8]) );
  MUX21X1 U131 ( .IN1(vec_in_i_AQ_mux_0[9]), .IN2(single_out_i_AQ[9]), .S(n30), 
        .Q(in_a_i_inner_prod_mux[9]) );
  MUX21X1 U132 ( .IN1(vec_in_i_AQ_mux_0[10]), .IN2(single_out_i_AQ[10]), .S(
        n30), .Q(in_a_i_inner_prod_mux[10]) );
  MUX21X1 U133 ( .IN1(vec_in_i_AQ_mux_0[11]), .IN2(single_out_i_AQ[11]), .S(
        n30), .Q(in_a_i_inner_prod_mux[11]) );
  MUX21X1 U134 ( .IN1(vec_in_r_AQ_mux_0[0]), .IN2(single_out_r_AQ[0]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[0]) );
  MUX21X1 U135 ( .IN1(vec_in_r_AQ_mux_0[1]), .IN2(single_out_r_AQ[1]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[1]) );
  MUX21X1 U136 ( .IN1(vec_in_r_AQ_mux_0[2]), .IN2(single_out_r_AQ[2]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[2]) );
  MUX21X1 U137 ( .IN1(vec_in_r_AQ_mux_0[3]), .IN2(single_out_r_AQ[3]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[3]) );
  MUX21X1 U138 ( .IN1(vec_in_r_AQ_mux_0[4]), .IN2(single_out_r_AQ[4]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[4]) );
  MUX21X1 U139 ( .IN1(vec_in_r_AQ_mux_0[5]), .IN2(single_out_r_AQ[5]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[5]) );
  MUX21X1 U140 ( .IN1(vec_in_r_AQ_mux_0[6]), .IN2(single_out_r_AQ[6]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[6]) );
  MUX21X1 U141 ( .IN1(vec_in_r_AQ_mux_0[7]), .IN2(single_out_r_AQ[7]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[7]) );
  MUX21X1 U142 ( .IN1(vec_in_r_AQ_mux_0[8]), .IN2(single_out_r_AQ[8]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[8]) );
  MUX21X1 U143 ( .IN1(vec_in_r_AQ_mux_0[9]), .IN2(single_out_r_AQ[9]), .S(n31), 
        .Q(in_a_r_inner_prod_mux[9]) );
  MUX21X1 U144 ( .IN1(vec_in_r_AQ_mux_0[10]), .IN2(single_out_r_AQ[10]), .S(
        n31), .Q(in_a_r_inner_prod_mux[10]) );
  MUX21X1 U145 ( .IN1(vec_in_r_AQ_mux_0[11]), .IN2(single_out_r_AQ[11]), .S(
        n31), .Q(in_a_r_inner_prod_mux[11]) );
  NAND2X1 U146 ( .IN1(n36), .IN2(n35), .QN(n37) );
  NAND2X1 U147 ( .IN1(vec_in_AQ_sel[0]), .IN2(n36), .QN(n38) );
  AO222X1 U148 ( .IN1(\in_A_i[3][0] ), .IN2(n25), .IN3(\out_i_vec_sub[3][0] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][0] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][0] ) );
  AO222X1 U154 ( .IN1(\in_A_i[3][1] ), .IN2(n25), .IN3(\out_i_vec_sub[3][1] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][1] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][1] ) );
  AO222X1 U155 ( .IN1(\in_A_i[3][2] ), .IN2(n25), .IN3(\out_i_vec_sub[3][2] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][2] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][2] ) );
  AO222X1 U156 ( .IN1(\in_A_i[3][3] ), .IN2(n25), .IN3(\out_i_vec_sub[3][3] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][3] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][3] ) );
  AO222X1 U157 ( .IN1(\in_A_i[3][4] ), .IN2(n25), .IN3(\out_i_vec_sub[3][4] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][4] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][4] ) );
  AO222X1 U161 ( .IN1(\in_A_i[3][5] ), .IN2(n25), .IN3(\out_i_vec_sub[3][5] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][5] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][5] ) );
  AO222X1 U162 ( .IN1(\in_A_i[3][6] ), .IN2(n25), .IN3(\out_i_vec_sub[3][6] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][6] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][6] ) );
  AO222X1 U164 ( .IN1(\in_A_i[3][7] ), .IN2(n25), .IN3(\out_i_vec_sub[3][7] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][7] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][7] ) );
  AO222X1 U166 ( .IN1(\in_A_i[3][8] ), .IN2(n25), .IN3(\out_i_vec_sub[3][8] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][8] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][8] ) );
  AO222X1 U167 ( .IN1(\in_A_i[3][9] ), .IN2(n25), .IN3(\out_i_vec_sub[3][9] ), 
        .IN4(n17), .IN5(\out_i_vec_mult[3][9] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][9] ) );
  AO222X1 U168 ( .IN1(\in_A_i[3][10] ), .IN2(n25), .IN3(\out_i_vec_sub[3][10] ), .IN4(n17), .IN5(\out_i_vec_mult[3][10] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][10] ) );
  AO222X1 U169 ( .IN1(\in_A_i[3][11] ), .IN2(n25), .IN3(\out_i_vec_sub[3][11] ), .IN4(n17), .IN5(\out_i_vec_mult[3][11] ), .IN6(n9), .Q(
        \vec_in_i_AQ_mux[3][11] ) );
  AO222X1 U170 ( .IN1(\in_A_i[2][0] ), .IN2(n24), .IN3(\out_i_vec_sub[2][0] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][0] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][0] ) );
  AO222X1 U171 ( .IN1(\in_A_i[2][1] ), .IN2(n24), .IN3(\out_i_vec_sub[2][1] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][1] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][1] ) );
  AO222X1 U172 ( .IN1(\in_A_i[2][2] ), .IN2(n24), .IN3(\out_i_vec_sub[2][2] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][2] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][2] ) );
  AO222X1 U173 ( .IN1(\in_A_i[2][3] ), .IN2(n24), .IN3(\out_i_vec_sub[2][3] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][3] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][3] ) );
  AO222X1 U174 ( .IN1(\in_A_i[2][4] ), .IN2(n24), .IN3(\out_i_vec_sub[2][4] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][4] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][4] ) );
  AO222X1 U175 ( .IN1(\in_A_i[2][5] ), .IN2(n24), .IN3(\out_i_vec_sub[2][5] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][5] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][5] ) );
  AO222X1 U176 ( .IN1(\in_A_i[2][6] ), .IN2(n24), .IN3(\out_i_vec_sub[2][6] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][6] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][6] ) );
  AO222X1 U177 ( .IN1(\in_A_i[2][7] ), .IN2(n24), .IN3(\out_i_vec_sub[2][7] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][7] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][7] ) );
  AO222X1 U178 ( .IN1(\in_A_i[2][8] ), .IN2(n24), .IN3(\out_i_vec_sub[2][8] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][8] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][8] ) );
  AO222X1 U179 ( .IN1(\in_A_i[2][9] ), .IN2(n24), .IN3(\out_i_vec_sub[2][9] ), 
        .IN4(n16), .IN5(\out_i_vec_mult[2][9] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][9] ) );
  AO222X1 U180 ( .IN1(\in_A_i[2][10] ), .IN2(n24), .IN3(\out_i_vec_sub[2][10] ), .IN4(n16), .IN5(\out_i_vec_mult[2][10] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][10] ) );
  AO222X1 U181 ( .IN1(\in_A_i[2][11] ), .IN2(n24), .IN3(\out_i_vec_sub[2][11] ), .IN4(n16), .IN5(\out_i_vec_mult[2][11] ), .IN6(n8), .Q(
        \vec_in_i_AQ_mux[2][11] ) );
  AO222X1 U182 ( .IN1(\in_A_i[1][0] ), .IN2(n23), .IN3(\out_i_vec_sub[1][0] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][0] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][0] ) );
  AO222X1 U183 ( .IN1(\in_A_i[1][1] ), .IN2(n23), .IN3(\out_i_vec_sub[1][1] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][1] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][1] ) );
  AO222X1 U184 ( .IN1(\in_A_i[1][2] ), .IN2(n23), .IN3(\out_i_vec_sub[1][2] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][2] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][2] ) );
  AO222X1 U185 ( .IN1(\in_A_i[1][3] ), .IN2(n23), .IN3(\out_i_vec_sub[1][3] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][3] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][3] ) );
  AO222X1 U186 ( .IN1(\in_A_i[1][4] ), .IN2(n23), .IN3(\out_i_vec_sub[1][4] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][4] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][4] ) );
  AO222X1 U187 ( .IN1(\in_A_i[1][5] ), .IN2(n23), .IN3(\out_i_vec_sub[1][5] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][5] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][5] ) );
  AO222X1 U188 ( .IN1(\in_A_i[1][6] ), .IN2(n23), .IN3(\out_i_vec_sub[1][6] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][6] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][6] ) );
  AO222X1 U189 ( .IN1(\in_A_i[1][7] ), .IN2(n23), .IN3(\out_i_vec_sub[1][7] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][7] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][7] ) );
  AO222X1 U190 ( .IN1(\in_A_i[1][8] ), .IN2(n23), .IN3(\out_i_vec_sub[1][8] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][8] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][8] ) );
  AO222X1 U191 ( .IN1(\in_A_i[1][9] ), .IN2(n23), .IN3(\out_i_vec_sub[1][9] ), 
        .IN4(n15), .IN5(\out_i_vec_mult[1][9] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][9] ) );
  AO222X1 U192 ( .IN1(\in_A_i[1][10] ), .IN2(n23), .IN3(\out_i_vec_sub[1][10] ), .IN4(n15), .IN5(\out_i_vec_mult[1][10] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][10] ) );
  AO222X1 U193 ( .IN1(\in_A_i[1][11] ), .IN2(n23), .IN3(\out_i_vec_sub[1][11] ), .IN4(n15), .IN5(\out_i_vec_mult[1][11] ), .IN6(n7), .Q(
        \vec_in_i_AQ_mux[1][11] ) );
  AO222X1 U194 ( .IN1(\in_A_i[0][0] ), .IN2(n22), .IN3(\out_i_vec_sub[0][0] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][0] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][0] ) );
  AO222X1 U195 ( .IN1(\in_A_i[0][1] ), .IN2(n22), .IN3(\out_i_vec_sub[0][1] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][1] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][1] ) );
  AO222X1 U196 ( .IN1(\in_A_i[0][2] ), .IN2(n22), .IN3(\out_i_vec_sub[0][2] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][2] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][2] ) );
  AO222X1 U197 ( .IN1(\in_A_i[0][3] ), .IN2(n22), .IN3(\out_i_vec_sub[0][3] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][3] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][3] ) );
  AO222X1 U198 ( .IN1(\in_A_i[0][4] ), .IN2(n22), .IN3(\out_i_vec_sub[0][4] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][4] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][4] ) );
  AO222X1 U199 ( .IN1(\in_A_i[0][5] ), .IN2(n22), .IN3(\out_i_vec_sub[0][5] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][5] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][5] ) );
  AO222X1 U200 ( .IN1(\in_A_i[0][6] ), .IN2(n22), .IN3(\out_i_vec_sub[0][6] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][6] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][6] ) );
  AO222X1 U201 ( .IN1(\in_A_i[0][7] ), .IN2(n22), .IN3(\out_i_vec_sub[0][7] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][7] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][7] ) );
  AO222X1 U202 ( .IN1(\in_A_i[0][8] ), .IN2(n22), .IN3(\out_i_vec_sub[0][8] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][8] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][8] ) );
  AO222X1 U203 ( .IN1(\in_A_i[0][9] ), .IN2(n22), .IN3(\out_i_vec_sub[0][9] ), 
        .IN4(n14), .IN5(\out_i_vec_mult[0][9] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][9] ) );
  AO222X1 U204 ( .IN1(\in_A_i[0][10] ), .IN2(n22), .IN3(\out_i_vec_sub[0][10] ), .IN4(n14), .IN5(\out_i_vec_mult[0][10] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][10] ) );
  AO222X1 U205 ( .IN1(\in_A_i[0][11] ), .IN2(n22), .IN3(\out_i_vec_sub[0][11] ), .IN4(n14), .IN5(\out_i_vec_mult[0][11] ), .IN6(n6), .Q(
        \vec_in_i_AQ_mux[0][11] ) );
  AO222X1 U206 ( .IN1(\in_A_r[3][0] ), .IN2(n21), .IN3(\out_r_vec_sub[3][0] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][0] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][0] ) );
  AO222X1 U207 ( .IN1(\in_A_r[3][1] ), .IN2(n21), .IN3(\out_r_vec_sub[3][1] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][1] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][1] ) );
  AO222X1 U208 ( .IN1(\in_A_r[3][2] ), .IN2(n21), .IN3(\out_r_vec_sub[3][2] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][2] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][2] ) );
  AO222X1 U209 ( .IN1(\in_A_r[3][3] ), .IN2(n21), .IN3(\out_r_vec_sub[3][3] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][3] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][3] ) );
  AO222X1 U210 ( .IN1(\in_A_r[3][4] ), .IN2(n21), .IN3(\out_r_vec_sub[3][4] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][4] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][4] ) );
  AO222X1 U211 ( .IN1(\in_A_r[3][5] ), .IN2(n21), .IN3(\out_r_vec_sub[3][5] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][5] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][5] ) );
  AO222X1 U212 ( .IN1(\in_A_r[3][6] ), .IN2(n21), .IN3(\out_r_vec_sub[3][6] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][6] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][6] ) );
  AO222X1 U213 ( .IN1(\in_A_r[3][7] ), .IN2(n21), .IN3(\out_r_vec_sub[3][7] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][7] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][7] ) );
  AO222X1 U214 ( .IN1(\in_A_r[3][8] ), .IN2(n21), .IN3(\out_r_vec_sub[3][8] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][8] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][8] ) );
  AO222X1 U215 ( .IN1(\in_A_r[3][9] ), .IN2(n21), .IN3(\out_r_vec_sub[3][9] ), 
        .IN4(n13), .IN5(\out_r_vec_mult[3][9] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][9] ) );
  AO222X1 U216 ( .IN1(\in_A_r[3][10] ), .IN2(n21), .IN3(\out_r_vec_sub[3][10] ), .IN4(n13), .IN5(\out_r_vec_mult[3][10] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][10] ) );
  AO222X1 U217 ( .IN1(\in_A_r[3][11] ), .IN2(n21), .IN3(\out_r_vec_sub[3][11] ), .IN4(n13), .IN5(\out_r_vec_mult[3][11] ), .IN6(n5), .Q(
        \vec_in_r_AQ_mux[3][11] ) );
  AO222X1 U218 ( .IN1(\in_A_r[2][0] ), .IN2(n20), .IN3(\out_r_vec_sub[2][0] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][0] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][0] ) );
  AO222X1 U219 ( .IN1(\in_A_r[2][1] ), .IN2(n20), .IN3(\out_r_vec_sub[2][1] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][1] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][1] ) );
  AO222X1 U220 ( .IN1(\in_A_r[2][2] ), .IN2(n20), .IN3(\out_r_vec_sub[2][2] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][2] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][2] ) );
  AO222X1 U225 ( .IN1(\in_A_r[2][3] ), .IN2(n20), .IN3(\out_r_vec_sub[2][3] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][3] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][3] ) );
  AO222X1 U226 ( .IN1(\in_A_r[2][4] ), .IN2(n20), .IN3(\out_r_vec_sub[2][4] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][4] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][4] ) );
  AO222X1 U227 ( .IN1(\in_A_r[2][5] ), .IN2(n20), .IN3(\out_r_vec_sub[2][5] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][5] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][5] ) );
  AO222X1 U228 ( .IN1(\in_A_r[2][6] ), .IN2(n20), .IN3(\out_r_vec_sub[2][6] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][6] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][6] ) );
  AO222X1 U229 ( .IN1(\in_A_r[2][7] ), .IN2(n20), .IN3(\out_r_vec_sub[2][7] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][7] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][7] ) );
  AO222X1 U230 ( .IN1(\in_A_r[2][8] ), .IN2(n20), .IN3(\out_r_vec_sub[2][8] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][8] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][8] ) );
  AO222X1 U231 ( .IN1(\in_A_r[2][9] ), .IN2(n20), .IN3(\out_r_vec_sub[2][9] ), 
        .IN4(n12), .IN5(\out_r_vec_mult[2][9] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][9] ) );
  AO222X1 U232 ( .IN1(\in_A_r[2][10] ), .IN2(n20), .IN3(\out_r_vec_sub[2][10] ), .IN4(n12), .IN5(\out_r_vec_mult[2][10] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][10] ) );
  AO222X1 U233 ( .IN1(\in_A_r[2][11] ), .IN2(n20), .IN3(\out_r_vec_sub[2][11] ), .IN4(n12), .IN5(\out_r_vec_mult[2][11] ), .IN6(n4), .Q(
        \vec_in_r_AQ_mux[2][11] ) );
  AO222X1 U234 ( .IN1(\in_A_r[1][0] ), .IN2(n19), .IN3(\out_r_vec_sub[1][0] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][0] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][0] ) );
  AO222X1 U235 ( .IN1(\in_A_r[1][1] ), .IN2(n19), .IN3(\out_r_vec_sub[1][1] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][1] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][1] ) );
  AO222X1 U236 ( .IN1(\in_A_r[1][2] ), .IN2(n19), .IN3(\out_r_vec_sub[1][2] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][2] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][2] ) );
  AO222X1 U237 ( .IN1(\in_A_r[1][3] ), .IN2(n19), .IN3(\out_r_vec_sub[1][3] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][3] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][3] ) );
  AO222X1 U238 ( .IN1(\in_A_r[1][4] ), .IN2(n19), .IN3(\out_r_vec_sub[1][4] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][4] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][4] ) );
  AO222X1 U239 ( .IN1(\in_A_r[1][5] ), .IN2(n19), .IN3(\out_r_vec_sub[1][5] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][5] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][5] ) );
  AO222X1 U240 ( .IN1(\in_A_r[1][6] ), .IN2(n19), .IN3(\out_r_vec_sub[1][6] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][6] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][6] ) );
  AO222X1 U241 ( .IN1(\in_A_r[1][7] ), .IN2(n19), .IN3(\out_r_vec_sub[1][7] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][7] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][7] ) );
  AO222X1 U242 ( .IN1(\in_A_r[1][8] ), .IN2(n19), .IN3(\out_r_vec_sub[1][8] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][8] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][8] ) );
  AO222X1 U243 ( .IN1(\in_A_r[1][9] ), .IN2(n19), .IN3(\out_r_vec_sub[1][9] ), 
        .IN4(n11), .IN5(\out_r_vec_mult[1][9] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][9] ) );
  AO222X1 U244 ( .IN1(\in_A_r[1][10] ), .IN2(n19), .IN3(\out_r_vec_sub[1][10] ), .IN4(n11), .IN5(\out_r_vec_mult[1][10] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][10] ) );
  AO222X1 U245 ( .IN1(\in_A_r[1][11] ), .IN2(n19), .IN3(\out_r_vec_sub[1][11] ), .IN4(n11), .IN5(\out_r_vec_mult[1][11] ), .IN6(n3), .Q(
        \vec_in_r_AQ_mux[1][11] ) );
  AO222X1 U246 ( .IN1(\in_A_r[0][0] ), .IN2(n18), .IN3(\out_r_vec_sub[0][0] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][0] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][0] ) );
  AO222X1 U247 ( .IN1(\in_A_r[0][1] ), .IN2(n18), .IN3(\out_r_vec_sub[0][1] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][1] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][1] ) );
  AO222X1 U248 ( .IN1(\in_A_r[0][2] ), .IN2(n18), .IN3(\out_r_vec_sub[0][2] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][2] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][2] ) );
  AO222X1 U249 ( .IN1(\in_A_r[0][3] ), .IN2(n18), .IN3(\out_r_vec_sub[0][3] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][3] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][3] ) );
  AO222X1 U250 ( .IN1(\in_A_r[0][4] ), .IN2(n18), .IN3(\out_r_vec_sub[0][4] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][4] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][4] ) );
  AO222X1 U251 ( .IN1(\in_A_r[0][5] ), .IN2(n18), .IN3(\out_r_vec_sub[0][5] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][5] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][5] ) );
  AO222X1 U252 ( .IN1(\in_A_r[0][6] ), .IN2(n18), .IN3(\out_r_vec_sub[0][6] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][6] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][6] ) );
  AO222X1 U253 ( .IN1(\in_A_r[0][7] ), .IN2(n18), .IN3(\out_r_vec_sub[0][7] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][7] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][7] ) );
  AO222X1 U254 ( .IN1(\in_A_r[0][8] ), .IN2(n18), .IN3(\out_r_vec_sub[0][8] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][8] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][8] ) );
  AO222X1 U255 ( .IN1(\in_A_r[0][9] ), .IN2(n18), .IN3(\out_r_vec_sub[0][9] ), 
        .IN4(n10), .IN5(\out_r_vec_mult[0][9] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][9] ) );
  AO222X1 U256 ( .IN1(\in_A_r[0][10] ), .IN2(n18), .IN3(\out_r_vec_sub[0][10] ), .IN4(n10), .IN5(\out_r_vec_mult[0][10] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][10] ) );
  AO222X1 U257 ( .IN1(\in_A_r[0][11] ), .IN2(n18), .IN3(\out_r_vec_sub[0][11] ), .IN4(n10), .IN5(\out_r_vec_mult[0][11] ), .IN6(n2), .Q(
        \vec_in_r_AQ_mux[0][11] ) );
endmodule


module qr_decomp_ctl_1 ( clk, rst, start, done_inner_prod, done_inv_sqrt, 
        out_inv_sqrt, reduced_matrix, done, start_inner_prod, start_inv_sqrt, 
        w_in_a_vec_sub, row_sel_AQ2, row_sel_R, wr_en_R, row_sel_AQ_out, 
        red_mat_reg_out, col_sel_AQ_int, col_sel_AQ2_int, in_a_r_mult, 
        col_sel_R_int, w_col_sel_AQ_int, wr_en_AQ_int, vec_in_AQ_sel, 
        col_sel_AQ2_sel, wr_en_AQ_sel, col_sel_R_sel, w_col_sel_AQ_sel, 
        in_a_inner_prod_sel, in_b_inner_prod_sel, single_in_R_sel, 
        in_b_vec_mult_sel );
  input [11:0] out_inv_sqrt;
  output [1:0] row_sel_AQ2;
  output [1:0] row_sel_R;
  output [1:0] row_sel_AQ_out;
  output [1:0] col_sel_AQ_int;
  output [1:0] col_sel_AQ2_int;
  output [11:0] in_a_r_mult;
  output [1:0] col_sel_R_int;
  output [1:0] w_col_sel_AQ_int;
  output [1:0] vec_in_AQ_sel;
  input clk, rst, start, done_inner_prod, done_inv_sqrt, reduced_matrix;
  output done, start_inner_prod, start_inv_sqrt, w_in_a_vec_sub, wr_en_R,
         red_mat_reg_out, wr_en_AQ_int, col_sel_AQ2_sel, wr_en_AQ_sel,
         col_sel_R_sel, w_col_sel_AQ_sel, in_a_inner_prod_sel,
         in_b_inner_prod_sel, single_in_R_sel, in_b_vec_mult_sel;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n40, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n39, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n89, n94, n183, n184;
  wire   [2:0] mult_counter;
  wire   [3:0] state;

  DFFARX1 \state_reg[0]  ( .D(n182), .CLK(clk), .RSTB(n38), .Q(state[0]), .QN(
        n66) );
  DFFARX1 \state_reg[2]  ( .D(n173), .CLK(clk), .RSTB(n37), .Q(state[2]), .QN(
        n64) );
  DFFARX1 col_sel_AQ2_sel_reg ( .D(n172), .CLK(clk), .RSTB(n36), .Q(
        col_sel_AQ2_sel) );
  DFFARX1 col_sel_R_sel_reg ( .D(n171), .CLK(clk), .RSTB(n35), .Q(
        col_sel_R_sel) );
  DFFARX1 pre_red_mat_reg_reg ( .D(n170), .CLK(clk), .RSTB(n34), .Q(
        red_mat_reg_out) );
  DFFARX1 \state_reg[3]  ( .D(n180), .CLK(clk), .RSTB(n33), .Q(state[3]) );
  DFFARX1 \state_reg[1]  ( .D(n174), .CLK(clk), .RSTB(n32), .Q(state[1]), .QN(
        n65) );
  DFFX1 \in_a_r_mult_reg[0]  ( .D(n159), .CLK(clk), .Q(in_a_r_mult[0]) );
  DFFX1 \in_a_r_mult_reg[1]  ( .D(n158), .CLK(clk), .Q(in_a_r_mult[1]) );
  DFFX1 \in_a_r_mult_reg[2]  ( .D(n157), .CLK(clk), .Q(in_a_r_mult[2]) );
  DFFX1 \in_a_r_mult_reg[3]  ( .D(n156), .CLK(clk), .Q(in_a_r_mult[3]) );
  DFFX1 \in_a_r_mult_reg[4]  ( .D(n155), .CLK(clk), .Q(in_a_r_mult[4]) );
  DFFX1 \in_a_r_mult_reg[5]  ( .D(n154), .CLK(clk), .Q(in_a_r_mult[5]) );
  DFFX1 \in_a_r_mult_reg[6]  ( .D(n153), .CLK(clk), .Q(in_a_r_mult[6]) );
  DFFX1 \in_a_r_mult_reg[7]  ( .D(n152), .CLK(clk), .Q(in_a_r_mult[7]) );
  DFFX1 \in_a_r_mult_reg[8]  ( .D(n151), .CLK(clk), .Q(in_a_r_mult[8]) );
  DFFX1 \in_a_r_mult_reg[9]  ( .D(n150), .CLK(clk), .Q(in_a_r_mult[9]) );
  DFFX1 \in_a_r_mult_reg[10]  ( .D(n149), .CLK(clk), .Q(in_a_r_mult[10]) );
  DFFX1 \in_a_r_mult_reg[11]  ( .D(n148), .CLK(clk), .Q(in_a_r_mult[11]) );
  DFFARX1 done_reg ( .D(n147), .CLK(clk), .RSTB(n31), .Q(done) );
  DFFARX1 \mult_counter_reg[0]  ( .D(n165), .CLK(clk), .RSTB(n30), .Q(
        mult_counter[0]) );
  DFFARX1 \mult_counter_reg[1]  ( .D(n164), .CLK(clk), .RSTB(n29), .Q(
        mult_counter[1]) );
  DFFARX1 \mult_counter_reg[2]  ( .D(n179), .CLK(clk), .RSTB(n28), .Q(
        mult_counter[2]) );
  DFFARX1 \k_reg[0]  ( .D(n175), .CLK(clk), .RSTB(n27), .Q(col_sel_AQ_int[0])
         );
  DFFARX1 \row_sel_R_reg[0]  ( .D(n163), .CLK(clk), .RSTB(n26), .Q(
        row_sel_R[0]) );
  DFFARX1 \k_reg[1]  ( .D(n176), .CLK(clk), .RSTB(n25), .Q(col_sel_AQ_int[1])
         );
  DFFARX1 \j_reg[1]  ( .D(n178), .CLK(clk), .RSTB(n24), .Q(col_sel_AQ2_int[1])
         );
  DFFARX1 \j_reg[0]  ( .D(n177), .CLK(clk), .RSTB(n23), .Q(col_sel_AQ2_int[0]), 
        .QN(n40) );
  DFFARX1 \row_sel_R_reg[1]  ( .D(n166), .CLK(clk), .RSTB(n22), .Q(
        row_sel_R[1]) );
  DFFASX1 in_b_inner_prod_sel_reg ( .D(n168), .CLK(clk), .SETB(n21), .Q(
        in_b_inner_prod_sel) );
  DFFASX1 in_a_inner_prod_sel_reg ( .D(n169), .CLK(clk), .SETB(n20), .Q(
        in_a_inner_prod_sel) );
  DFFARX1 \row_sel_AQ_reg[0]  ( .D(n160), .CLK(clk), .RSTB(n19), .Q(
        row_sel_AQ_out[0]) );
  DFFARX1 \row_sel_AQ2_reg[0]  ( .D(n146), .CLK(clk), .RSTB(n18), .Q(
        row_sel_AQ2[0]) );
  DFFARX1 \row_sel_AQ_reg[1]  ( .D(n181), .CLK(clk), .RSTB(n17), .Q(
        row_sel_AQ_out[1]) );
  DFFARX1 \row_sel_AQ2_reg[1]  ( .D(n145), .CLK(clk), .RSTB(n16), .Q(
        row_sel_AQ2[1]) );
  DFFARX1 \col_sel_R_int_reg[1]  ( .D(n161), .CLK(clk), .RSTB(n15), .Q(
        col_sel_R_int[1]) );
  DFFARX1 \col_sel_R_int_reg[0]  ( .D(n162), .CLK(clk), .RSTB(n14), .Q(
        col_sel_R_int[0]) );
  DFFASX1 in_b_vec_mult_sel_reg ( .D(n167), .CLK(clk), .SETB(n13), .Q(
        in_b_vec_mult_sel) );
  DFFARX1 start_inner_prod_reg ( .D(n144), .CLK(clk), .RSTB(n12), .Q(
        start_inner_prod), .QN(n39) );
  DFFARX1 start_inv_sqrt_reg ( .D(n143), .CLK(clk), .RSTB(n11), .Q(
        start_inv_sqrt) );
  DFFARX1 single_in_R_sel_reg ( .D(n142), .CLK(clk), .RSTB(n10), .Q(
        single_in_R_sel) );
  DFFARX1 \vec_in_AQ_sel_reg[1]  ( .D(n141), .CLK(clk), .RSTB(n9), .Q(
        vec_in_AQ_sel[1]) );
  DFFARX1 \vec_in_AQ_sel_reg[0]  ( .D(n140), .CLK(clk), .RSTB(n8), .Q(
        vec_in_AQ_sel[0]) );
  DFFARX1 \w_col_sel_AQ_int_reg[1]  ( .D(n139), .CLK(clk), .RSTB(n7), .Q(
        w_col_sel_AQ_int[1]) );
  DFFARX1 \w_col_sel_AQ_int_reg[0]  ( .D(n138), .CLK(clk), .RSTB(n6), .Q(
        w_col_sel_AQ_int[0]) );
  DFFARX1 w_col_sel_AQ_sel_reg ( .D(n137), .CLK(clk), .RSTB(n5), .Q(
        w_col_sel_AQ_sel) );
  DFFARX1 wr_en_AQ_int_reg ( .D(n136), .CLK(clk), .RSTB(n4), .Q(wr_en_AQ_int)
         );
  DFFARX1 wr_en_R_reg ( .D(n135), .CLK(clk), .RSTB(n3), .Q(wr_en_R) );
  DFFARX1 wr_en_AQ_sel_reg ( .D(n134), .CLK(clk), .RSTB(n2), .Q(wr_en_AQ_sel)
         );
  DFFARX1 w_in_a_vec_sub_reg ( .D(n133), .CLK(clk), .RSTB(n1), .Q(
        w_in_a_vec_sub) );
  AO21X1 U100 ( .IN1(w_in_a_vec_sub), .IN2(n67), .IN3(n62), .Q(n133) );
  AO21X1 U101 ( .IN1(wr_en_AQ_sel), .IN2(n68), .IN3(n94), .Q(n134) );
  AO22X1 U102 ( .IN1(wr_en_R), .IN2(n58), .IN3(n69), .IN4(n70), .Q(n135) );
  NAND4X0 U103 ( .IN1(n67), .IN2(n73), .IN3(n74), .IN4(n75), .QN(n70) );
  AOI21X1 U104 ( .IN1(n89), .IN2(mult_counter[2]), .IN3(n76), .QN(n75) );
  AO22X1 U105 ( .IN1(wr_en_AQ_int), .IN2(n57), .IN3(n77), .IN4(n78), .Q(n136)
         );
  AO21X1 U106 ( .IN1(w_col_sel_AQ_sel), .IN2(n68), .IN3(n94), .Q(n137) );
  AO222X1 U107 ( .IN1(col_sel_AQ_int[0]), .IN2(n81), .IN3(col_sel_AQ2_int[0]), 
        .IN4(n61), .IN5(w_col_sel_AQ_int[0]), .IN6(n79), .Q(n138) );
  AO222X1 U108 ( .IN1(col_sel_AQ_int[1]), .IN2(n81), .IN3(col_sel_AQ2_int[1]), 
        .IN4(n61), .IN5(w_col_sel_AQ_int[1]), .IN6(n79), .Q(n139) );
  AO22X1 U109 ( .IN1(n50), .IN2(n45), .IN3(vec_in_AQ_sel[0]), .IN4(n82), .Q(
        n140) );
  AO22X1 U110 ( .IN1(n63), .IN2(n45), .IN3(vec_in_AQ_sel[1]), .IN4(n82), .Q(
        n141) );
  AO21X1 U111 ( .IN1(single_in_R_sel), .IN2(n83), .IN3(n61), .Q(n142) );
  AO22X1 U112 ( .IN1(n84), .IN2(n85), .IN3(start_inv_sqrt), .IN4(n51), .Q(n143) );
  NAND3X0 U113 ( .IN1(n86), .IN2(n68), .IN3(n87), .QN(n85) );
  AO21X1 U116 ( .IN1(row_sel_AQ2[1]), .IN2(n91), .IN3(n92), .Q(n145) );
  AO21X1 U117 ( .IN1(row_sel_AQ2[0]), .IN2(n91), .IN3(n93), .Q(n146) );
  AO21X1 U118 ( .IN1(done), .IN2(n68), .IN3(n76), .Q(n147) );
  AO21X1 U131 ( .IN1(row_sel_AQ_out[0]), .IN2(n91), .IN3(n93), .Q(n160) );
  AO222X1 U132 ( .IN1(n95), .IN2(col_sel_AQ_int[1]), .IN3(n96), .IN4(
        col_sel_AQ2_int[1]), .IN5(col_sel_R_int[1]), .IN6(n97), .Q(n161) );
  AO222X1 U133 ( .IN1(n95), .IN2(col_sel_AQ_int[0]), .IN3(n96), .IN4(
        col_sel_AQ2_int[0]), .IN5(col_sel_R_int[0]), .IN6(n97), .Q(n162) );
  AO22X1 U134 ( .IN1(n49), .IN2(col_sel_AQ_int[0]), .IN3(row_sel_R[0]), .IN4(
        n83), .Q(n163) );
  AO22X1 U135 ( .IN1(mult_counter[1]), .IN2(n98), .IN3(mult_counter[0]), .IN4(
        n78), .Q(n164) );
  AO22X1 U136 ( .IN1(n98), .IN2(mult_counter[0]), .IN3(n99), .IN4(n46), .Q(
        n165) );
  AO22X1 U137 ( .IN1(n49), .IN2(col_sel_AQ_int[1]), .IN3(row_sel_R[1]), .IN4(
        n83), .Q(n166) );
  AO21X1 U138 ( .IN1(in_b_vec_mult_sel), .IN2(n97), .IN3(n95), .Q(n167) );
  AO21X1 U139 ( .IN1(in_b_inner_prod_sel), .IN2(n100), .IN3(n59), .Q(n168) );
  NAND3X0 U140 ( .IN1(n103), .IN2(n100), .IN3(in_a_inner_prod_sel), .QN(n102)
         );
  NAND4X0 U141 ( .IN1(n104), .IN2(n56), .IN3(mult_counter[2]), .IN4(n105), 
        .QN(n100) );
  AO22X1 U142 ( .IN1(reduced_matrix), .IN2(n94), .IN3(red_mat_reg_out), .IN4(
        n107), .Q(n170) );
  AO21X1 U143 ( .IN1(col_sel_R_sel), .IN2(n68), .IN3(n94), .Q(n171) );
  AO21X1 U144 ( .IN1(col_sel_AQ2_sel), .IN2(n68), .IN3(n94), .Q(n172) );
  AO22X1 U145 ( .IN1(n48), .IN2(state[2]), .IN3(n108), .IN4(n109), .Q(n173) );
  OR4X1 U146 ( .IN1(n99), .IN2(n61), .IN3(n110), .IN4(n106), .Q(n108) );
  AO22X1 U147 ( .IN1(n48), .IN2(state[1]), .IN3(n111), .IN4(n109), .Q(n174) );
  AO22X1 U148 ( .IN1(n113), .IN2(col_sel_AQ_int[0]), .IN3(n114), .IN4(n56), 
        .Q(n175) );
  AO22X1 U149 ( .IN1(n113), .IN2(col_sel_AQ_int[1]), .IN3(n115), .IN4(n56), 
        .Q(n176) );
  AND2X1 U150 ( .IN1(n68), .IN2(n117), .Q(n113) );
  NAND3X0 U151 ( .IN1(n56), .IN2(mult_counter[2]), .IN3(n104), .QN(n117) );
  AO221X1 U152 ( .IN1(n118), .IN2(n119), .IN3(n52), .IN4(col_sel_AQ2_int[0]), 
        .IN5(n54), .Q(n177) );
  AO22X1 U153 ( .IN1(col_sel_AQ2_int[1]), .IN2(n121), .IN3(n122), .IN4(n90), 
        .Q(n178) );
  AO22X1 U154 ( .IN1(n116), .IN2(n119), .IN3(n110), .IN4(col_sel_AQ2_int[0]), 
        .Q(n122) );
  AO21X1 U155 ( .IN1(n104), .IN2(n56), .IN3(n89), .Q(n119) );
  XOR2X1 U156 ( .IN1(col_sel_AQ_int[1]), .IN2(col_sel_AQ_int[0]), .Q(n116) );
  NAND3X0 U157 ( .IN1(n90), .IN2(n40), .IN3(n110), .QN(n120) );
  AO21X1 U158 ( .IN1(mult_counter[2]), .IN2(n55), .IN3(n183), .Q(n90) );
  AO22X1 U159 ( .IN1(n98), .IN2(mult_counter[2]), .IN3(mult_counter[1]), .IN4(
        n78), .Q(n179) );
  AO22X1 U160 ( .IN1(n48), .IN2(state[3]), .IN3(n123), .IN4(n124), .Q(n180) );
  AO21X1 U161 ( .IN1(row_sel_AQ_out[1]), .IN2(n91), .IN3(n92), .Q(n181) );
  AND2X1 U162 ( .IN1(n125), .IN2(n60), .Q(n92) );
  XOR2X1 U163 ( .IN1(row_sel_AQ_out[1]), .IN2(row_sel_AQ_out[0]), .Q(n125) );
  AND3X1 U164 ( .IN1(n126), .IN2(n107), .IN3(n79), .Q(n91) );
  AO22X1 U165 ( .IN1(n48), .IN2(state[0]), .IN3(n128), .IN4(n109), .Q(n182) );
  NAND3X0 U166 ( .IN1(n112), .IN2(n68), .IN3(n127), .QN(n128) );
  AND2X1 U167 ( .IN1(col_sel_AQ_int[0]), .IN2(n105), .Q(n124) );
  OR2X1 U168 ( .IN1(red_mat_reg_out), .IN2(col_sel_AQ_int[1]), .Q(n105) );
  NAND3X0 U169 ( .IN1(n97), .IN2(n80), .IN3(n129), .QN(n109) );
  AOI221X1 U170 ( .IN1(done_inner_prod), .IN2(n84), .IN3(row_sel_AQ_out[0]), 
        .IN4(n130), .IN5(n94), .QN(n129) );
  NAND3X0 U171 ( .IN1(n65), .IN2(n64), .IN3(n131), .QN(n68) );
  NAND3X0 U172 ( .IN1(state[2]), .IN2(n65), .IN3(n132), .QN(n74) );
  AND3X1 U173 ( .IN1(n65), .IN2(n64), .IN3(n132), .Q(n81) );
  AND3X1 U174 ( .IN1(n131), .IN2(n64), .IN3(state[1]), .Q(n84) );
  AOI21X1 U175 ( .IN1(mult_counter[2]), .IN2(n78), .IN3(n76), .QN(n80) );
  AND4X1 U176 ( .IN1(state[3]), .IN2(n66), .IN3(n65), .IN4(n64), .Q(n76) );
  NAND3X0 U177 ( .IN1(state[2]), .IN2(state[1]), .IN3(n132), .QN(n67) );
  NAND3X0 U178 ( .IN1(n131), .IN2(n65), .IN3(state[2]), .QN(n71) );
  NAND3X0 U179 ( .IN1(state[1]), .IN2(n131), .IN3(state[2]), .QN(n72) );
  NAND3X0 U180 ( .IN1(state[1]), .IN2(n64), .IN3(n132), .QN(n86) );
  INVX0 U3 ( .INP(n97), .ZN(n47) );
  INVX0 U4 ( .INP(n127), .ZN(n55) );
  INVX0 U5 ( .INP(n82), .ZN(n45) );
  NOR2X0 U6 ( .IN1(n49), .IN2(n62), .QN(n97) );
  NOR2X0 U7 ( .IN1(n78), .IN2(n47), .QN(n98) );
  NOR2X0 U8 ( .IN1(n47), .IN2(n183), .QN(n82) );
  NOR2X0 U9 ( .IN1(n56), .IN2(n106), .QN(n127) );
  INVX0 U10 ( .INP(n79), .ZN(n60) );
  NOR2X0 U11 ( .IN1(n60), .IN2(n183), .QN(n101) );
  NOR2X0 U12 ( .IN1(n71), .IN2(n124), .QN(n106) );
  NOR2X0 U13 ( .IN1(n97), .IN2(n72), .QN(n96) );
  INVX0 U14 ( .INP(n109), .ZN(n48) );
  NOR2X0 U15 ( .IN1(n86), .IN2(n97), .QN(n95) );
  INVX0 U16 ( .INP(n73), .ZN(n62) );
  NOR2X0 U17 ( .IN1(n81), .IN2(n61), .QN(n79) );
  INVX0 U18 ( .INP(n68), .ZN(n183) );
  NAND2X0 U19 ( .IN1(n71), .IN2(n67), .QN(n78) );
  INVX0 U20 ( .INP(n67), .ZN(n56) );
  INVX0 U21 ( .INP(n72), .ZN(n63) );
  NOR2X0 U22 ( .IN1(n67), .IN2(n104), .QN(n110) );
  INVX0 U23 ( .INP(n74), .ZN(n61) );
  INVX0 U24 ( .INP(n71), .ZN(n89) );
  INVX0 U25 ( .INP(n107), .ZN(n94) );
  INVX0 U26 ( .INP(n86), .ZN(n50) );
  NAND2X0 U27 ( .IN1(n86), .IN2(n72), .QN(n99) );
  NOR2X0 U28 ( .IN1(n84), .IN2(n63), .QN(n112) );
  INVX0 U29 ( .INP(n83), .ZN(n49) );
  NOR2X0 U30 ( .IN1(col_sel_AQ_int[0]), .IN2(n113), .QN(n114) );
  INVX0 U31 ( .INP(n120), .ZN(n54) );
  NOR2X0 U32 ( .IN1(col_sel_AQ_int[0]), .IN2(n52), .QN(n118) );
  INVX0 U33 ( .INP(n90), .ZN(n52) );
  NOR2X0 U34 ( .IN1(n113), .IN2(n184), .QN(n115) );
  INVX0 U35 ( .INP(n116), .ZN(n184) );
  OA21X1 U36 ( .IN1(row_sel_AQ_out[1]), .IN2(red_mat_reg_out), .IN3(n60), .Q(
        n130) );
  NAND2X0 U37 ( .IN1(mult_counter[2]), .IN2(n55), .QN(n126) );
  NOR2X0 U38 ( .IN1(n79), .IN2(row_sel_AQ_out[0]), .QN(n93) );
  NAND2X0 U39 ( .IN1(done_inner_prod), .IN2(n63), .QN(n73) );
  NAND2X0 U40 ( .IN1(n101), .IN2(n102), .QN(n169) );
  NAND2X0 U41 ( .IN1(n106), .IN2(mult_counter[2]), .QN(n103) );
  NOR2X0 U42 ( .IN1(n48), .IN2(n71), .QN(n123) );
  NAND2X0 U43 ( .IN1(n112), .IN2(n79), .QN(n111) );
  INVX0 U44 ( .INP(n98), .ZN(n46) );
  NAND2X0 U45 ( .IN1(n90), .IN2(n120), .QN(n121) );
  OAI22X1 U46 ( .IN1(n39), .IN2(n53), .IN3(n41), .IN4(n88), .QN(n144) );
  NOR2X0 U47 ( .IN1(n78), .IN2(n94), .QN(n41) );
  NOR2X0 U48 ( .IN1(n90), .IN2(n60), .QN(n88) );
  INVX0 U49 ( .INP(n88), .ZN(n53) );
  INVX0 U50 ( .INP(n43), .ZN(n44) );
  INVX0 U51 ( .INP(rst), .ZN(n42) );
  NOR2X0 U52 ( .IN1(state[3]), .IN2(state[0]), .QN(n131) );
  NOR2X0 U53 ( .IN1(n66), .IN2(state[3]), .QN(n132) );
  NAND2X0 U54 ( .IN1(start), .IN2(n183), .QN(n107) );
  OA21X1 U55 ( .IN1(red_mat_reg_out), .IN2(col_sel_AQ2_int[1]), .IN3(
        col_sel_AQ2_int[0]), .Q(n104) );
  NAND2X0 U56 ( .IN1(done_inv_sqrt), .IN2(n50), .QN(n83) );
  NAND2X0 U57 ( .IN1(n71), .IN2(n72), .QN(n69) );
  INVX0 U58 ( .INP(n70), .ZN(n58) );
  INVX0 U59 ( .INP(n85), .ZN(n51) );
  NAND2X0 U60 ( .IN1(n84), .IN2(done_inner_prod), .QN(n87) );
  INVX0 U61 ( .INP(n77), .ZN(n57) );
  NAND2X0 U62 ( .IN1(n79), .IN2(n80), .QN(n77) );
  INVX0 U63 ( .INP(n101), .ZN(n59) );
  INVX0 U64 ( .INP(rst), .ZN(n1) );
  INVX0 U65 ( .INP(rst), .ZN(n2) );
  INVX0 U66 ( .INP(rst), .ZN(n3) );
  INVX0 U67 ( .INP(rst), .ZN(n4) );
  INVX0 U68 ( .INP(rst), .ZN(n5) );
  INVX0 U69 ( .INP(rst), .ZN(n6) );
  INVX0 U70 ( .INP(rst), .ZN(n7) );
  INVX0 U71 ( .INP(rst), .ZN(n8) );
  INVX0 U72 ( .INP(rst), .ZN(n9) );
  INVX0 U73 ( .INP(rst), .ZN(n10) );
  INVX0 U74 ( .INP(rst), .ZN(n11) );
  INVX0 U75 ( .INP(rst), .ZN(n12) );
  INVX0 U76 ( .INP(rst), .ZN(n14) );
  INVX0 U77 ( .INP(rst), .ZN(n15) );
  INVX0 U78 ( .INP(rst), .ZN(n16) );
  INVX0 U79 ( .INP(rst), .ZN(n17) );
  INVX0 U80 ( .INP(rst), .ZN(n18) );
  INVX0 U81 ( .INP(rst), .ZN(n19) );
  INVX0 U82 ( .INP(rst), .ZN(n22) );
  INVX0 U83 ( .INP(rst), .ZN(n23) );
  INVX0 U84 ( .INP(rst), .ZN(n24) );
  INVX0 U85 ( .INP(rst), .ZN(n25) );
  INVX0 U86 ( .INP(rst), .ZN(n26) );
  INVX0 U87 ( .INP(rst), .ZN(n27) );
  INVX0 U88 ( .INP(rst), .ZN(n28) );
  INVX0 U89 ( .INP(rst), .ZN(n29) );
  INVX0 U90 ( .INP(rst), .ZN(n30) );
  INVX0 U91 ( .INP(rst), .ZN(n31) );
  INVX0 U92 ( .INP(rst), .ZN(n32) );
  INVX0 U93 ( .INP(rst), .ZN(n33) );
  INVX0 U94 ( .INP(rst), .ZN(n34) );
  INVX0 U95 ( .INP(rst), .ZN(n35) );
  INVX0 U96 ( .INP(rst), .ZN(n36) );
  INVX0 U97 ( .INP(rst), .ZN(n37) );
  INVX0 U98 ( .INP(rst), .ZN(n38) );
  INVX0 U99 ( .INP(rst), .ZN(n13) );
  INVX0 U114 ( .INP(rst), .ZN(n20) );
  INVX0 U115 ( .INP(rst), .ZN(n21) );
  NAND2X1 U119 ( .IN1(n42), .IN2(n89), .QN(n43) );
  MUX21X1 U120 ( .IN1(in_a_r_mult[0]), .IN2(out_inv_sqrt[0]), .S(n44), .Q(n159) );
  MUX21X1 U121 ( .IN1(in_a_r_mult[1]), .IN2(out_inv_sqrt[1]), .S(n44), .Q(n158) );
  MUX21X1 U122 ( .IN1(in_a_r_mult[2]), .IN2(out_inv_sqrt[2]), .S(n44), .Q(n157) );
  MUX21X1 U123 ( .IN1(in_a_r_mult[3]), .IN2(out_inv_sqrt[3]), .S(n44), .Q(n156) );
  MUX21X1 U124 ( .IN1(in_a_r_mult[4]), .IN2(out_inv_sqrt[4]), .S(n44), .Q(n155) );
  MUX21X1 U125 ( .IN1(in_a_r_mult[5]), .IN2(out_inv_sqrt[5]), .S(n44), .Q(n154) );
  MUX21X1 U126 ( .IN1(in_a_r_mult[6]), .IN2(out_inv_sqrt[6]), .S(n44), .Q(n153) );
  MUX21X1 U127 ( .IN1(in_a_r_mult[7]), .IN2(out_inv_sqrt[7]), .S(n44), .Q(n152) );
  MUX21X1 U128 ( .IN1(in_a_r_mult[8]), .IN2(out_inv_sqrt[8]), .S(n44), .Q(n151) );
  MUX21X1 U129 ( .IN1(in_a_r_mult[9]), .IN2(out_inv_sqrt[9]), .S(n44), .Q(n150) );
  MUX21X1 U130 ( .IN1(in_a_r_mult[10]), .IN2(out_inv_sqrt[10]), .S(n44), .Q(
        n149) );
  MUX21X1 U181 ( .IN1(in_a_r_mult[11]), .IN2(out_inv_sqrt[11]), .S(n44), .Q(
        n148) );
endmodule


module qr_decomp_USE_NEWTON1 ( .in_A_r({\in_A_r[0][11] , \in_A_r[0][10] , 
        \in_A_r[0][9] , \in_A_r[0][8] , \in_A_r[0][7] , \in_A_r[0][6] , 
        \in_A_r[0][5] , \in_A_r[0][4] , \in_A_r[0][3] , \in_A_r[0][2] , 
        \in_A_r[0][1] , \in_A_r[0][0] , \in_A_r[1][11] , \in_A_r[1][10] , 
        \in_A_r[1][9] , \in_A_r[1][8] , \in_A_r[1][7] , \in_A_r[1][6] , 
        \in_A_r[1][5] , \in_A_r[1][4] , \in_A_r[1][3] , \in_A_r[1][2] , 
        \in_A_r[1][1] , \in_A_r[1][0] , \in_A_r[2][11] , \in_A_r[2][10] , 
        \in_A_r[2][9] , \in_A_r[2][8] , \in_A_r[2][7] , \in_A_r[2][6] , 
        \in_A_r[2][5] , \in_A_r[2][4] , \in_A_r[2][3] , \in_A_r[2][2] , 
        \in_A_r[2][1] , \in_A_r[2][0] , \in_A_r[3][11] , \in_A_r[3][10] , 
        \in_A_r[3][9] , \in_A_r[3][8] , \in_A_r[3][7] , \in_A_r[3][6] , 
        \in_A_r[3][5] , \in_A_r[3][4] , \in_A_r[3][3] , \in_A_r[3][2] , 
        \in_A_r[3][1] , \in_A_r[3][0] }), .in_A_i({\in_A_i[0][11] , 
        \in_A_i[0][10] , \in_A_i[0][9] , \in_A_i[0][8] , \in_A_i[0][7] , 
        \in_A_i[0][6] , \in_A_i[0][5] , \in_A_i[0][4] , \in_A_i[0][3] , 
        \in_A_i[0][2] , \in_A_i[0][1] , \in_A_i[0][0] , \in_A_i[1][11] , 
        \in_A_i[1][10] , \in_A_i[1][9] , \in_A_i[1][8] , \in_A_i[1][7] , 
        \in_A_i[1][6] , \in_A_i[1][5] , \in_A_i[1][4] , \in_A_i[1][3] , 
        \in_A_i[1][2] , \in_A_i[1][1] , \in_A_i[1][0] , \in_A_i[2][11] , 
        \in_A_i[2][10] , \in_A_i[2][9] , \in_A_i[2][8] , \in_A_i[2][7] , 
        \in_A_i[2][6] , \in_A_i[2][5] , \in_A_i[2][4] , \in_A_i[2][3] , 
        \in_A_i[2][2] , \in_A_i[2][1] , \in_A_i[2][0] , \in_A_i[3][11] , 
        \in_A_i[3][10] , \in_A_i[3][9] , \in_A_i[3][8] , \in_A_i[3][7] , 
        \in_A_i[3][6] , \in_A_i[3][5] , \in_A_i[3][4] , \in_A_i[3][3] , 
        \in_A_i[3][2] , \in_A_i[3][1] , \in_A_i[3][0] }), .out_Q_r({
        \out_Q_r[0][11] , \out_Q_r[0][10] , \out_Q_r[0][9] , \out_Q_r[0][8] , 
        \out_Q_r[0][7] , \out_Q_r[0][6] , \out_Q_r[0][5] , \out_Q_r[0][4] , 
        \out_Q_r[0][3] , \out_Q_r[0][2] , \out_Q_r[0][1] , \out_Q_r[0][0] , 
        \out_Q_r[1][11] , \out_Q_r[1][10] , \out_Q_r[1][9] , \out_Q_r[1][8] , 
        \out_Q_r[1][7] , \out_Q_r[1][6] , \out_Q_r[1][5] , \out_Q_r[1][4] , 
        \out_Q_r[1][3] , \out_Q_r[1][2] , \out_Q_r[1][1] , \out_Q_r[1][0] , 
        \out_Q_r[2][11] , \out_Q_r[2][10] , \out_Q_r[2][9] , \out_Q_r[2][8] , 
        \out_Q_r[2][7] , \out_Q_r[2][6] , \out_Q_r[2][5] , \out_Q_r[2][4] , 
        \out_Q_r[2][3] , \out_Q_r[2][2] , \out_Q_r[2][1] , \out_Q_r[2][0] , 
        \out_Q_r[3][11] , \out_Q_r[3][10] , \out_Q_r[3][9] , \out_Q_r[3][8] , 
        \out_Q_r[3][7] , \out_Q_r[3][6] , \out_Q_r[3][5] , \out_Q_r[3][4] , 
        \out_Q_r[3][3] , \out_Q_r[3][2] , \out_Q_r[3][1] , \out_Q_r[3][0] }), 
    .out_Q_i({\out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] , 
        \out_Q_i[0][8] , \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] , 
        \out_Q_i[0][4] , \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] , 
        \out_Q_i[0][0] , \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] , 
        \out_Q_i[1][8] , \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] , 
        \out_Q_i[1][4] , \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] , 
        \out_Q_i[1][0] , \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] , 
        \out_Q_i[2][8] , \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] , 
        \out_Q_i[2][4] , \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] , 
        \out_Q_i[2][0] , \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] , 
        \out_Q_i[3][8] , \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] , 
        \out_Q_i[3][4] , \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] , 
        \out_Q_i[3][0] }), .out_R_r({\out_R_r[0][11] , \out_R_r[0][10] , 
        \out_R_r[0][9] , \out_R_r[0][8] , \out_R_r[0][7] , \out_R_r[0][6] , 
        \out_R_r[0][5] , \out_R_r[0][4] , \out_R_r[0][3] , \out_R_r[0][2] , 
        \out_R_r[0][1] , \out_R_r[0][0] , \out_R_r[1][11] , \out_R_r[1][10] , 
        \out_R_r[1][9] , \out_R_r[1][8] , \out_R_r[1][7] , \out_R_r[1][6] , 
        \out_R_r[1][5] , \out_R_r[1][4] , \out_R_r[1][3] , \out_R_r[1][2] , 
        \out_R_r[1][1] , \out_R_r[1][0] , \out_R_r[2][11] , \out_R_r[2][10] , 
        \out_R_r[2][9] , \out_R_r[2][8] , \out_R_r[2][7] , \out_R_r[2][6] , 
        \out_R_r[2][5] , \out_R_r[2][4] , \out_R_r[2][3] , \out_R_r[2][2] , 
        \out_R_r[2][1] , \out_R_r[2][0] , \out_R_r[3][11] , \out_R_r[3][10] , 
        \out_R_r[3][9] , \out_R_r[3][8] , \out_R_r[3][7] , \out_R_r[3][6] , 
        \out_R_r[3][5] , \out_R_r[3][4] , \out_R_r[3][3] , \out_R_r[3][2] , 
        \out_R_r[3][1] , \out_R_r[3][0] }), .out_R_i({\out_R_i[0][11] , 
        \out_R_i[0][10] , \out_R_i[0][9] , \out_R_i[0][8] , \out_R_i[0][7] , 
        \out_R_i[0][6] , \out_R_i[0][5] , \out_R_i[0][4] , \out_R_i[0][3] , 
        \out_R_i[0][2] , \out_R_i[0][1] , \out_R_i[0][0] , \out_R_i[1][11] , 
        \out_R_i[1][10] , \out_R_i[1][9] , \out_R_i[1][8] , \out_R_i[1][7] , 
        \out_R_i[1][6] , \out_R_i[1][5] , \out_R_i[1][4] , \out_R_i[1][3] , 
        \out_R_i[1][2] , \out_R_i[1][1] , \out_R_i[1][0] , \out_R_i[2][11] , 
        \out_R_i[2][10] , \out_R_i[2][9] , \out_R_i[2][8] , \out_R_i[2][7] , 
        \out_R_i[2][6] , \out_R_i[2][5] , \out_R_i[2][4] , \out_R_i[2][3] , 
        \out_R_i[2][2] , \out_R_i[2][1] , \out_R_i[2][0] , \out_R_i[3][11] , 
        \out_R_i[3][10] , \out_R_i[3][9] , \out_R_i[3][8] , \out_R_i[3][7] , 
        \out_R_i[3][6] , \out_R_i[3][5] , \out_R_i[3][4] , \out_R_i[3][3] , 
        \out_R_i[3][2] , \out_R_i[3][1] , \out_R_i[3][0] }), wr_A, col_sel_AQ, 
        col_sel_R, reduced_matrix, clk, rst, start, done );
  input [1:0] col_sel_AQ;
  input [1:0] col_sel_R;
  input \in_A_r[0][11] , \in_A_r[0][10] , \in_A_r[0][9] , \in_A_r[0][8] ,
         \in_A_r[0][7] , \in_A_r[0][6] , \in_A_r[0][5] , \in_A_r[0][4] ,
         \in_A_r[0][3] , \in_A_r[0][2] , \in_A_r[0][1] , \in_A_r[0][0] ,
         \in_A_r[1][11] , \in_A_r[1][10] , \in_A_r[1][9] , \in_A_r[1][8] ,
         \in_A_r[1][7] , \in_A_r[1][6] , \in_A_r[1][5] , \in_A_r[1][4] ,
         \in_A_r[1][3] , \in_A_r[1][2] , \in_A_r[1][1] , \in_A_r[1][0] ,
         \in_A_r[2][11] , \in_A_r[2][10] , \in_A_r[2][9] , \in_A_r[2][8] ,
         \in_A_r[2][7] , \in_A_r[2][6] , \in_A_r[2][5] , \in_A_r[2][4] ,
         \in_A_r[2][3] , \in_A_r[2][2] , \in_A_r[2][1] , \in_A_r[2][0] ,
         \in_A_r[3][11] , \in_A_r[3][10] , \in_A_r[3][9] , \in_A_r[3][8] ,
         \in_A_r[3][7] , \in_A_r[3][6] , \in_A_r[3][5] , \in_A_r[3][4] ,
         \in_A_r[3][3] , \in_A_r[3][2] , \in_A_r[3][1] , \in_A_r[3][0] ,
         \in_A_i[0][11] , \in_A_i[0][10] , \in_A_i[0][9] , \in_A_i[0][8] ,
         \in_A_i[0][7] , \in_A_i[0][6] , \in_A_i[0][5] , \in_A_i[0][4] ,
         \in_A_i[0][3] , \in_A_i[0][2] , \in_A_i[0][1] , \in_A_i[0][0] ,
         \in_A_i[1][11] , \in_A_i[1][10] , \in_A_i[1][9] , \in_A_i[1][8] ,
         \in_A_i[1][7] , \in_A_i[1][6] , \in_A_i[1][5] , \in_A_i[1][4] ,
         \in_A_i[1][3] , \in_A_i[1][2] , \in_A_i[1][1] , \in_A_i[1][0] ,
         \in_A_i[2][11] , \in_A_i[2][10] , \in_A_i[2][9] , \in_A_i[2][8] ,
         \in_A_i[2][7] , \in_A_i[2][6] , \in_A_i[2][5] , \in_A_i[2][4] ,
         \in_A_i[2][3] , \in_A_i[2][2] , \in_A_i[2][1] , \in_A_i[2][0] ,
         \in_A_i[3][11] , \in_A_i[3][10] , \in_A_i[3][9] , \in_A_i[3][8] ,
         \in_A_i[3][7] , \in_A_i[3][6] , \in_A_i[3][5] , \in_A_i[3][4] ,
         \in_A_i[3][3] , \in_A_i[3][2] , \in_A_i[3][1] , \in_A_i[3][0] , wr_A,
         reduced_matrix, clk, rst, start;
  output \out_Q_r[0][11] , \out_Q_r[0][10] , \out_Q_r[0][9] , \out_Q_r[0][8] ,
         \out_Q_r[0][7] , \out_Q_r[0][6] , \out_Q_r[0][5] , \out_Q_r[0][4] ,
         \out_Q_r[0][3] , \out_Q_r[0][2] , \out_Q_r[0][1] , \out_Q_r[0][0] ,
         \out_Q_r[1][11] , \out_Q_r[1][10] , \out_Q_r[1][9] , \out_Q_r[1][8] ,
         \out_Q_r[1][7] , \out_Q_r[1][6] , \out_Q_r[1][5] , \out_Q_r[1][4] ,
         \out_Q_r[1][3] , \out_Q_r[1][2] , \out_Q_r[1][1] , \out_Q_r[1][0] ,
         \out_Q_r[2][11] , \out_Q_r[2][10] , \out_Q_r[2][9] , \out_Q_r[2][8] ,
         \out_Q_r[2][7] , \out_Q_r[2][6] , \out_Q_r[2][5] , \out_Q_r[2][4] ,
         \out_Q_r[2][3] , \out_Q_r[2][2] , \out_Q_r[2][1] , \out_Q_r[2][0] ,
         \out_Q_r[3][11] , \out_Q_r[3][10] , \out_Q_r[3][9] , \out_Q_r[3][8] ,
         \out_Q_r[3][7] , \out_Q_r[3][6] , \out_Q_r[3][5] , \out_Q_r[3][4] ,
         \out_Q_r[3][3] , \out_Q_r[3][2] , \out_Q_r[3][1] , \out_Q_r[3][0] ,
         \out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] , \out_Q_i[0][8] ,
         \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] , \out_Q_i[0][4] ,
         \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] , \out_Q_i[0][0] ,
         \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] , \out_Q_i[1][8] ,
         \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] , \out_Q_i[1][4] ,
         \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] , \out_Q_i[1][0] ,
         \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] , \out_Q_i[2][8] ,
         \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] , \out_Q_i[2][4] ,
         \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] , \out_Q_i[2][0] ,
         \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] , \out_Q_i[3][8] ,
         \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] , \out_Q_i[3][4] ,
         \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] , \out_Q_i[3][0] ,
         \out_R_r[0][11] , \out_R_r[0][10] , \out_R_r[0][9] , \out_R_r[0][8] ,
         \out_R_r[0][7] , \out_R_r[0][6] , \out_R_r[0][5] , \out_R_r[0][4] ,
         \out_R_r[0][3] , \out_R_r[0][2] , \out_R_r[0][1] , \out_R_r[0][0] ,
         \out_R_r[1][11] , \out_R_r[1][10] , \out_R_r[1][9] , \out_R_r[1][8] ,
         \out_R_r[1][7] , \out_R_r[1][6] , \out_R_r[1][5] , \out_R_r[1][4] ,
         \out_R_r[1][3] , \out_R_r[1][2] , \out_R_r[1][1] , \out_R_r[1][0] ,
         \out_R_r[2][11] , \out_R_r[2][10] , \out_R_r[2][9] , \out_R_r[2][8] ,
         \out_R_r[2][7] , \out_R_r[2][6] , \out_R_r[2][5] , \out_R_r[2][4] ,
         \out_R_r[2][3] , \out_R_r[2][2] , \out_R_r[2][1] , \out_R_r[2][0] ,
         \out_R_r[3][11] , \out_R_r[3][10] , \out_R_r[3][9] , \out_R_r[3][8] ,
         \out_R_r[3][7] , \out_R_r[3][6] , \out_R_r[3][5] , \out_R_r[3][4] ,
         \out_R_r[3][3] , \out_R_r[3][2] , \out_R_r[3][1] , \out_R_r[3][0] ,
         \out_R_i[0][11] , \out_R_i[0][10] , \out_R_i[0][9] , \out_R_i[0][8] ,
         \out_R_i[0][7] , \out_R_i[0][6] , \out_R_i[0][5] , \out_R_i[0][4] ,
         \out_R_i[0][3] , \out_R_i[0][2] , \out_R_i[0][1] , \out_R_i[0][0] ,
         \out_R_i[1][11] , \out_R_i[1][10] , \out_R_i[1][9] , \out_R_i[1][8] ,
         \out_R_i[1][7] , \out_R_i[1][6] , \out_R_i[1][5] , \out_R_i[1][4] ,
         \out_R_i[1][3] , \out_R_i[1][2] , \out_R_i[1][1] , \out_R_i[1][0] ,
         \out_R_i[2][11] , \out_R_i[2][10] , \out_R_i[2][9] , \out_R_i[2][8] ,
         \out_R_i[2][7] , \out_R_i[2][6] , \out_R_i[2][5] , \out_R_i[2][4] ,
         \out_R_i[2][3] , \out_R_i[2][2] , \out_R_i[2][1] , \out_R_i[2][0] ,
         \out_R_i[3][11] , \out_R_i[3][10] , \out_R_i[3][9] , \out_R_i[3][8] ,
         \out_R_i[3][7] , \out_R_i[3][6] , \out_R_i[3][5] , \out_R_i[3][4] ,
         \out_R_i[3][3] , \out_R_i[3][2] , \out_R_i[3][1] , \out_R_i[3][0] ,
         done;
  wire   \vec_in_r_AQ_mux[0][11] , \vec_in_r_AQ_mux[0][10] ,
         \vec_in_r_AQ_mux[0][9] , \vec_in_r_AQ_mux[0][8] ,
         \vec_in_r_AQ_mux[0][7] , \vec_in_r_AQ_mux[0][6] ,
         \vec_in_r_AQ_mux[0][5] , \vec_in_r_AQ_mux[0][4] ,
         \vec_in_r_AQ_mux[0][3] , \vec_in_r_AQ_mux[0][2] ,
         \vec_in_r_AQ_mux[0][1] , \vec_in_r_AQ_mux[0][0] ,
         \vec_in_r_AQ_mux[1][11] , \vec_in_r_AQ_mux[1][10] ,
         \vec_in_r_AQ_mux[1][9] , \vec_in_r_AQ_mux[1][8] ,
         \vec_in_r_AQ_mux[1][7] , \vec_in_r_AQ_mux[1][6] ,
         \vec_in_r_AQ_mux[1][5] , \vec_in_r_AQ_mux[1][4] ,
         \vec_in_r_AQ_mux[1][3] , \vec_in_r_AQ_mux[1][2] ,
         \vec_in_r_AQ_mux[1][1] , \vec_in_r_AQ_mux[1][0] ,
         \vec_in_r_AQ_mux[2][11] , \vec_in_r_AQ_mux[2][10] ,
         \vec_in_r_AQ_mux[2][9] , \vec_in_r_AQ_mux[2][8] ,
         \vec_in_r_AQ_mux[2][7] , \vec_in_r_AQ_mux[2][6] ,
         \vec_in_r_AQ_mux[2][5] , \vec_in_r_AQ_mux[2][4] ,
         \vec_in_r_AQ_mux[2][3] , \vec_in_r_AQ_mux[2][2] ,
         \vec_in_r_AQ_mux[2][1] , \vec_in_r_AQ_mux[2][0] ,
         \vec_in_r_AQ_mux[3][11] , \vec_in_r_AQ_mux[3][10] ,
         \vec_in_r_AQ_mux[3][9] , \vec_in_r_AQ_mux[3][8] ,
         \vec_in_r_AQ_mux[3][7] , \vec_in_r_AQ_mux[3][6] ,
         \vec_in_r_AQ_mux[3][5] , \vec_in_r_AQ_mux[3][4] ,
         \vec_in_r_AQ_mux[3][3] , \vec_in_r_AQ_mux[3][2] ,
         \vec_in_r_AQ_mux[3][1] , \vec_in_r_AQ_mux[3][0] ,
         \vec_in_i_AQ_mux[0][11] , \vec_in_i_AQ_mux[0][10] ,
         \vec_in_i_AQ_mux[0][9] , \vec_in_i_AQ_mux[0][8] ,
         \vec_in_i_AQ_mux[0][7] , \vec_in_i_AQ_mux[0][6] ,
         \vec_in_i_AQ_mux[0][5] , \vec_in_i_AQ_mux[0][4] ,
         \vec_in_i_AQ_mux[0][3] , \vec_in_i_AQ_mux[0][2] ,
         \vec_in_i_AQ_mux[0][1] , \vec_in_i_AQ_mux[0][0] ,
         \vec_in_i_AQ_mux[1][11] , \vec_in_i_AQ_mux[1][10] ,
         \vec_in_i_AQ_mux[1][9] , \vec_in_i_AQ_mux[1][8] ,
         \vec_in_i_AQ_mux[1][7] , \vec_in_i_AQ_mux[1][6] ,
         \vec_in_i_AQ_mux[1][5] , \vec_in_i_AQ_mux[1][4] ,
         \vec_in_i_AQ_mux[1][3] , \vec_in_i_AQ_mux[1][2] ,
         \vec_in_i_AQ_mux[1][1] , \vec_in_i_AQ_mux[1][0] ,
         \vec_in_i_AQ_mux[2][11] , \vec_in_i_AQ_mux[2][10] ,
         \vec_in_i_AQ_mux[2][9] , \vec_in_i_AQ_mux[2][8] ,
         \vec_in_i_AQ_mux[2][7] , \vec_in_i_AQ_mux[2][6] ,
         \vec_in_i_AQ_mux[2][5] , \vec_in_i_AQ_mux[2][4] ,
         \vec_in_i_AQ_mux[2][3] , \vec_in_i_AQ_mux[2][2] ,
         \vec_in_i_AQ_mux[2][1] , \vec_in_i_AQ_mux[2][0] ,
         \vec_in_i_AQ_mux[3][11] , \vec_in_i_AQ_mux[3][10] ,
         \vec_in_i_AQ_mux[3][9] , \vec_in_i_AQ_mux[3][8] ,
         \vec_in_i_AQ_mux[3][7] , \vec_in_i_AQ_mux[3][6] ,
         \vec_in_i_AQ_mux[3][5] , \vec_in_i_AQ_mux[3][4] ,
         \vec_in_i_AQ_mux[3][3] , \vec_in_i_AQ_mux[3][2] ,
         \vec_in_i_AQ_mux[3][1] , \vec_in_i_AQ_mux[3][0] ,
         \vec_out_r_AQ[0][11] , \vec_out_r_AQ[0][10] , \vec_out_r_AQ[0][9] ,
         \vec_out_r_AQ[0][8] , \vec_out_r_AQ[0][7] , \vec_out_r_AQ[0][6] ,
         \vec_out_r_AQ[0][5] , \vec_out_r_AQ[0][4] , \vec_out_r_AQ[0][3] ,
         \vec_out_r_AQ[0][2] , \vec_out_r_AQ[0][1] , \vec_out_r_AQ[0][0] ,
         \vec_out_r_AQ[1][11] , \vec_out_r_AQ[1][10] , \vec_out_r_AQ[1][9] ,
         \vec_out_r_AQ[1][8] , \vec_out_r_AQ[1][7] , \vec_out_r_AQ[1][6] ,
         \vec_out_r_AQ[1][5] , \vec_out_r_AQ[1][4] , \vec_out_r_AQ[1][3] ,
         \vec_out_r_AQ[1][2] , \vec_out_r_AQ[1][1] , \vec_out_r_AQ[1][0] ,
         \vec_out_r_AQ[2][11] , \vec_out_r_AQ[2][10] , \vec_out_r_AQ[2][9] ,
         \vec_out_r_AQ[2][8] , \vec_out_r_AQ[2][7] , \vec_out_r_AQ[2][6] ,
         \vec_out_r_AQ[2][5] , \vec_out_r_AQ[2][4] , \vec_out_r_AQ[2][3] ,
         \vec_out_r_AQ[2][2] , \vec_out_r_AQ[2][1] , \vec_out_r_AQ[2][0] ,
         \vec_out_r_AQ[3][11] , \vec_out_r_AQ[3][10] , \vec_out_r_AQ[3][9] ,
         \vec_out_r_AQ[3][8] , \vec_out_r_AQ[3][7] , \vec_out_r_AQ[3][6] ,
         \vec_out_r_AQ[3][5] , \vec_out_r_AQ[3][4] , \vec_out_r_AQ[3][3] ,
         \vec_out_r_AQ[3][2] , \vec_out_r_AQ[3][1] , \vec_out_r_AQ[3][0] ,
         \vec_out_i_AQ[0][11] , \vec_out_i_AQ[0][10] , \vec_out_i_AQ[0][9] ,
         \vec_out_i_AQ[0][8] , \vec_out_i_AQ[0][7] , \vec_out_i_AQ[0][6] ,
         \vec_out_i_AQ[0][5] , \vec_out_i_AQ[0][4] , \vec_out_i_AQ[0][3] ,
         \vec_out_i_AQ[0][2] , \vec_out_i_AQ[0][1] , \vec_out_i_AQ[0][0] ,
         \vec_out_i_AQ[1][11] , \vec_out_i_AQ[1][10] , \vec_out_i_AQ[1][9] ,
         \vec_out_i_AQ[1][8] , \vec_out_i_AQ[1][7] , \vec_out_i_AQ[1][6] ,
         \vec_out_i_AQ[1][5] , \vec_out_i_AQ[1][4] , \vec_out_i_AQ[1][3] ,
         \vec_out_i_AQ[1][2] , \vec_out_i_AQ[1][1] , \vec_out_i_AQ[1][0] ,
         \vec_out_i_AQ[2][11] , \vec_out_i_AQ[2][10] , \vec_out_i_AQ[2][9] ,
         \vec_out_i_AQ[2][8] , \vec_out_i_AQ[2][7] , \vec_out_i_AQ[2][6] ,
         \vec_out_i_AQ[2][5] , \vec_out_i_AQ[2][4] , \vec_out_i_AQ[2][3] ,
         \vec_out_i_AQ[2][2] , \vec_out_i_AQ[2][1] , \vec_out_i_AQ[2][0] ,
         \vec_out_i_AQ[3][11] , \vec_out_i_AQ[3][10] , \vec_out_i_AQ[3][9] ,
         \vec_out_i_AQ[3][8] , \vec_out_i_AQ[3][7] , \vec_out_i_AQ[3][6] ,
         \vec_out_i_AQ[3][5] , \vec_out_i_AQ[3][4] , \vec_out_i_AQ[3][3] ,
         \vec_out_i_AQ[3][2] , \vec_out_i_AQ[3][1] , \vec_out_i_AQ[3][0] ,
         wr_en_AQ_mux, wr_en_R, red_mat_reg, start_inner_prod, done_inner_prod,
         \out_r_vec_mult[0][11] , \out_r_vec_mult[0][10] ,
         \out_r_vec_mult[0][9] , \out_r_vec_mult[0][8] ,
         \out_r_vec_mult[0][7] , \out_r_vec_mult[0][6] ,
         \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] ,
         \out_r_vec_mult[0][3] , \out_r_vec_mult[0][2] ,
         \out_r_vec_mult[0][1] , \out_r_vec_mult[0][0] ,
         \out_r_vec_mult[1][11] , \out_r_vec_mult[1][10] ,
         \out_r_vec_mult[1][9] , \out_r_vec_mult[1][8] ,
         \out_r_vec_mult[1][7] , \out_r_vec_mult[1][6] ,
         \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] ,
         \out_r_vec_mult[1][3] , \out_r_vec_mult[1][2] ,
         \out_r_vec_mult[1][1] , \out_r_vec_mult[1][0] ,
         \out_r_vec_mult[2][11] , \out_r_vec_mult[2][10] ,
         \out_r_vec_mult[2][9] , \out_r_vec_mult[2][8] ,
         \out_r_vec_mult[2][7] , \out_r_vec_mult[2][6] ,
         \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] ,
         \out_r_vec_mult[2][3] , \out_r_vec_mult[2][2] ,
         \out_r_vec_mult[2][1] , \out_r_vec_mult[2][0] ,
         \out_r_vec_mult[3][11] , \out_r_vec_mult[3][10] ,
         \out_r_vec_mult[3][9] , \out_r_vec_mult[3][8] ,
         \out_r_vec_mult[3][7] , \out_r_vec_mult[3][6] ,
         \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] ,
         \out_r_vec_mult[3][3] , \out_r_vec_mult[3][2] ,
         \out_r_vec_mult[3][1] , \out_r_vec_mult[3][0] ,
         \out_i_vec_mult[0][11] , \out_i_vec_mult[0][10] ,
         \out_i_vec_mult[0][9] , \out_i_vec_mult[0][8] ,
         \out_i_vec_mult[0][7] , \out_i_vec_mult[0][6] ,
         \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] ,
         \out_i_vec_mult[0][3] , \out_i_vec_mult[0][2] ,
         \out_i_vec_mult[0][1] , \out_i_vec_mult[0][0] ,
         \out_i_vec_mult[1][11] , \out_i_vec_mult[1][10] ,
         \out_i_vec_mult[1][9] , \out_i_vec_mult[1][8] ,
         \out_i_vec_mult[1][7] , \out_i_vec_mult[1][6] ,
         \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] ,
         \out_i_vec_mult[1][3] , \out_i_vec_mult[1][2] ,
         \out_i_vec_mult[1][1] , \out_i_vec_mult[1][0] ,
         \out_i_vec_mult[2][11] , \out_i_vec_mult[2][10] ,
         \out_i_vec_mult[2][9] , \out_i_vec_mult[2][8] ,
         \out_i_vec_mult[2][7] , \out_i_vec_mult[2][6] ,
         \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] ,
         \out_i_vec_mult[2][3] , \out_i_vec_mult[2][2] ,
         \out_i_vec_mult[2][1] , \out_i_vec_mult[2][0] ,
         \out_i_vec_mult[3][11] , \out_i_vec_mult[3][10] ,
         \out_i_vec_mult[3][9] , \out_i_vec_mult[3][8] ,
         \out_i_vec_mult[3][7] , \out_i_vec_mult[3][6] ,
         \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] ,
         \out_i_vec_mult[3][3] , \out_i_vec_mult[3][2] ,
         \out_i_vec_mult[3][1] , \out_i_vec_mult[3][0] ,
         \out_r_vec_sub[0][11] , \out_r_vec_sub[0][10] , \out_r_vec_sub[0][9] ,
         \out_r_vec_sub[0][8] , \out_r_vec_sub[0][7] , \out_r_vec_sub[0][6] ,
         \out_r_vec_sub[0][5] , \out_r_vec_sub[0][4] , \out_r_vec_sub[0][3] ,
         \out_r_vec_sub[0][2] , \out_r_vec_sub[0][1] , \out_r_vec_sub[0][0] ,
         \out_r_vec_sub[1][11] , \out_r_vec_sub[1][10] , \out_r_vec_sub[1][9] ,
         \out_r_vec_sub[1][8] , \out_r_vec_sub[1][7] , \out_r_vec_sub[1][6] ,
         \out_r_vec_sub[1][5] , \out_r_vec_sub[1][4] , \out_r_vec_sub[1][3] ,
         \out_r_vec_sub[1][2] , \out_r_vec_sub[1][1] , \out_r_vec_sub[1][0] ,
         \out_r_vec_sub[2][11] , \out_r_vec_sub[2][10] , \out_r_vec_sub[2][9] ,
         \out_r_vec_sub[2][8] , \out_r_vec_sub[2][7] , \out_r_vec_sub[2][6] ,
         \out_r_vec_sub[2][5] , \out_r_vec_sub[2][4] , \out_r_vec_sub[2][3] ,
         \out_r_vec_sub[2][2] , \out_r_vec_sub[2][1] , \out_r_vec_sub[2][0] ,
         \out_r_vec_sub[3][11] , \out_r_vec_sub[3][10] , \out_r_vec_sub[3][9] ,
         \out_r_vec_sub[3][8] , \out_r_vec_sub[3][7] , \out_r_vec_sub[3][6] ,
         \out_r_vec_sub[3][5] , \out_r_vec_sub[3][4] , \out_r_vec_sub[3][3] ,
         \out_r_vec_sub[3][2] , \out_r_vec_sub[3][1] , \out_r_vec_sub[3][0] ,
         \out_i_vec_sub[0][11] , \out_i_vec_sub[0][10] , \out_i_vec_sub[0][9] ,
         \out_i_vec_sub[0][8] , \out_i_vec_sub[0][7] , \out_i_vec_sub[0][6] ,
         \out_i_vec_sub[0][5] , \out_i_vec_sub[0][4] , \out_i_vec_sub[0][3] ,
         \out_i_vec_sub[0][2] , \out_i_vec_sub[0][1] , \out_i_vec_sub[0][0] ,
         \out_i_vec_sub[1][11] , \out_i_vec_sub[1][10] , \out_i_vec_sub[1][9] ,
         \out_i_vec_sub[1][8] , \out_i_vec_sub[1][7] , \out_i_vec_sub[1][6] ,
         \out_i_vec_sub[1][5] , \out_i_vec_sub[1][4] , \out_i_vec_sub[1][3] ,
         \out_i_vec_sub[1][2] , \out_i_vec_sub[1][1] , \out_i_vec_sub[1][0] ,
         \out_i_vec_sub[2][11] , \out_i_vec_sub[2][10] , \out_i_vec_sub[2][9] ,
         \out_i_vec_sub[2][8] , \out_i_vec_sub[2][7] , \out_i_vec_sub[2][6] ,
         \out_i_vec_sub[2][5] , \out_i_vec_sub[2][4] , \out_i_vec_sub[2][3] ,
         \out_i_vec_sub[2][2] , \out_i_vec_sub[2][1] , \out_i_vec_sub[2][0] ,
         \out_i_vec_sub[3][11] , \out_i_vec_sub[3][10] , \out_i_vec_sub[3][9] ,
         \out_i_vec_sub[3][8] , \out_i_vec_sub[3][7] , \out_i_vec_sub[3][6] ,
         \out_i_vec_sub[3][5] , \out_i_vec_sub[3][4] , \out_i_vec_sub[3][3] ,
         \out_i_vec_sub[3][2] , \out_i_vec_sub[3][1] , \out_i_vec_sub[3][0] ,
         w_in_a_vec_sub, start_inv_sqrt, done_inv_sqrt, col_sel_AQ2_sel,
         wr_en_AQ_int, wr_en_AQ_sel, single_in_R_sel, col_sel_R_sel,
         in_b_vec_mult_sel, w_col_sel_AQ_sel, in_a_inner_prod_sel,
         in_b_inner_prod_sel;
  wire   [1:0] w_col_sel_AQ_mux;
  wire   [11:0] single_out_r_AQ;
  wire   [11:0] single_out_i_AQ;
  wire   [1:0] col_sel_AQ_int;
  wire   [1:0] row_sel_AQ;
  wire   [11:0] single_out_r_AQ2;
  wire   [11:0] single_out_i_AQ2;
  wire   [1:0] col_sel_AQ2_mux;
  wire   [1:0] row_sel_AQ2;
  wire   [11:0] single_in_r_R_mux;
  wire   [11:0] single_in_i_R_mux;
  wire   [1:0] col_sel_R_mux;
  wire   [1:0] row_sel_R;
  wire   [11:0] in_a_r_inner_prod_mux;
  wire   [11:0] in_a_i_inner_prod_mux;
  wire   [11:0] in_b_r_inner_prod_mux;
  wire   [11:0] in_b_i_inner_prod_mux;
  wire   [11:0] out_inner_prod_r;
  wire   [11:0] out_inner_prod_i;
  wire   [11:0] in_b_r_vec_mult_mux;
  wire   [11:0] in_b_i_vec_mult_mux;
  wire   [11:0] in_a_r_mult;
  wire   [11:0] out_mult;
  wire   [11:0] out_inv_sqrt;
  wire   [1:0] vec_in_AQ_sel;
  wire   [1:0] col_sel_AQ2_int;
  wire   [1:0] col_sel_R_int;
  wire   [1:0] w_col_sel_AQ_int;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;
  assign \out_R_i[3][11]  = 1'b0;
  assign \out_R_i[3][10]  = 1'b0;
  assign \out_R_i[3][9]  = 1'b0;
  assign \out_R_i[3][8]  = 1'b0;
  assign \out_R_i[3][7]  = 1'b0;
  assign \out_R_i[3][6]  = 1'b0;
  assign \out_R_i[3][5]  = 1'b0;
  assign \out_R_i[3][4]  = 1'b0;
  assign \out_R_i[3][3]  = 1'b0;
  assign \out_R_i[3][2]  = 1'b0;
  assign \out_R_i[3][1]  = 1'b0;
  assign \out_R_i[3][0]  = 1'b0;

  mat_regs_WORD_WIDTH12_N4_LOG2_N2 A_Q_mat ( .vector_in_r({
        \vec_in_r_AQ_mux[0][11] , \vec_in_r_AQ_mux[0][10] , 
        \vec_in_r_AQ_mux[0][9] , \vec_in_r_AQ_mux[0][8] , 
        \vec_in_r_AQ_mux[0][7] , \vec_in_r_AQ_mux[0][6] , 
        \vec_in_r_AQ_mux[0][5] , \vec_in_r_AQ_mux[0][4] , 
        \vec_in_r_AQ_mux[0][3] , \vec_in_r_AQ_mux[0][2] , 
        \vec_in_r_AQ_mux[0][1] , \vec_in_r_AQ_mux[0][0] , 
        \vec_in_r_AQ_mux[1][11] , \vec_in_r_AQ_mux[1][10] , 
        \vec_in_r_AQ_mux[1][9] , \vec_in_r_AQ_mux[1][8] , 
        \vec_in_r_AQ_mux[1][7] , \vec_in_r_AQ_mux[1][6] , 
        \vec_in_r_AQ_mux[1][5] , \vec_in_r_AQ_mux[1][4] , 
        \vec_in_r_AQ_mux[1][3] , \vec_in_r_AQ_mux[1][2] , 
        \vec_in_r_AQ_mux[1][1] , \vec_in_r_AQ_mux[1][0] , 
        \vec_in_r_AQ_mux[2][11] , \vec_in_r_AQ_mux[2][10] , 
        \vec_in_r_AQ_mux[2][9] , \vec_in_r_AQ_mux[2][8] , 
        \vec_in_r_AQ_mux[2][7] , \vec_in_r_AQ_mux[2][6] , 
        \vec_in_r_AQ_mux[2][5] , \vec_in_r_AQ_mux[2][4] , 
        \vec_in_r_AQ_mux[2][3] , \vec_in_r_AQ_mux[2][2] , 
        \vec_in_r_AQ_mux[2][1] , \vec_in_r_AQ_mux[2][0] , 
        \vec_in_r_AQ_mux[3][11] , \vec_in_r_AQ_mux[3][10] , 
        \vec_in_r_AQ_mux[3][9] , \vec_in_r_AQ_mux[3][8] , 
        \vec_in_r_AQ_mux[3][7] , \vec_in_r_AQ_mux[3][6] , 
        \vec_in_r_AQ_mux[3][5] , \vec_in_r_AQ_mux[3][4] , 
        \vec_in_r_AQ_mux[3][3] , \vec_in_r_AQ_mux[3][2] , 
        \vec_in_r_AQ_mux[3][1] , \vec_in_r_AQ_mux[3][0] }), .vector_in_i({
        \vec_in_i_AQ_mux[0][11] , \vec_in_i_AQ_mux[0][10] , 
        \vec_in_i_AQ_mux[0][9] , \vec_in_i_AQ_mux[0][8] , 
        \vec_in_i_AQ_mux[0][7] , \vec_in_i_AQ_mux[0][6] , 
        \vec_in_i_AQ_mux[0][5] , \vec_in_i_AQ_mux[0][4] , 
        \vec_in_i_AQ_mux[0][3] , \vec_in_i_AQ_mux[0][2] , 
        \vec_in_i_AQ_mux[0][1] , \vec_in_i_AQ_mux[0][0] , 
        \vec_in_i_AQ_mux[1][11] , \vec_in_i_AQ_mux[1][10] , 
        \vec_in_i_AQ_mux[1][9] , \vec_in_i_AQ_mux[1][8] , 
        \vec_in_i_AQ_mux[1][7] , \vec_in_i_AQ_mux[1][6] , 
        \vec_in_i_AQ_mux[1][5] , \vec_in_i_AQ_mux[1][4] , 
        \vec_in_i_AQ_mux[1][3] , \vec_in_i_AQ_mux[1][2] , 
        \vec_in_i_AQ_mux[1][1] , \vec_in_i_AQ_mux[1][0] , 
        \vec_in_i_AQ_mux[2][11] , \vec_in_i_AQ_mux[2][10] , 
        \vec_in_i_AQ_mux[2][9] , \vec_in_i_AQ_mux[2][8] , 
        \vec_in_i_AQ_mux[2][7] , \vec_in_i_AQ_mux[2][6] , 
        \vec_in_i_AQ_mux[2][5] , \vec_in_i_AQ_mux[2][4] , 
        \vec_in_i_AQ_mux[2][3] , \vec_in_i_AQ_mux[2][2] , 
        \vec_in_i_AQ_mux[2][1] , \vec_in_i_AQ_mux[2][0] , 
        \vec_in_i_AQ_mux[3][11] , \vec_in_i_AQ_mux[3][10] , 
        \vec_in_i_AQ_mux[3][9] , \vec_in_i_AQ_mux[3][8] , 
        \vec_in_i_AQ_mux[3][7] , \vec_in_i_AQ_mux[3][6] , 
        \vec_in_i_AQ_mux[3][5] , \vec_in_i_AQ_mux[3][4] , 
        \vec_in_i_AQ_mux[3][3] , \vec_in_i_AQ_mux[3][2] , 
        \vec_in_i_AQ_mux[3][1] , \vec_in_i_AQ_mux[3][0] }), .w_col_sel(
        w_col_sel_AQ_mux), .vector_out_r({\vec_out_r_AQ[0][11] , 
        \vec_out_r_AQ[0][10] , \vec_out_r_AQ[0][9] , \vec_out_r_AQ[0][8] , 
        \vec_out_r_AQ[0][7] , \vec_out_r_AQ[0][6] , \vec_out_r_AQ[0][5] , 
        \vec_out_r_AQ[0][4] , \vec_out_r_AQ[0][3] , \vec_out_r_AQ[0][2] , 
        \vec_out_r_AQ[0][1] , \vec_out_r_AQ[0][0] , \vec_out_r_AQ[1][11] , 
        \vec_out_r_AQ[1][10] , \vec_out_r_AQ[1][9] , \vec_out_r_AQ[1][8] , 
        \vec_out_r_AQ[1][7] , \vec_out_r_AQ[1][6] , \vec_out_r_AQ[1][5] , 
        \vec_out_r_AQ[1][4] , \vec_out_r_AQ[1][3] , \vec_out_r_AQ[1][2] , 
        \vec_out_r_AQ[1][1] , \vec_out_r_AQ[1][0] , \vec_out_r_AQ[2][11] , 
        \vec_out_r_AQ[2][10] , \vec_out_r_AQ[2][9] , \vec_out_r_AQ[2][8] , 
        \vec_out_r_AQ[2][7] , \vec_out_r_AQ[2][6] , \vec_out_r_AQ[2][5] , 
        \vec_out_r_AQ[2][4] , \vec_out_r_AQ[2][3] , \vec_out_r_AQ[2][2] , 
        \vec_out_r_AQ[2][1] , \vec_out_r_AQ[2][0] , \vec_out_r_AQ[3][11] , 
        \vec_out_r_AQ[3][10] , \vec_out_r_AQ[3][9] , \vec_out_r_AQ[3][8] , 
        \vec_out_r_AQ[3][7] , \vec_out_r_AQ[3][6] , \vec_out_r_AQ[3][5] , 
        \vec_out_r_AQ[3][4] , \vec_out_r_AQ[3][3] , \vec_out_r_AQ[3][2] , 
        \vec_out_r_AQ[3][1] , \vec_out_r_AQ[3][0] }), .vector_out_i({
        \vec_out_i_AQ[0][11] , \vec_out_i_AQ[0][10] , \vec_out_i_AQ[0][9] , 
        \vec_out_i_AQ[0][8] , \vec_out_i_AQ[0][7] , \vec_out_i_AQ[0][6] , 
        \vec_out_i_AQ[0][5] , \vec_out_i_AQ[0][4] , \vec_out_i_AQ[0][3] , 
        \vec_out_i_AQ[0][2] , \vec_out_i_AQ[0][1] , \vec_out_i_AQ[0][0] , 
        \vec_out_i_AQ[1][11] , \vec_out_i_AQ[1][10] , \vec_out_i_AQ[1][9] , 
        \vec_out_i_AQ[1][8] , \vec_out_i_AQ[1][7] , \vec_out_i_AQ[1][6] , 
        \vec_out_i_AQ[1][5] , \vec_out_i_AQ[1][4] , \vec_out_i_AQ[1][3] , 
        \vec_out_i_AQ[1][2] , \vec_out_i_AQ[1][1] , \vec_out_i_AQ[1][0] , 
        \vec_out_i_AQ[2][11] , \vec_out_i_AQ[2][10] , \vec_out_i_AQ[2][9] , 
        \vec_out_i_AQ[2][8] , \vec_out_i_AQ[2][7] , \vec_out_i_AQ[2][6] , 
        \vec_out_i_AQ[2][5] , \vec_out_i_AQ[2][4] , \vec_out_i_AQ[2][3] , 
        \vec_out_i_AQ[2][2] , \vec_out_i_AQ[2][1] , \vec_out_i_AQ[2][0] , 
        \vec_out_i_AQ[3][11] , \vec_out_i_AQ[3][10] , \vec_out_i_AQ[3][9] , 
        \vec_out_i_AQ[3][8] , \vec_out_i_AQ[3][7] , \vec_out_i_AQ[3][6] , 
        \vec_out_i_AQ[3][5] , \vec_out_i_AQ[3][4] , \vec_out_i_AQ[3][3] , 
        \vec_out_i_AQ[3][2] , \vec_out_i_AQ[3][1] , \vec_out_i_AQ[3][0] }), 
        .single_out_r(single_out_r_AQ), .single_out_i(single_out_i_AQ), 
        .col_sel(col_sel_AQ_int), .row_sel(row_sel_AQ), .vector_out_r2({
        \out_Q_r[0][11] , \out_Q_r[0][10] , \out_Q_r[0][9] , \out_Q_r[0][8] , 
        \out_Q_r[0][7] , \out_Q_r[0][6] , \out_Q_r[0][5] , \out_Q_r[0][4] , 
        \out_Q_r[0][3] , \out_Q_r[0][2] , \out_Q_r[0][1] , \out_Q_r[0][0] , 
        \out_Q_r[1][11] , \out_Q_r[1][10] , \out_Q_r[1][9] , \out_Q_r[1][8] , 
        \out_Q_r[1][7] , \out_Q_r[1][6] , \out_Q_r[1][5] , \out_Q_r[1][4] , 
        \out_Q_r[1][3] , \out_Q_r[1][2] , \out_Q_r[1][1] , \out_Q_r[1][0] , 
        \out_Q_r[2][11] , \out_Q_r[2][10] , \out_Q_r[2][9] , \out_Q_r[2][8] , 
        \out_Q_r[2][7] , \out_Q_r[2][6] , \out_Q_r[2][5] , \out_Q_r[2][4] , 
        \out_Q_r[2][3] , \out_Q_r[2][2] , \out_Q_r[2][1] , \out_Q_r[2][0] , 
        \out_Q_r[3][11] , \out_Q_r[3][10] , \out_Q_r[3][9] , \out_Q_r[3][8] , 
        \out_Q_r[3][7] , \out_Q_r[3][6] , \out_Q_r[3][5] , \out_Q_r[3][4] , 
        \out_Q_r[3][3] , \out_Q_r[3][2] , \out_Q_r[3][1] , \out_Q_r[3][0] }), 
        .vector_out_i2({\out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] , 
        \out_Q_i[0][8] , \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] , 
        \out_Q_i[0][4] , \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] , 
        \out_Q_i[0][0] , \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] , 
        \out_Q_i[1][8] , \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] , 
        \out_Q_i[1][4] , \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] , 
        \out_Q_i[1][0] , \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] , 
        \out_Q_i[2][8] , \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] , 
        \out_Q_i[2][4] , \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] , 
        \out_Q_i[2][0] , \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] , 
        \out_Q_i[3][8] , \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] , 
        \out_Q_i[3][4] , \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] , 
        \out_Q_i[3][0] }), .single_out_r2(single_out_r_AQ2), .single_out_i2(
        single_out_i_AQ2), .col_sel2(col_sel_AQ2_mux), .row_sel2(row_sel_AQ2), 
        .clk(clk), .wr_enable(wr_en_AQ_mux) );
  r_mat_regs_WORD_WIDTH12_N4_LOG2_N2 R_mat ( .single_in_r(single_in_r_R_mux), 
        .single_in_i(single_in_i_R_mux), .vector_out_r({\out_R_r[0][11] , 
        \out_R_r[0][10] , \out_R_r[0][9] , \out_R_r[0][8] , \out_R_r[0][7] , 
        \out_R_r[0][6] , \out_R_r[0][5] , \out_R_r[0][4] , \out_R_r[0][3] , 
        \out_R_r[0][2] , \out_R_r[0][1] , \out_R_r[0][0] , \out_R_r[1][11] , 
        \out_R_r[1][10] , \out_R_r[1][9] , \out_R_r[1][8] , \out_R_r[1][7] , 
        \out_R_r[1][6] , \out_R_r[1][5] , \out_R_r[1][4] , \out_R_r[1][3] , 
        \out_R_r[1][2] , \out_R_r[1][1] , \out_R_r[1][0] , \out_R_r[2][11] , 
        \out_R_r[2][10] , \out_R_r[2][9] , \out_R_r[2][8] , \out_R_r[2][7] , 
        \out_R_r[2][6] , \out_R_r[2][5] , \out_R_r[2][4] , \out_R_r[2][3] , 
        \out_R_r[2][2] , \out_R_r[2][1] , \out_R_r[2][0] , \out_R_r[3][11] , 
        \out_R_r[3][10] , \out_R_r[3][9] , \out_R_r[3][8] , \out_R_r[3][7] , 
        \out_R_r[3][6] , \out_R_r[3][5] , \out_R_r[3][4] , \out_R_r[3][3] , 
        \out_R_r[3][2] , \out_R_r[3][1] , \out_R_r[3][0] }), .vector_out_i({
        \out_R_i[0][11] , \out_R_i[0][10] , \out_R_i[0][9] , \out_R_i[0][8] , 
        \out_R_i[0][7] , \out_R_i[0][6] , \out_R_i[0][5] , \out_R_i[0][4] , 
        \out_R_i[0][3] , \out_R_i[0][2] , \out_R_i[0][1] , \out_R_i[0][0] , 
        \out_R_i[1][11] , \out_R_i[1][10] , \out_R_i[1][9] , \out_R_i[1][8] , 
        \out_R_i[1][7] , \out_R_i[1][6] , \out_R_i[1][5] , \out_R_i[1][4] , 
        \out_R_i[1][3] , \out_R_i[1][2] , \out_R_i[1][1] , \out_R_i[1][0] , 
        \out_R_i[2][11] , \out_R_i[2][10] , \out_R_i[2][9] , \out_R_i[2][8] , 
        \out_R_i[2][7] , \out_R_i[2][6] , \out_R_i[2][5] , \out_R_i[2][4] , 
        \out_R_i[2][3] , \out_R_i[2][2] , \out_R_i[2][1] , \out_R_i[2][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}), .col_sel(
        col_sel_R_mux), .row_sel(row_sel_R), .clk(clk), .wr_enable(wr_en_R) );
  inner_prod_INT_BITS4_WORD_WIDTH12_N4 inner_prod_inst ( .clk(clk), .rst(rst), 
        .in_a_r(in_a_r_inner_prod_mux), .in_a_i(in_a_i_inner_prod_mux), 
        .in_b_r(in_b_r_inner_prod_mux), .in_b_i(in_b_i_inner_prod_mux), 
        .out_r(out_inner_prod_r), .out_i(out_inner_prod_i), .reduced_matrix(
        red_mat_reg), .start(start_inner_prod), .done(done_inner_prod) );
  vec_mult_N4_WORD_WIDTH12_INT_BITS4 vec_mult_inst ( .in_a_r({
        \vec_out_r_AQ[0][11] , \vec_out_r_AQ[0][10] , \vec_out_r_AQ[0][9] , 
        \vec_out_r_AQ[0][8] , \vec_out_r_AQ[0][7] , \vec_out_r_AQ[0][6] , 
        \vec_out_r_AQ[0][5] , \vec_out_r_AQ[0][4] , \vec_out_r_AQ[0][3] , 
        \vec_out_r_AQ[0][2] , \vec_out_r_AQ[0][1] , \vec_out_r_AQ[0][0] , 
        \vec_out_r_AQ[1][11] , \vec_out_r_AQ[1][10] , \vec_out_r_AQ[1][9] , 
        \vec_out_r_AQ[1][8] , \vec_out_r_AQ[1][7] , \vec_out_r_AQ[1][6] , 
        \vec_out_r_AQ[1][5] , \vec_out_r_AQ[1][4] , \vec_out_r_AQ[1][3] , 
        \vec_out_r_AQ[1][2] , \vec_out_r_AQ[1][1] , \vec_out_r_AQ[1][0] , 
        \vec_out_r_AQ[2][11] , \vec_out_r_AQ[2][10] , \vec_out_r_AQ[2][9] , 
        \vec_out_r_AQ[2][8] , \vec_out_r_AQ[2][7] , \vec_out_r_AQ[2][6] , 
        \vec_out_r_AQ[2][5] , \vec_out_r_AQ[2][4] , \vec_out_r_AQ[2][3] , 
        \vec_out_r_AQ[2][2] , \vec_out_r_AQ[2][1] , \vec_out_r_AQ[2][0] , 
        \vec_out_r_AQ[3][11] , \vec_out_r_AQ[3][10] , \vec_out_r_AQ[3][9] , 
        \vec_out_r_AQ[3][8] , \vec_out_r_AQ[3][7] , \vec_out_r_AQ[3][6] , 
        \vec_out_r_AQ[3][5] , \vec_out_r_AQ[3][4] , \vec_out_r_AQ[3][3] , 
        \vec_out_r_AQ[3][2] , \vec_out_r_AQ[3][1] , \vec_out_r_AQ[3][0] }), 
        .in_a_i({\vec_out_i_AQ[0][11] , \vec_out_i_AQ[0][10] , 
        \vec_out_i_AQ[0][9] , \vec_out_i_AQ[0][8] , \vec_out_i_AQ[0][7] , 
        \vec_out_i_AQ[0][6] , \vec_out_i_AQ[0][5] , \vec_out_i_AQ[0][4] , 
        \vec_out_i_AQ[0][3] , \vec_out_i_AQ[0][2] , \vec_out_i_AQ[0][1] , 
        \vec_out_i_AQ[0][0] , \vec_out_i_AQ[1][11] , \vec_out_i_AQ[1][10] , 
        \vec_out_i_AQ[1][9] , \vec_out_i_AQ[1][8] , \vec_out_i_AQ[1][7] , 
        \vec_out_i_AQ[1][6] , \vec_out_i_AQ[1][5] , \vec_out_i_AQ[1][4] , 
        \vec_out_i_AQ[1][3] , \vec_out_i_AQ[1][2] , \vec_out_i_AQ[1][1] , 
        \vec_out_i_AQ[1][0] , \vec_out_i_AQ[2][11] , \vec_out_i_AQ[2][10] , 
        \vec_out_i_AQ[2][9] , \vec_out_i_AQ[2][8] , \vec_out_i_AQ[2][7] , 
        \vec_out_i_AQ[2][6] , \vec_out_i_AQ[2][5] , \vec_out_i_AQ[2][4] , 
        \vec_out_i_AQ[2][3] , \vec_out_i_AQ[2][2] , \vec_out_i_AQ[2][1] , 
        \vec_out_i_AQ[2][0] , \vec_out_i_AQ[3][11] , \vec_out_i_AQ[3][10] , 
        \vec_out_i_AQ[3][9] , \vec_out_i_AQ[3][8] , \vec_out_i_AQ[3][7] , 
        \vec_out_i_AQ[3][6] , \vec_out_i_AQ[3][5] , \vec_out_i_AQ[3][4] , 
        \vec_out_i_AQ[3][3] , \vec_out_i_AQ[3][2] , \vec_out_i_AQ[3][1] , 
        \vec_out_i_AQ[3][0] }), .in_b_r(in_b_r_vec_mult_mux), .in_b_i(
        in_b_i_vec_mult_mux), .out_r({\out_r_vec_mult[0][11] , 
        \out_r_vec_mult[0][10] , \out_r_vec_mult[0][9] , 
        \out_r_vec_mult[0][8] , \out_r_vec_mult[0][7] , \out_r_vec_mult[0][6] , 
        \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] , \out_r_vec_mult[0][3] , 
        \out_r_vec_mult[0][2] , \out_r_vec_mult[0][1] , \out_r_vec_mult[0][0] , 
        \out_r_vec_mult[1][11] , \out_r_vec_mult[1][10] , 
        \out_r_vec_mult[1][9] , \out_r_vec_mult[1][8] , \out_r_vec_mult[1][7] , 
        \out_r_vec_mult[1][6] , \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] , 
        \out_r_vec_mult[1][3] , \out_r_vec_mult[1][2] , \out_r_vec_mult[1][1] , 
        \out_r_vec_mult[1][0] , \out_r_vec_mult[2][11] , 
        \out_r_vec_mult[2][10] , \out_r_vec_mult[2][9] , 
        \out_r_vec_mult[2][8] , \out_r_vec_mult[2][7] , \out_r_vec_mult[2][6] , 
        \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] , \out_r_vec_mult[2][3] , 
        \out_r_vec_mult[2][2] , \out_r_vec_mult[2][1] , \out_r_vec_mult[2][0] , 
        \out_r_vec_mult[3][11] , \out_r_vec_mult[3][10] , 
        \out_r_vec_mult[3][9] , \out_r_vec_mult[3][8] , \out_r_vec_mult[3][7] , 
        \out_r_vec_mult[3][6] , \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] , 
        \out_r_vec_mult[3][3] , \out_r_vec_mult[3][2] , \out_r_vec_mult[3][1] , 
        \out_r_vec_mult[3][0] }), .out_i({\out_i_vec_mult[0][11] , 
        \out_i_vec_mult[0][10] , \out_i_vec_mult[0][9] , 
        \out_i_vec_mult[0][8] , \out_i_vec_mult[0][7] , \out_i_vec_mult[0][6] , 
        \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] , \out_i_vec_mult[0][3] , 
        \out_i_vec_mult[0][2] , \out_i_vec_mult[0][1] , \out_i_vec_mult[0][0] , 
        \out_i_vec_mult[1][11] , \out_i_vec_mult[1][10] , 
        \out_i_vec_mult[1][9] , \out_i_vec_mult[1][8] , \out_i_vec_mult[1][7] , 
        \out_i_vec_mult[1][6] , \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] , 
        \out_i_vec_mult[1][3] , \out_i_vec_mult[1][2] , \out_i_vec_mult[1][1] , 
        \out_i_vec_mult[1][0] , \out_i_vec_mult[2][11] , 
        \out_i_vec_mult[2][10] , \out_i_vec_mult[2][9] , 
        \out_i_vec_mult[2][8] , \out_i_vec_mult[2][7] , \out_i_vec_mult[2][6] , 
        \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] , \out_i_vec_mult[2][3] , 
        \out_i_vec_mult[2][2] , \out_i_vec_mult[2][1] , \out_i_vec_mult[2][0] , 
        \out_i_vec_mult[3][11] , \out_i_vec_mult[3][10] , 
        \out_i_vec_mult[3][9] , \out_i_vec_mult[3][8] , \out_i_vec_mult[3][7] , 
        \out_i_vec_mult[3][6] , \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] , 
        \out_i_vec_mult[3][3] , \out_i_vec_mult[3][2] , \out_i_vec_mult[3][1] , 
        \out_i_vec_mult[3][0] }), .clk(clk) );
  vec_sub_N4_WORD_WIDTH12 vec_sub_inst ( .in_a_r({\out_Q_r[0][11] , 
        \out_Q_r[0][10] , \out_Q_r[0][9] , \out_Q_r[0][8] , \out_Q_r[0][7] , 
        \out_Q_r[0][6] , \out_Q_r[0][5] , \out_Q_r[0][4] , \out_Q_r[0][3] , 
        \out_Q_r[0][2] , \out_Q_r[0][1] , \out_Q_r[0][0] , \out_Q_r[1][11] , 
        \out_Q_r[1][10] , \out_Q_r[1][9] , \out_Q_r[1][8] , \out_Q_r[1][7] , 
        \out_Q_r[1][6] , \out_Q_r[1][5] , \out_Q_r[1][4] , \out_Q_r[1][3] , 
        \out_Q_r[1][2] , \out_Q_r[1][1] , \out_Q_r[1][0] , \out_Q_r[2][11] , 
        \out_Q_r[2][10] , \out_Q_r[2][9] , \out_Q_r[2][8] , \out_Q_r[2][7] , 
        \out_Q_r[2][6] , \out_Q_r[2][5] , \out_Q_r[2][4] , \out_Q_r[2][3] , 
        \out_Q_r[2][2] , \out_Q_r[2][1] , \out_Q_r[2][0] , \out_Q_r[3][11] , 
        \out_Q_r[3][10] , \out_Q_r[3][9] , \out_Q_r[3][8] , \out_Q_r[3][7] , 
        \out_Q_r[3][6] , \out_Q_r[3][5] , \out_Q_r[3][4] , \out_Q_r[3][3] , 
        \out_Q_r[3][2] , \out_Q_r[3][1] , \out_Q_r[3][0] }), .in_a_i({
        \out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] , \out_Q_i[0][8] , 
        \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] , \out_Q_i[0][4] , 
        \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] , \out_Q_i[0][0] , 
        \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] , \out_Q_i[1][8] , 
        \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] , \out_Q_i[1][4] , 
        \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] , \out_Q_i[1][0] , 
        \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] , \out_Q_i[2][8] , 
        \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] , \out_Q_i[2][4] , 
        \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] , \out_Q_i[2][0] , 
        \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] , \out_Q_i[3][8] , 
        \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] , \out_Q_i[3][4] , 
        \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] , \out_Q_i[3][0] }), 
        .in_b_r({\out_r_vec_mult[0][11] , \out_r_vec_mult[0][10] , 
        \out_r_vec_mult[0][9] , \out_r_vec_mult[0][8] , \out_r_vec_mult[0][7] , 
        \out_r_vec_mult[0][6] , \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] , 
        \out_r_vec_mult[0][3] , \out_r_vec_mult[0][2] , \out_r_vec_mult[0][1] , 
        \out_r_vec_mult[0][0] , \out_r_vec_mult[1][11] , 
        \out_r_vec_mult[1][10] , \out_r_vec_mult[1][9] , 
        \out_r_vec_mult[1][8] , \out_r_vec_mult[1][7] , \out_r_vec_mult[1][6] , 
        \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] , \out_r_vec_mult[1][3] , 
        \out_r_vec_mult[1][2] , \out_r_vec_mult[1][1] , \out_r_vec_mult[1][0] , 
        \out_r_vec_mult[2][11] , \out_r_vec_mult[2][10] , 
        \out_r_vec_mult[2][9] , \out_r_vec_mult[2][8] , \out_r_vec_mult[2][7] , 
        \out_r_vec_mult[2][6] , \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] , 
        \out_r_vec_mult[2][3] , \out_r_vec_mult[2][2] , \out_r_vec_mult[2][1] , 
        \out_r_vec_mult[2][0] , \out_r_vec_mult[3][11] , 
        \out_r_vec_mult[3][10] , \out_r_vec_mult[3][9] , 
        \out_r_vec_mult[3][8] , \out_r_vec_mult[3][7] , \out_r_vec_mult[3][6] , 
        \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] , \out_r_vec_mult[3][3] , 
        \out_r_vec_mult[3][2] , \out_r_vec_mult[3][1] , \out_r_vec_mult[3][0] }), .in_b_i({\out_i_vec_mult[0][11] , \out_i_vec_mult[0][10] , 
        \out_i_vec_mult[0][9] , \out_i_vec_mult[0][8] , \out_i_vec_mult[0][7] , 
        \out_i_vec_mult[0][6] , \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] , 
        \out_i_vec_mult[0][3] , \out_i_vec_mult[0][2] , \out_i_vec_mult[0][1] , 
        \out_i_vec_mult[0][0] , \out_i_vec_mult[1][11] , 
        \out_i_vec_mult[1][10] , \out_i_vec_mult[1][9] , 
        \out_i_vec_mult[1][8] , \out_i_vec_mult[1][7] , \out_i_vec_mult[1][6] , 
        \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] , \out_i_vec_mult[1][3] , 
        \out_i_vec_mult[1][2] , \out_i_vec_mult[1][1] , \out_i_vec_mult[1][0] , 
        \out_i_vec_mult[2][11] , \out_i_vec_mult[2][10] , 
        \out_i_vec_mult[2][9] , \out_i_vec_mult[2][8] , \out_i_vec_mult[2][7] , 
        \out_i_vec_mult[2][6] , \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] , 
        \out_i_vec_mult[2][3] , \out_i_vec_mult[2][2] , \out_i_vec_mult[2][1] , 
        \out_i_vec_mult[2][0] , \out_i_vec_mult[3][11] , 
        \out_i_vec_mult[3][10] , \out_i_vec_mult[3][9] , 
        \out_i_vec_mult[3][8] , \out_i_vec_mult[3][7] , \out_i_vec_mult[3][6] , 
        \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] , \out_i_vec_mult[3][3] , 
        \out_i_vec_mult[3][2] , \out_i_vec_mult[3][1] , \out_i_vec_mult[3][0] }), .out_r({\out_r_vec_sub[0][11] , \out_r_vec_sub[0][10] , 
        \out_r_vec_sub[0][9] , \out_r_vec_sub[0][8] , \out_r_vec_sub[0][7] , 
        \out_r_vec_sub[0][6] , \out_r_vec_sub[0][5] , \out_r_vec_sub[0][4] , 
        \out_r_vec_sub[0][3] , \out_r_vec_sub[0][2] , \out_r_vec_sub[0][1] , 
        \out_r_vec_sub[0][0] , \out_r_vec_sub[1][11] , \out_r_vec_sub[1][10] , 
        \out_r_vec_sub[1][9] , \out_r_vec_sub[1][8] , \out_r_vec_sub[1][7] , 
        \out_r_vec_sub[1][6] , \out_r_vec_sub[1][5] , \out_r_vec_sub[1][4] , 
        \out_r_vec_sub[1][3] , \out_r_vec_sub[1][2] , \out_r_vec_sub[1][1] , 
        \out_r_vec_sub[1][0] , \out_r_vec_sub[2][11] , \out_r_vec_sub[2][10] , 
        \out_r_vec_sub[2][9] , \out_r_vec_sub[2][8] , \out_r_vec_sub[2][7] , 
        \out_r_vec_sub[2][6] , \out_r_vec_sub[2][5] , \out_r_vec_sub[2][4] , 
        \out_r_vec_sub[2][3] , \out_r_vec_sub[2][2] , \out_r_vec_sub[2][1] , 
        \out_r_vec_sub[2][0] , \out_r_vec_sub[3][11] , \out_r_vec_sub[3][10] , 
        \out_r_vec_sub[3][9] , \out_r_vec_sub[3][8] , \out_r_vec_sub[3][7] , 
        \out_r_vec_sub[3][6] , \out_r_vec_sub[3][5] , \out_r_vec_sub[3][4] , 
        \out_r_vec_sub[3][3] , \out_r_vec_sub[3][2] , \out_r_vec_sub[3][1] , 
        \out_r_vec_sub[3][0] }), .out_i({\out_i_vec_sub[0][11] , 
        \out_i_vec_sub[0][10] , \out_i_vec_sub[0][9] , \out_i_vec_sub[0][8] , 
        \out_i_vec_sub[0][7] , \out_i_vec_sub[0][6] , \out_i_vec_sub[0][5] , 
        \out_i_vec_sub[0][4] , \out_i_vec_sub[0][3] , \out_i_vec_sub[0][2] , 
        \out_i_vec_sub[0][1] , \out_i_vec_sub[0][0] , \out_i_vec_sub[1][11] , 
        \out_i_vec_sub[1][10] , \out_i_vec_sub[1][9] , \out_i_vec_sub[1][8] , 
        \out_i_vec_sub[1][7] , \out_i_vec_sub[1][6] , \out_i_vec_sub[1][5] , 
        \out_i_vec_sub[1][4] , \out_i_vec_sub[1][3] , \out_i_vec_sub[1][2] , 
        \out_i_vec_sub[1][1] , \out_i_vec_sub[1][0] , \out_i_vec_sub[2][11] , 
        \out_i_vec_sub[2][10] , \out_i_vec_sub[2][9] , \out_i_vec_sub[2][8] , 
        \out_i_vec_sub[2][7] , \out_i_vec_sub[2][6] , \out_i_vec_sub[2][5] , 
        \out_i_vec_sub[2][4] , \out_i_vec_sub[2][3] , \out_i_vec_sub[2][2] , 
        \out_i_vec_sub[2][1] , \out_i_vec_sub[2][0] , \out_i_vec_sub[3][11] , 
        \out_i_vec_sub[3][10] , \out_i_vec_sub[3][9] , \out_i_vec_sub[3][8] , 
        \out_i_vec_sub[3][7] , \out_i_vec_sub[3][6] , \out_i_vec_sub[3][5] , 
        \out_i_vec_sub[3][4] , \out_i_vec_sub[3][3] , \out_i_vec_sub[3][2] , 
        \out_i_vec_sub[3][1] , \out_i_vec_sub[3][0] }), .w_in_a(w_in_a_vec_sub), .clk(clk) );
  mult_with_reg_WORD_WIDTH12_INT_BITS4_USE_SAT1 r_mult ( .in_a(in_a_r_mult), 
        .in_b(out_inner_prod_r), .clk(clk), .\output (out_mult) );
  inv_sqrt_INT_BITS4_WORD_WIDTH12_LOG_WORD_WIDTH4_USE_NEWTON1_SMALLER_POW2_WW16 inv_sqrt_inst ( 
        .\input (out_inner_prod_r), .\output (out_inv_sqrt), .clk(clk), .rst(
        rst), .start(start_inv_sqrt), .done(done_inv_sqrt) );
  qr_decomp_ctl_mux_1 muxes ( .in_A_r({\in_A_r[0][11] , \in_A_r[0][10] , 
        \in_A_r[0][9] , \in_A_r[0][8] , \in_A_r[0][7] , \in_A_r[0][6] , 
        \in_A_r[0][5] , \in_A_r[0][4] , \in_A_r[0][3] , \in_A_r[0][2] , 
        \in_A_r[0][1] , \in_A_r[0][0] , \in_A_r[1][11] , \in_A_r[1][10] , 
        \in_A_r[1][9] , \in_A_r[1][8] , \in_A_r[1][7] , \in_A_r[1][6] , 
        \in_A_r[1][5] , \in_A_r[1][4] , \in_A_r[1][3] , \in_A_r[1][2] , 
        \in_A_r[1][1] , \in_A_r[1][0] , \in_A_r[2][11] , \in_A_r[2][10] , 
        \in_A_r[2][9] , \in_A_r[2][8] , \in_A_r[2][7] , \in_A_r[2][6] , 
        \in_A_r[2][5] , \in_A_r[2][4] , \in_A_r[2][3] , \in_A_r[2][2] , 
        \in_A_r[2][1] , \in_A_r[2][0] , \in_A_r[3][11] , \in_A_r[3][10] , 
        \in_A_r[3][9] , \in_A_r[3][8] , \in_A_r[3][7] , \in_A_r[3][6] , 
        \in_A_r[3][5] , \in_A_r[3][4] , \in_A_r[3][3] , \in_A_r[3][2] , 
        \in_A_r[3][1] , \in_A_r[3][0] }), .out_r_vec_mult({
        \out_r_vec_mult[0][11] , \out_r_vec_mult[0][10] , 
        \out_r_vec_mult[0][9] , \out_r_vec_mult[0][8] , \out_r_vec_mult[0][7] , 
        \out_r_vec_mult[0][6] , \out_r_vec_mult[0][5] , \out_r_vec_mult[0][4] , 
        \out_r_vec_mult[0][3] , \out_r_vec_mult[0][2] , \out_r_vec_mult[0][1] , 
        \out_r_vec_mult[0][0] , \out_r_vec_mult[1][11] , 
        \out_r_vec_mult[1][10] , \out_r_vec_mult[1][9] , 
        \out_r_vec_mult[1][8] , \out_r_vec_mult[1][7] , \out_r_vec_mult[1][6] , 
        \out_r_vec_mult[1][5] , \out_r_vec_mult[1][4] , \out_r_vec_mult[1][3] , 
        \out_r_vec_mult[1][2] , \out_r_vec_mult[1][1] , \out_r_vec_mult[1][0] , 
        \out_r_vec_mult[2][11] , \out_r_vec_mult[2][10] , 
        \out_r_vec_mult[2][9] , \out_r_vec_mult[2][8] , \out_r_vec_mult[2][7] , 
        \out_r_vec_mult[2][6] , \out_r_vec_mult[2][5] , \out_r_vec_mult[2][4] , 
        \out_r_vec_mult[2][3] , \out_r_vec_mult[2][2] , \out_r_vec_mult[2][1] , 
        \out_r_vec_mult[2][0] , \out_r_vec_mult[3][11] , 
        \out_r_vec_mult[3][10] , \out_r_vec_mult[3][9] , 
        \out_r_vec_mult[3][8] , \out_r_vec_mult[3][7] , \out_r_vec_mult[3][6] , 
        \out_r_vec_mult[3][5] , \out_r_vec_mult[3][4] , \out_r_vec_mult[3][3] , 
        \out_r_vec_mult[3][2] , \out_r_vec_mult[3][1] , \out_r_vec_mult[3][0] }), .out_r_vec_sub({\out_r_vec_sub[0][11] , \out_r_vec_sub[0][10] , 
        \out_r_vec_sub[0][9] , \out_r_vec_sub[0][8] , \out_r_vec_sub[0][7] , 
        \out_r_vec_sub[0][6] , \out_r_vec_sub[0][5] , \out_r_vec_sub[0][4] , 
        \out_r_vec_sub[0][3] , \out_r_vec_sub[0][2] , \out_r_vec_sub[0][1] , 
        \out_r_vec_sub[0][0] , \out_r_vec_sub[1][11] , \out_r_vec_sub[1][10] , 
        \out_r_vec_sub[1][9] , \out_r_vec_sub[1][8] , \out_r_vec_sub[1][7] , 
        \out_r_vec_sub[1][6] , \out_r_vec_sub[1][5] , \out_r_vec_sub[1][4] , 
        \out_r_vec_sub[1][3] , \out_r_vec_sub[1][2] , \out_r_vec_sub[1][1] , 
        \out_r_vec_sub[1][0] , \out_r_vec_sub[2][11] , \out_r_vec_sub[2][10] , 
        \out_r_vec_sub[2][9] , \out_r_vec_sub[2][8] , \out_r_vec_sub[2][7] , 
        \out_r_vec_sub[2][6] , \out_r_vec_sub[2][5] , \out_r_vec_sub[2][4] , 
        \out_r_vec_sub[2][3] , \out_r_vec_sub[2][2] , \out_r_vec_sub[2][1] , 
        \out_r_vec_sub[2][0] , \out_r_vec_sub[3][11] , \out_r_vec_sub[3][10] , 
        \out_r_vec_sub[3][9] , \out_r_vec_sub[3][8] , \out_r_vec_sub[3][7] , 
        \out_r_vec_sub[3][6] , \out_r_vec_sub[3][5] , \out_r_vec_sub[3][4] , 
        \out_r_vec_sub[3][3] , \out_r_vec_sub[3][2] , \out_r_vec_sub[3][1] , 
        \out_r_vec_sub[3][0] }), .vec_in_r_AQ_mux({\vec_in_r_AQ_mux[0][11] , 
        \vec_in_r_AQ_mux[0][10] , \vec_in_r_AQ_mux[0][9] , 
        \vec_in_r_AQ_mux[0][8] , \vec_in_r_AQ_mux[0][7] , 
        \vec_in_r_AQ_mux[0][6] , \vec_in_r_AQ_mux[0][5] , 
        \vec_in_r_AQ_mux[0][4] , \vec_in_r_AQ_mux[0][3] , 
        \vec_in_r_AQ_mux[0][2] , \vec_in_r_AQ_mux[0][1] , 
        \vec_in_r_AQ_mux[0][0] , \vec_in_r_AQ_mux[1][11] , 
        \vec_in_r_AQ_mux[1][10] , \vec_in_r_AQ_mux[1][9] , 
        \vec_in_r_AQ_mux[1][8] , \vec_in_r_AQ_mux[1][7] , 
        \vec_in_r_AQ_mux[1][6] , \vec_in_r_AQ_mux[1][5] , 
        \vec_in_r_AQ_mux[1][4] , \vec_in_r_AQ_mux[1][3] , 
        \vec_in_r_AQ_mux[1][2] , \vec_in_r_AQ_mux[1][1] , 
        \vec_in_r_AQ_mux[1][0] , \vec_in_r_AQ_mux[2][11] , 
        \vec_in_r_AQ_mux[2][10] , \vec_in_r_AQ_mux[2][9] , 
        \vec_in_r_AQ_mux[2][8] , \vec_in_r_AQ_mux[2][7] , 
        \vec_in_r_AQ_mux[2][6] , \vec_in_r_AQ_mux[2][5] , 
        \vec_in_r_AQ_mux[2][4] , \vec_in_r_AQ_mux[2][3] , 
        \vec_in_r_AQ_mux[2][2] , \vec_in_r_AQ_mux[2][1] , 
        \vec_in_r_AQ_mux[2][0] , \vec_in_r_AQ_mux[3][11] , 
        \vec_in_r_AQ_mux[3][10] , \vec_in_r_AQ_mux[3][9] , 
        \vec_in_r_AQ_mux[3][8] , \vec_in_r_AQ_mux[3][7] , 
        \vec_in_r_AQ_mux[3][6] , \vec_in_r_AQ_mux[3][5] , 
        \vec_in_r_AQ_mux[3][4] , \vec_in_r_AQ_mux[3][3] , 
        \vec_in_r_AQ_mux[3][2] , \vec_in_r_AQ_mux[3][1] , 
        \vec_in_r_AQ_mux[3][0] }), .in_A_i({\in_A_i[0][11] , \in_A_i[0][10] , 
        \in_A_i[0][9] , \in_A_i[0][8] , \in_A_i[0][7] , \in_A_i[0][6] , 
        \in_A_i[0][5] , \in_A_i[0][4] , \in_A_i[0][3] , \in_A_i[0][2] , 
        \in_A_i[0][1] , \in_A_i[0][0] , \in_A_i[1][11] , \in_A_i[1][10] , 
        \in_A_i[1][9] , \in_A_i[1][8] , \in_A_i[1][7] , \in_A_i[1][6] , 
        \in_A_i[1][5] , \in_A_i[1][4] , \in_A_i[1][3] , \in_A_i[1][2] , 
        \in_A_i[1][1] , \in_A_i[1][0] , \in_A_i[2][11] , \in_A_i[2][10] , 
        \in_A_i[2][9] , \in_A_i[2][8] , \in_A_i[2][7] , \in_A_i[2][6] , 
        \in_A_i[2][5] , \in_A_i[2][4] , \in_A_i[2][3] , \in_A_i[2][2] , 
        \in_A_i[2][1] , \in_A_i[2][0] , \in_A_i[3][11] , \in_A_i[3][10] , 
        \in_A_i[3][9] , \in_A_i[3][8] , \in_A_i[3][7] , \in_A_i[3][6] , 
        \in_A_i[3][5] , \in_A_i[3][4] , \in_A_i[3][3] , \in_A_i[3][2] , 
        \in_A_i[3][1] , \in_A_i[3][0] }), .out_i_vec_mult({
        \out_i_vec_mult[0][11] , \out_i_vec_mult[0][10] , 
        \out_i_vec_mult[0][9] , \out_i_vec_mult[0][8] , \out_i_vec_mult[0][7] , 
        \out_i_vec_mult[0][6] , \out_i_vec_mult[0][5] , \out_i_vec_mult[0][4] , 
        \out_i_vec_mult[0][3] , \out_i_vec_mult[0][2] , \out_i_vec_mult[0][1] , 
        \out_i_vec_mult[0][0] , \out_i_vec_mult[1][11] , 
        \out_i_vec_mult[1][10] , \out_i_vec_mult[1][9] , 
        \out_i_vec_mult[1][8] , \out_i_vec_mult[1][7] , \out_i_vec_mult[1][6] , 
        \out_i_vec_mult[1][5] , \out_i_vec_mult[1][4] , \out_i_vec_mult[1][3] , 
        \out_i_vec_mult[1][2] , \out_i_vec_mult[1][1] , \out_i_vec_mult[1][0] , 
        \out_i_vec_mult[2][11] , \out_i_vec_mult[2][10] , 
        \out_i_vec_mult[2][9] , \out_i_vec_mult[2][8] , \out_i_vec_mult[2][7] , 
        \out_i_vec_mult[2][6] , \out_i_vec_mult[2][5] , \out_i_vec_mult[2][4] , 
        \out_i_vec_mult[2][3] , \out_i_vec_mult[2][2] , \out_i_vec_mult[2][1] , 
        \out_i_vec_mult[2][0] , \out_i_vec_mult[3][11] , 
        \out_i_vec_mult[3][10] , \out_i_vec_mult[3][9] , 
        \out_i_vec_mult[3][8] , \out_i_vec_mult[3][7] , \out_i_vec_mult[3][6] , 
        \out_i_vec_mult[3][5] , \out_i_vec_mult[3][4] , \out_i_vec_mult[3][3] , 
        \out_i_vec_mult[3][2] , \out_i_vec_mult[3][1] , \out_i_vec_mult[3][0] }), .out_i_vec_sub({\out_i_vec_sub[0][11] , \out_i_vec_sub[0][10] , 
        \out_i_vec_sub[0][9] , \out_i_vec_sub[0][8] , \out_i_vec_sub[0][7] , 
        \out_i_vec_sub[0][6] , \out_i_vec_sub[0][5] , \out_i_vec_sub[0][4] , 
        \out_i_vec_sub[0][3] , \out_i_vec_sub[0][2] , \out_i_vec_sub[0][1] , 
        \out_i_vec_sub[0][0] , \out_i_vec_sub[1][11] , \out_i_vec_sub[1][10] , 
        \out_i_vec_sub[1][9] , \out_i_vec_sub[1][8] , \out_i_vec_sub[1][7] , 
        \out_i_vec_sub[1][6] , \out_i_vec_sub[1][5] , \out_i_vec_sub[1][4] , 
        \out_i_vec_sub[1][3] , \out_i_vec_sub[1][2] , \out_i_vec_sub[1][1] , 
        \out_i_vec_sub[1][0] , \out_i_vec_sub[2][11] , \out_i_vec_sub[2][10] , 
        \out_i_vec_sub[2][9] , \out_i_vec_sub[2][8] , \out_i_vec_sub[2][7] , 
        \out_i_vec_sub[2][6] , \out_i_vec_sub[2][5] , \out_i_vec_sub[2][4] , 
        \out_i_vec_sub[2][3] , \out_i_vec_sub[2][2] , \out_i_vec_sub[2][1] , 
        \out_i_vec_sub[2][0] , \out_i_vec_sub[3][11] , \out_i_vec_sub[3][10] , 
        \out_i_vec_sub[3][9] , \out_i_vec_sub[3][8] , \out_i_vec_sub[3][7] , 
        \out_i_vec_sub[3][6] , \out_i_vec_sub[3][5] , \out_i_vec_sub[3][4] , 
        \out_i_vec_sub[3][3] , \out_i_vec_sub[3][2] , \out_i_vec_sub[3][1] , 
        \out_i_vec_sub[3][0] }), .vec_in_i_AQ_mux({\vec_in_i_AQ_mux[0][11] , 
        \vec_in_i_AQ_mux[0][10] , \vec_in_i_AQ_mux[0][9] , 
        \vec_in_i_AQ_mux[0][8] , \vec_in_i_AQ_mux[0][7] , 
        \vec_in_i_AQ_mux[0][6] , \vec_in_i_AQ_mux[0][5] , 
        \vec_in_i_AQ_mux[0][4] , \vec_in_i_AQ_mux[0][3] , 
        \vec_in_i_AQ_mux[0][2] , \vec_in_i_AQ_mux[0][1] , 
        \vec_in_i_AQ_mux[0][0] , \vec_in_i_AQ_mux[1][11] , 
        \vec_in_i_AQ_mux[1][10] , \vec_in_i_AQ_mux[1][9] , 
        \vec_in_i_AQ_mux[1][8] , \vec_in_i_AQ_mux[1][7] , 
        \vec_in_i_AQ_mux[1][6] , \vec_in_i_AQ_mux[1][5] , 
        \vec_in_i_AQ_mux[1][4] , \vec_in_i_AQ_mux[1][3] , 
        \vec_in_i_AQ_mux[1][2] , \vec_in_i_AQ_mux[1][1] , 
        \vec_in_i_AQ_mux[1][0] , \vec_in_i_AQ_mux[2][11] , 
        \vec_in_i_AQ_mux[2][10] , \vec_in_i_AQ_mux[2][9] , 
        \vec_in_i_AQ_mux[2][8] , \vec_in_i_AQ_mux[2][7] , 
        \vec_in_i_AQ_mux[2][6] , \vec_in_i_AQ_mux[2][5] , 
        \vec_in_i_AQ_mux[2][4] , \vec_in_i_AQ_mux[2][3] , 
        \vec_in_i_AQ_mux[2][2] , \vec_in_i_AQ_mux[2][1] , 
        \vec_in_i_AQ_mux[2][0] , \vec_in_i_AQ_mux[3][11] , 
        \vec_in_i_AQ_mux[3][10] , \vec_in_i_AQ_mux[3][9] , 
        \vec_in_i_AQ_mux[3][8] , \vec_in_i_AQ_mux[3][7] , 
        \vec_in_i_AQ_mux[3][6] , \vec_in_i_AQ_mux[3][5] , 
        \vec_in_i_AQ_mux[3][4] , \vec_in_i_AQ_mux[3][3] , 
        \vec_in_i_AQ_mux[3][2] , \vec_in_i_AQ_mux[3][1] , 
        \vec_in_i_AQ_mux[3][0] }), .vec_in_AQ_sel(vec_in_AQ_sel), .col_sel_AQ(
        col_sel_AQ), .col_sel_AQ2_int(col_sel_AQ2_int), .col_sel_AQ2_mux(
        col_sel_AQ2_mux), .col_sel_AQ2_sel(col_sel_AQ2_sel), .wr_A(wr_A), 
        .wr_en_AQ_int(wr_en_AQ_int), .wr_en_AQ_mux(wr_en_AQ_mux), 
        .wr_en_AQ_sel(wr_en_AQ_sel), .out_mult(out_mult), .out_inner_prod_r(
        out_inner_prod_r), .single_in_r_R_mux(single_in_r_R_mux), 
        .out_inner_prod_i(out_inner_prod_i), .single_in_i_R_mux(
        single_in_i_R_mux), .single_in_R_sel(single_in_R_sel), .col_sel_R(
        col_sel_R), .col_sel_R_int(col_sel_R_int), .col_sel_R_mux(
        col_sel_R_mux), .col_sel_R_sel(col_sel_R_sel), .out_inv_sqrt(
        out_inv_sqrt), .in_b_r_vec_mult_mux(in_b_r_vec_mult_mux), 
        .in_b_i_vec_mult_mux(in_b_i_vec_mult_mux), .in_b_vec_mult_sel(
        in_b_vec_mult_sel), .w_col_sel_AQ_int(w_col_sel_AQ_int), 
        .w_col_sel_AQ_mux(w_col_sel_AQ_mux), .w_col_sel_AQ_sel(
        w_col_sel_AQ_sel), .vec_in_r_AQ_mux_0({\vec_in_r_AQ_mux[0][11] , 
        \vec_in_r_AQ_mux[0][10] , \vec_in_r_AQ_mux[0][9] , 
        \vec_in_r_AQ_mux[0][8] , \vec_in_r_AQ_mux[0][7] , 
        \vec_in_r_AQ_mux[0][6] , \vec_in_r_AQ_mux[0][5] , 
        \vec_in_r_AQ_mux[0][4] , \vec_in_r_AQ_mux[0][3] , 
        \vec_in_r_AQ_mux[0][2] , \vec_in_r_AQ_mux[0][1] , 
        \vec_in_r_AQ_mux[0][0] }), .single_out_r_AQ(single_out_r_AQ), 
        .vec_in_i_AQ_mux_0({\vec_in_i_AQ_mux[0][11] , \vec_in_i_AQ_mux[0][10] , 
        \vec_in_i_AQ_mux[0][9] , \vec_in_i_AQ_mux[0][8] , 
        \vec_in_i_AQ_mux[0][7] , \vec_in_i_AQ_mux[0][6] , 
        \vec_in_i_AQ_mux[0][5] , \vec_in_i_AQ_mux[0][4] , 
        \vec_in_i_AQ_mux[0][3] , \vec_in_i_AQ_mux[0][2] , 
        \vec_in_i_AQ_mux[0][1] , \vec_in_i_AQ_mux[0][0] }), .single_out_i_AQ(
        single_out_i_AQ), .in_a_r_inner_prod_mux(in_a_r_inner_prod_mux), 
        .in_a_i_inner_prod_mux(in_a_i_inner_prod_mux), .in_a_inner_prod_sel(
        in_a_inner_prod_sel), .out_r_vec_sub_0({\out_r_vec_sub[0][11] , 
        \out_r_vec_sub[0][10] , \out_r_vec_sub[0][9] , \out_r_vec_sub[0][8] , 
        \out_r_vec_sub[0][7] , \out_r_vec_sub[0][6] , \out_r_vec_sub[0][5] , 
        \out_r_vec_sub[0][4] , \out_r_vec_sub[0][3] , \out_r_vec_sub[0][2] , 
        \out_r_vec_sub[0][1] , \out_r_vec_sub[0][0] }), .single_out_r_AQ2(
        single_out_r_AQ2), .out_i_vec_sub_0({\out_i_vec_sub[0][11] , 
        \out_i_vec_sub[0][10] , \out_i_vec_sub[0][9] , \out_i_vec_sub[0][8] , 
        \out_i_vec_sub[0][7] , \out_i_vec_sub[0][6] , \out_i_vec_sub[0][5] , 
        \out_i_vec_sub[0][4] , \out_i_vec_sub[0][3] , \out_i_vec_sub[0][2] , 
        \out_i_vec_sub[0][1] , \out_i_vec_sub[0][0] }), .single_out_i_AQ2(
        single_out_i_AQ2), .in_b_r_inner_prod_mux(in_b_r_inner_prod_mux), 
        .in_b_i_inner_prod_mux(in_b_i_inner_prod_mux), .in_b_inner_prod_sel(
        in_b_inner_prod_sel) );
  qr_decomp_ctl_1 the_ctl ( .clk(clk), .rst(rst), .start(start), 
        .done_inner_prod(done_inner_prod), .done_inv_sqrt(done_inv_sqrt), 
        .out_inv_sqrt(out_inv_sqrt), .reduced_matrix(reduced_matrix), .done(
        done), .start_inner_prod(start_inner_prod), .start_inv_sqrt(
        start_inv_sqrt), .w_in_a_vec_sub(w_in_a_vec_sub), .row_sel_AQ2(
        row_sel_AQ2), .row_sel_R(row_sel_R), .wr_en_R(wr_en_R), 
        .row_sel_AQ_out(row_sel_AQ), .red_mat_reg_out(red_mat_reg), 
        .col_sel_AQ_int(col_sel_AQ_int), .col_sel_AQ2_int(col_sel_AQ2_int), 
        .in_a_r_mult(in_a_r_mult), .col_sel_R_int(col_sel_R_int), 
        .w_col_sel_AQ_int(w_col_sel_AQ_int), .wr_en_AQ_int(wr_en_AQ_int), 
        .vec_in_AQ_sel(vec_in_AQ_sel), .col_sel_AQ2_sel(col_sel_AQ2_sel), 
        .wr_en_AQ_sel(wr_en_AQ_sel), .col_sel_R_sel(col_sel_R_sel), 
        .w_col_sel_AQ_sel(w_col_sel_AQ_sel), .in_a_inner_prod_sel(
        in_a_inner_prod_sel), .in_b_inner_prod_sel(in_b_inner_prod_sel), 
        .single_in_R_sel(single_in_R_sel), .in_b_vec_mult_sel(
        in_b_vec_mult_sel) );
endmodule


module qr_wrapper_1 ( clk, rst, reduced_matrix, start, request_out, valid_out, 
        ready, .in_A_r({\in_A_r[0][11] , \in_A_r[0][10] , \in_A_r[0][9] , 
        \in_A_r[0][8] , \in_A_r[0][7] , \in_A_r[0][6] , \in_A_r[0][5] , 
        \in_A_r[0][4] , \in_A_r[0][3] , \in_A_r[0][2] , \in_A_r[0][1] , 
        \in_A_r[0][0] , \in_A_r[1][11] , \in_A_r[1][10] , \in_A_r[1][9] , 
        \in_A_r[1][8] , \in_A_r[1][7] , \in_A_r[1][6] , \in_A_r[1][5] , 
        \in_A_r[1][4] , \in_A_r[1][3] , \in_A_r[1][2] , \in_A_r[1][1] , 
        \in_A_r[1][0] , \in_A_r[2][11] , \in_A_r[2][10] , \in_A_r[2][9] , 
        \in_A_r[2][8] , \in_A_r[2][7] , \in_A_r[2][6] , \in_A_r[2][5] , 
        \in_A_r[2][4] , \in_A_r[2][3] , \in_A_r[2][2] , \in_A_r[2][1] , 
        \in_A_r[2][0] , \in_A_r[3][11] , \in_A_r[3][10] , \in_A_r[3][9] , 
        \in_A_r[3][8] , \in_A_r[3][7] , \in_A_r[3][6] , \in_A_r[3][5] , 
        \in_A_r[3][4] , \in_A_r[3][3] , \in_A_r[3][2] , \in_A_r[3][1] , 
        \in_A_r[3][0] }), .in_A_i({\in_A_i[0][11] , \in_A_i[0][10] , 
        \in_A_i[0][9] , \in_A_i[0][8] , \in_A_i[0][7] , \in_A_i[0][6] , 
        \in_A_i[0][5] , \in_A_i[0][4] , \in_A_i[0][3] , \in_A_i[0][2] , 
        \in_A_i[0][1] , \in_A_i[0][0] , \in_A_i[1][11] , \in_A_i[1][10] , 
        \in_A_i[1][9] , \in_A_i[1][8] , \in_A_i[1][7] , \in_A_i[1][6] , 
        \in_A_i[1][5] , \in_A_i[1][4] , \in_A_i[1][3] , \in_A_i[1][2] , 
        \in_A_i[1][1] , \in_A_i[1][0] , \in_A_i[2][11] , \in_A_i[2][10] , 
        \in_A_i[2][9] , \in_A_i[2][8] , \in_A_i[2][7] , \in_A_i[2][6] , 
        \in_A_i[2][5] , \in_A_i[2][4] , \in_A_i[2][3] , \in_A_i[2][2] , 
        \in_A_i[2][1] , \in_A_i[2][0] , \in_A_i[3][11] , \in_A_i[3][10] , 
        \in_A_i[3][9] , \in_A_i[3][8] , \in_A_i[3][7] , \in_A_i[3][6] , 
        \in_A_i[3][5] , \in_A_i[3][4] , \in_A_i[3][3] , \in_A_i[3][2] , 
        \in_A_i[3][1] , \in_A_i[3][0] }), .out_Q_r({\out_Q_r[0][11] , 
        \out_Q_r[0][10] , \out_Q_r[0][9] , \out_Q_r[0][8] , \out_Q_r[0][7] , 
        \out_Q_r[0][6] , \out_Q_r[0][5] , \out_Q_r[0][4] , \out_Q_r[0][3] , 
        \out_Q_r[0][2] , \out_Q_r[0][1] , \out_Q_r[0][0] , \out_Q_r[1][11] , 
        \out_Q_r[1][10] , \out_Q_r[1][9] , \out_Q_r[1][8] , \out_Q_r[1][7] , 
        \out_Q_r[1][6] , \out_Q_r[1][5] , \out_Q_r[1][4] , \out_Q_r[1][3] , 
        \out_Q_r[1][2] , \out_Q_r[1][1] , \out_Q_r[1][0] , \out_Q_r[2][11] , 
        \out_Q_r[2][10] , \out_Q_r[2][9] , \out_Q_r[2][8] , \out_Q_r[2][7] , 
        \out_Q_r[2][6] , \out_Q_r[2][5] , \out_Q_r[2][4] , \out_Q_r[2][3] , 
        \out_Q_r[2][2] , \out_Q_r[2][1] , \out_Q_r[2][0] , \out_Q_r[3][11] , 
        \out_Q_r[3][10] , \out_Q_r[3][9] , \out_Q_r[3][8] , \out_Q_r[3][7] , 
        \out_Q_r[3][6] , \out_Q_r[3][5] , \out_Q_r[3][4] , \out_Q_r[3][3] , 
        \out_Q_r[3][2] , \out_Q_r[3][1] , \out_Q_r[3][0] }), .out_Q_i({
        \out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] , \out_Q_i[0][8] , 
        \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] , \out_Q_i[0][4] , 
        \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] , \out_Q_i[0][0] , 
        \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] , \out_Q_i[1][8] , 
        \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] , \out_Q_i[1][4] , 
        \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] , \out_Q_i[1][0] , 
        \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] , \out_Q_i[2][8] , 
        \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] , \out_Q_i[2][4] , 
        \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] , \out_Q_i[2][0] , 
        \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] , \out_Q_i[3][8] , 
        \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] , \out_Q_i[3][4] , 
        \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] , \out_Q_i[3][0] }), 
    .out_R_r({\out_R_r[0][11] , \out_R_r[0][10] , \out_R_r[0][9] , 
        \out_R_r[0][8] , \out_R_r[0][7] , \out_R_r[0][6] , \out_R_r[0][5] , 
        \out_R_r[0][4] , \out_R_r[0][3] , \out_R_r[0][2] , \out_R_r[0][1] , 
        \out_R_r[0][0] , \out_R_r[1][11] , \out_R_r[1][10] , \out_R_r[1][9] , 
        \out_R_r[1][8] , \out_R_r[1][7] , \out_R_r[1][6] , \out_R_r[1][5] , 
        \out_R_r[1][4] , \out_R_r[1][3] , \out_R_r[1][2] , \out_R_r[1][1] , 
        \out_R_r[1][0] , \out_R_r[2][11] , \out_R_r[2][10] , \out_R_r[2][9] , 
        \out_R_r[2][8] , \out_R_r[2][7] , \out_R_r[2][6] , \out_R_r[2][5] , 
        \out_R_r[2][4] , \out_R_r[2][3] , \out_R_r[2][2] , \out_R_r[2][1] , 
        \out_R_r[2][0] , \out_R_r[3][11] , \out_R_r[3][10] , \out_R_r[3][9] , 
        \out_R_r[3][8] , \out_R_r[3][7] , \out_R_r[3][6] , \out_R_r[3][5] , 
        \out_R_r[3][4] , \out_R_r[3][3] , \out_R_r[3][2] , \out_R_r[3][1] , 
        \out_R_r[3][0] }), .out_R_i({\out_R_i[0][11] , \out_R_i[0][10] , 
        \out_R_i[0][9] , \out_R_i[0][8] , \out_R_i[0][7] , \out_R_i[0][6] , 
        \out_R_i[0][5] , \out_R_i[0][4] , \out_R_i[0][3] , \out_R_i[0][2] , 
        \out_R_i[0][1] , \out_R_i[0][0] , \out_R_i[1][11] , \out_R_i[1][10] , 
        \out_R_i[1][9] , \out_R_i[1][8] , \out_R_i[1][7] , \out_R_i[1][6] , 
        \out_R_i[1][5] , \out_R_i[1][4] , \out_R_i[1][3] , \out_R_i[1][2] , 
        \out_R_i[1][1] , \out_R_i[1][0] , \out_R_i[2][11] , \out_R_i[2][10] , 
        \out_R_i[2][9] , \out_R_i[2][8] , \out_R_i[2][7] , \out_R_i[2][6] , 
        \out_R_i[2][5] , \out_R_i[2][4] , \out_R_i[2][3] , \out_R_i[2][2] , 
        \out_R_i[2][1] , \out_R_i[2][0] , \out_R_i[3][11] , \out_R_i[3][10] , 
        \out_R_i[3][9] , \out_R_i[3][8] , \out_R_i[3][7] , \out_R_i[3][6] , 
        \out_R_i[3][5] , \out_R_i[3][4] , \out_R_i[3][3] , \out_R_i[3][2] , 
        \out_R_i[3][1] , \out_R_i[3][0] }) );
  input clk, rst, reduced_matrix, start, request_out, \in_A_r[0][11] ,
         \in_A_r[0][10] , \in_A_r[0][9] , \in_A_r[0][8] , \in_A_r[0][7] ,
         \in_A_r[0][6] , \in_A_r[0][5] , \in_A_r[0][4] , \in_A_r[0][3] ,
         \in_A_r[0][2] , \in_A_r[0][1] , \in_A_r[0][0] , \in_A_r[1][11] ,
         \in_A_r[1][10] , \in_A_r[1][9] , \in_A_r[1][8] , \in_A_r[1][7] ,
         \in_A_r[1][6] , \in_A_r[1][5] , \in_A_r[1][4] , \in_A_r[1][3] ,
         \in_A_r[1][2] , \in_A_r[1][1] , \in_A_r[1][0] , \in_A_r[2][11] ,
         \in_A_r[2][10] , \in_A_r[2][9] , \in_A_r[2][8] , \in_A_r[2][7] ,
         \in_A_r[2][6] , \in_A_r[2][5] , \in_A_r[2][4] , \in_A_r[2][3] ,
         \in_A_r[2][2] , \in_A_r[2][1] , \in_A_r[2][0] , \in_A_r[3][11] ,
         \in_A_r[3][10] , \in_A_r[3][9] , \in_A_r[3][8] , \in_A_r[3][7] ,
         \in_A_r[3][6] , \in_A_r[3][5] , \in_A_r[3][4] , \in_A_r[3][3] ,
         \in_A_r[3][2] , \in_A_r[3][1] , \in_A_r[3][0] , \in_A_i[0][11] ,
         \in_A_i[0][10] , \in_A_i[0][9] , \in_A_i[0][8] , \in_A_i[0][7] ,
         \in_A_i[0][6] , \in_A_i[0][5] , \in_A_i[0][4] , \in_A_i[0][3] ,
         \in_A_i[0][2] , \in_A_i[0][1] , \in_A_i[0][0] , \in_A_i[1][11] ,
         \in_A_i[1][10] , \in_A_i[1][9] , \in_A_i[1][8] , \in_A_i[1][7] ,
         \in_A_i[1][6] , \in_A_i[1][5] , \in_A_i[1][4] , \in_A_i[1][3] ,
         \in_A_i[1][2] , \in_A_i[1][1] , \in_A_i[1][0] , \in_A_i[2][11] ,
         \in_A_i[2][10] , \in_A_i[2][9] , \in_A_i[2][8] , \in_A_i[2][7] ,
         \in_A_i[2][6] , \in_A_i[2][5] , \in_A_i[2][4] , \in_A_i[2][3] ,
         \in_A_i[2][2] , \in_A_i[2][1] , \in_A_i[2][0] , \in_A_i[3][11] ,
         \in_A_i[3][10] , \in_A_i[3][9] , \in_A_i[3][8] , \in_A_i[3][7] ,
         \in_A_i[3][6] , \in_A_i[3][5] , \in_A_i[3][4] , \in_A_i[3][3] ,
         \in_A_i[3][2] , \in_A_i[3][1] , \in_A_i[3][0] ;
  output valid_out, ready, \out_Q_r[0][11] , \out_Q_r[0][10] , \out_Q_r[0][9] ,
         \out_Q_r[0][8] , \out_Q_r[0][7] , \out_Q_r[0][6] , \out_Q_r[0][5] ,
         \out_Q_r[0][4] , \out_Q_r[0][3] , \out_Q_r[0][2] , \out_Q_r[0][1] ,
         \out_Q_r[0][0] , \out_Q_r[1][11] , \out_Q_r[1][10] , \out_Q_r[1][9] ,
         \out_Q_r[1][8] , \out_Q_r[1][7] , \out_Q_r[1][6] , \out_Q_r[1][5] ,
         \out_Q_r[1][4] , \out_Q_r[1][3] , \out_Q_r[1][2] , \out_Q_r[1][1] ,
         \out_Q_r[1][0] , \out_Q_r[2][11] , \out_Q_r[2][10] , \out_Q_r[2][9] ,
         \out_Q_r[2][8] , \out_Q_r[2][7] , \out_Q_r[2][6] , \out_Q_r[2][5] ,
         \out_Q_r[2][4] , \out_Q_r[2][3] , \out_Q_r[2][2] , \out_Q_r[2][1] ,
         \out_Q_r[2][0] , \out_Q_r[3][11] , \out_Q_r[3][10] , \out_Q_r[3][9] ,
         \out_Q_r[3][8] , \out_Q_r[3][7] , \out_Q_r[3][6] , \out_Q_r[3][5] ,
         \out_Q_r[3][4] , \out_Q_r[3][3] , \out_Q_r[3][2] , \out_Q_r[3][1] ,
         \out_Q_r[3][0] , \out_Q_i[0][11] , \out_Q_i[0][10] , \out_Q_i[0][9] ,
         \out_Q_i[0][8] , \out_Q_i[0][7] , \out_Q_i[0][6] , \out_Q_i[0][5] ,
         \out_Q_i[0][4] , \out_Q_i[0][3] , \out_Q_i[0][2] , \out_Q_i[0][1] ,
         \out_Q_i[0][0] , \out_Q_i[1][11] , \out_Q_i[1][10] , \out_Q_i[1][9] ,
         \out_Q_i[1][8] , \out_Q_i[1][7] , \out_Q_i[1][6] , \out_Q_i[1][5] ,
         \out_Q_i[1][4] , \out_Q_i[1][3] , \out_Q_i[1][2] , \out_Q_i[1][1] ,
         \out_Q_i[1][0] , \out_Q_i[2][11] , \out_Q_i[2][10] , \out_Q_i[2][9] ,
         \out_Q_i[2][8] , \out_Q_i[2][7] , \out_Q_i[2][6] , \out_Q_i[2][5] ,
         \out_Q_i[2][4] , \out_Q_i[2][3] , \out_Q_i[2][2] , \out_Q_i[2][1] ,
         \out_Q_i[2][0] , \out_Q_i[3][11] , \out_Q_i[3][10] , \out_Q_i[3][9] ,
         \out_Q_i[3][8] , \out_Q_i[3][7] , \out_Q_i[3][6] , \out_Q_i[3][5] ,
         \out_Q_i[3][4] , \out_Q_i[3][3] , \out_Q_i[3][2] , \out_Q_i[3][1] ,
         \out_Q_i[3][0] , \out_R_r[0][11] , \out_R_r[0][10] , \out_R_r[0][9] ,
         \out_R_r[0][8] , \out_R_r[0][7] , \out_R_r[0][6] , \out_R_r[0][5] ,
         \out_R_r[0][4] , \out_R_r[0][3] , \out_R_r[0][2] , \out_R_r[0][1] ,
         \out_R_r[0][0] , \out_R_r[1][11] , \out_R_r[1][10] , \out_R_r[1][9] ,
         \out_R_r[1][8] , \out_R_r[1][7] , \out_R_r[1][6] , \out_R_r[1][5] ,
         \out_R_r[1][4] , \out_R_r[1][3] , \out_R_r[1][2] , \out_R_r[1][1] ,
         \out_R_r[1][0] , \out_R_r[2][11] , \out_R_r[2][10] , \out_R_r[2][9] ,
         \out_R_r[2][8] , \out_R_r[2][7] , \out_R_r[2][6] , \out_R_r[2][5] ,
         \out_R_r[2][4] , \out_R_r[2][3] , \out_R_r[2][2] , \out_R_r[2][1] ,
         \out_R_r[2][0] , \out_R_r[3][11] , \out_R_r[3][10] , \out_R_r[3][9] ,
         \out_R_r[3][8] , \out_R_r[3][7] , \out_R_r[3][6] , \out_R_r[3][5] ,
         \out_R_r[3][4] , \out_R_r[3][3] , \out_R_r[3][2] , \out_R_r[3][1] ,
         \out_R_r[3][0] , \out_R_i[0][11] , \out_R_i[0][10] , \out_R_i[0][9] ,
         \out_R_i[0][8] , \out_R_i[0][7] , \out_R_i[0][6] , \out_R_i[0][5] ,
         \out_R_i[0][4] , \out_R_i[0][3] , \out_R_i[0][2] , \out_R_i[0][1] ,
         \out_R_i[0][0] , \out_R_i[1][11] , \out_R_i[1][10] , \out_R_i[1][9] ,
         \out_R_i[1][8] , \out_R_i[1][7] , \out_R_i[1][6] , \out_R_i[1][5] ,
         \out_R_i[1][4] , \out_R_i[1][3] , \out_R_i[1][2] , \out_R_i[1][1] ,
         \out_R_i[1][0] , \out_R_i[2][11] , \out_R_i[2][10] , \out_R_i[2][9] ,
         \out_R_i[2][8] , \out_R_i[2][7] , \out_R_i[2][6] , \out_R_i[2][5] ,
         \out_R_i[2][4] , \out_R_i[2][3] , \out_R_i[2][2] , \out_R_i[2][1] ,
         \out_R_i[2][0] , \out_R_i[3][11] , \out_R_i[3][10] , \out_R_i[3][9] ,
         \out_R_i[3][8] , \out_R_i[3][7] , \out_R_i[3][6] , \out_R_i[3][5] ,
         \out_R_i[3][4] , \out_R_i[3][3] , \out_R_i[3][2] , \out_R_i[3][1] ,
         \out_R_i[3][0] ;
  wire   wr_A_QR, red_mat_reg, start_QR, done_QR, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n19, n21, n23, n24, n25, n26, n27, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n12,
         n14, n15, n16, n17, n18, n20, n22, n28;
  wire   [1:0] col_sel_AQ;
  wire   [1:0] col_sel_R;
  wire   [1:0] state;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;
  assign \out_R_i[3][11]  = 1'b0;
  assign \out_R_i[3][10]  = 1'b0;
  assign \out_R_i[3][9]  = 1'b0;
  assign \out_R_i[3][8]  = 1'b0;
  assign \out_R_i[3][7]  = 1'b0;
  assign \out_R_i[3][6]  = 1'b0;
  assign \out_R_i[3][5]  = 1'b0;
  assign \out_R_i[3][4]  = 1'b0;
  assign \out_R_i[3][3]  = 1'b0;
  assign \out_R_i[3][2]  = 1'b0;
  assign \out_R_i[3][1]  = 1'b0;
  assign \out_R_i[3][0]  = 1'b0;

  DFFARX1 \col_sel_AQ_reg[0]  ( .D(n58), .CLK(clk), .RSTB(n11), .Q(
        col_sel_AQ[0]), .QN(n21) );
  DFFARX1 wr_A_QR_reg ( .D(n52), .CLK(clk), .RSTB(n10), .Q(wr_A_QR) );
  DFFARX1 \state_reg[0]  ( .D(n55), .CLK(clk), .RSTB(n9), .Q(state[0]) );
  DFFARX1 \state_reg[1]  ( .D(n56), .CLK(clk), .RSTB(n8), .Q(state[1]), .QN(
        n19) );
  DFFARX1 start_QR_reg ( .D(n50), .CLK(clk), .RSTB(n7), .Q(start_QR) );
  DFFARX1 \col_sel_AQ_reg[1]  ( .D(n57), .CLK(clk), .RSTB(n6), .Q(
        col_sel_AQ[1]) );
  DFFARX1 \col_sel_R_reg[0]  ( .D(n49), .CLK(clk), .RSTB(n5), .Q(col_sel_R[0])
         );
  DFFARX1 \col_sel_R_reg[1]  ( .D(n48), .CLK(clk), .RSTB(n4), .Q(col_sel_R[1])
         );
  DFFARX1 red_mat_reg_reg ( .D(n53), .CLK(clk), .RSTB(n3), .Q(red_mat_reg) );
  DFFARX1 ready_reg ( .D(n54), .CLK(clk), .RSTB(n2), .Q(ready) );
  DFFARX1 valid_out_reg ( .D(n51), .CLK(clk), .RSTB(n1), .Q(valid_out) );
  AO22X1 U35 ( .IN1(col_sel_R[1]), .IN2(n23), .IN3(n24), .IN4(col_sel_R[0]), 
        .Q(n48) );
  AO21X1 U36 ( .IN1(n26), .IN2(n25), .IN3(n27), .Q(n23) );
  AO22X1 U38 ( .IN1(n29), .IN2(n30), .IN3(start_QR), .IN4(n16), .Q(n50) );
  AO21X1 U39 ( .IN1(n31), .IN2(n29), .IN3(n32), .Q(n30) );
  AO22X1 U40 ( .IN1(n22), .IN2(n25), .IN3(valid_out), .IN4(n33), .Q(n51) );
  NAND3X0 U41 ( .IN1(n34), .IN2(n28), .IN3(request_out), .QN(n26) );
  AO22X1 U42 ( .IN1(n35), .IN2(n36), .IN3(wr_A_QR), .IN4(n15), .Q(n52) );
  NAND4X0 U43 ( .IN1(reduced_matrix), .IN2(start), .IN3(n34), .IN4(n25), .QN(
        n38) );
  OAI21X1 U44 ( .IN1(n39), .IN2(n28), .IN3(red_mat_reg), .QN(n37) );
  AO21X1 U45 ( .IN1(ready), .IN2(n39), .IN3(n40), .Q(n54) );
  NOR4X0 U46 ( .IN1(start), .IN2(request_out), .IN3(n18), .IN4(n20), .QN(n40)
         );
  AO22X1 U47 ( .IN1(n35), .IN2(n41), .IN3(n14), .IN4(state[0]), .Q(n55) );
  AO22X1 U48 ( .IN1(n14), .IN2(state[1]), .IN3(n42), .IN4(n41), .Q(n56) );
  AO21X1 U49 ( .IN1(n35), .IN2(n28), .IN3(n29), .Q(n42) );
  AO221X1 U50 ( .IN1(done_QR), .IN2(n32), .IN3(n35), .IN4(request_out), .IN5(
        n43), .Q(n41) );
  AO21X1 U51 ( .IN1(n31), .IN2(n18), .IN3(n36), .Q(n43) );
  AO22X1 U52 ( .IN1(n31), .IN2(n29), .IN3(start), .IN4(n35), .Q(n36) );
  AO22X1 U53 ( .IN1(n44), .IN2(col_sel_AQ[1]), .IN3(n45), .IN4(n17), .Q(n57)
         );
  XNOR2X1 U54 ( .IN1(col_sel_AQ[1]), .IN2(n21), .Q(n45) );
  AO22X1 U55 ( .IN1(n44), .IN2(col_sel_AQ[0]), .IN3(n17), .IN4(n21), .Q(n58)
         );
  AND2X1 U56 ( .IN1(n46), .IN2(n47), .Q(n44) );
  OAI21X1 U57 ( .IN1(start), .IN2(request_out), .IN3(n35), .QN(n47) );
  AND2X1 U58 ( .IN1(state[0]), .IN2(n19), .Q(n29) );
  qr_decomp_USE_NEWTON1 qr_decomp_inst ( .in_A_r({\in_A_r[0][11] , 
        \in_A_r[0][10] , \in_A_r[0][9] , \in_A_r[0][8] , \in_A_r[0][7] , 
        \in_A_r[0][6] , \in_A_r[0][5] , \in_A_r[0][4] , \in_A_r[0][3] , 
        \in_A_r[0][2] , \in_A_r[0][1] , \in_A_r[0][0] , \in_A_r[1][11] , 
        \in_A_r[1][10] , \in_A_r[1][9] , \in_A_r[1][8] , \in_A_r[1][7] , 
        \in_A_r[1][6] , \in_A_r[1][5] , \in_A_r[1][4] , \in_A_r[1][3] , 
        \in_A_r[1][2] , \in_A_r[1][1] , \in_A_r[1][0] , \in_A_r[2][11] , 
        \in_A_r[2][10] , \in_A_r[2][9] , \in_A_r[2][8] , \in_A_r[2][7] , 
        \in_A_r[2][6] , \in_A_r[2][5] , \in_A_r[2][4] , \in_A_r[2][3] , 
        \in_A_r[2][2] , \in_A_r[2][1] , \in_A_r[2][0] , \in_A_r[3][11] , 
        \in_A_r[3][10] , \in_A_r[3][9] , \in_A_r[3][8] , \in_A_r[3][7] , 
        \in_A_r[3][6] , \in_A_r[3][5] , \in_A_r[3][4] , \in_A_r[3][3] , 
        \in_A_r[3][2] , \in_A_r[3][1] , \in_A_r[3][0] }), .in_A_i({
        \in_A_i[0][11] , \in_A_i[0][10] , \in_A_i[0][9] , \in_A_i[0][8] , 
        \in_A_i[0][7] , \in_A_i[0][6] , \in_A_i[0][5] , \in_A_i[0][4] , 
        \in_A_i[0][3] , \in_A_i[0][2] , \in_A_i[0][1] , \in_A_i[0][0] , 
        \in_A_i[1][11] , \in_A_i[1][10] , \in_A_i[1][9] , \in_A_i[1][8] , 
        \in_A_i[1][7] , \in_A_i[1][6] , \in_A_i[1][5] , \in_A_i[1][4] , 
        \in_A_i[1][3] , \in_A_i[1][2] , \in_A_i[1][1] , \in_A_i[1][0] , 
        \in_A_i[2][11] , \in_A_i[2][10] , \in_A_i[2][9] , \in_A_i[2][8] , 
        \in_A_i[2][7] , \in_A_i[2][6] , \in_A_i[2][5] , \in_A_i[2][4] , 
        \in_A_i[2][3] , \in_A_i[2][2] , \in_A_i[2][1] , \in_A_i[2][0] , 
        \in_A_i[3][11] , \in_A_i[3][10] , \in_A_i[3][9] , \in_A_i[3][8] , 
        \in_A_i[3][7] , \in_A_i[3][6] , \in_A_i[3][5] , \in_A_i[3][4] , 
        \in_A_i[3][3] , \in_A_i[3][2] , \in_A_i[3][1] , \in_A_i[3][0] }), 
        .out_Q_r({\out_Q_r[0][11] , \out_Q_r[0][10] , \out_Q_r[0][9] , 
        \out_Q_r[0][8] , \out_Q_r[0][7] , \out_Q_r[0][6] , \out_Q_r[0][5] , 
        \out_Q_r[0][4] , \out_Q_r[0][3] , \out_Q_r[0][2] , \out_Q_r[0][1] , 
        \out_Q_r[0][0] , \out_Q_r[1][11] , \out_Q_r[1][10] , \out_Q_r[1][9] , 
        \out_Q_r[1][8] , \out_Q_r[1][7] , \out_Q_r[1][6] , \out_Q_r[1][5] , 
        \out_Q_r[1][4] , \out_Q_r[1][3] , \out_Q_r[1][2] , \out_Q_r[1][1] , 
        \out_Q_r[1][0] , \out_Q_r[2][11] , \out_Q_r[2][10] , \out_Q_r[2][9] , 
        \out_Q_r[2][8] , \out_Q_r[2][7] , \out_Q_r[2][6] , \out_Q_r[2][5] , 
        \out_Q_r[2][4] , \out_Q_r[2][3] , \out_Q_r[2][2] , \out_Q_r[2][1] , 
        \out_Q_r[2][0] , \out_Q_r[3][11] , \out_Q_r[3][10] , \out_Q_r[3][9] , 
        \out_Q_r[3][8] , \out_Q_r[3][7] , \out_Q_r[3][6] , \out_Q_r[3][5] , 
        \out_Q_r[3][4] , \out_Q_r[3][3] , \out_Q_r[3][2] , \out_Q_r[3][1] , 
        \out_Q_r[3][0] }), .out_Q_i({\out_Q_i[0][11] , \out_Q_i[0][10] , 
        \out_Q_i[0][9] , \out_Q_i[0][8] , \out_Q_i[0][7] , \out_Q_i[0][6] , 
        \out_Q_i[0][5] , \out_Q_i[0][4] , \out_Q_i[0][3] , \out_Q_i[0][2] , 
        \out_Q_i[0][1] , \out_Q_i[0][0] , \out_Q_i[1][11] , \out_Q_i[1][10] , 
        \out_Q_i[1][9] , \out_Q_i[1][8] , \out_Q_i[1][7] , \out_Q_i[1][6] , 
        \out_Q_i[1][5] , \out_Q_i[1][4] , \out_Q_i[1][3] , \out_Q_i[1][2] , 
        \out_Q_i[1][1] , \out_Q_i[1][0] , \out_Q_i[2][11] , \out_Q_i[2][10] , 
        \out_Q_i[2][9] , \out_Q_i[2][8] , \out_Q_i[2][7] , \out_Q_i[2][6] , 
        \out_Q_i[2][5] , \out_Q_i[2][4] , \out_Q_i[2][3] , \out_Q_i[2][2] , 
        \out_Q_i[2][1] , \out_Q_i[2][0] , \out_Q_i[3][11] , \out_Q_i[3][10] , 
        \out_Q_i[3][9] , \out_Q_i[3][8] , \out_Q_i[3][7] , \out_Q_i[3][6] , 
        \out_Q_i[3][5] , \out_Q_i[3][4] , \out_Q_i[3][3] , \out_Q_i[3][2] , 
        \out_Q_i[3][1] , \out_Q_i[3][0] }), .out_R_r({\out_R_r[0][11] , 
        \out_R_r[0][10] , \out_R_r[0][9] , \out_R_r[0][8] , \out_R_r[0][7] , 
        \out_R_r[0][6] , \out_R_r[0][5] , \out_R_r[0][4] , \out_R_r[0][3] , 
        \out_R_r[0][2] , \out_R_r[0][1] , \out_R_r[0][0] , \out_R_r[1][11] , 
        \out_R_r[1][10] , \out_R_r[1][9] , \out_R_r[1][8] , \out_R_r[1][7] , 
        \out_R_r[1][6] , \out_R_r[1][5] , \out_R_r[1][4] , \out_R_r[1][3] , 
        \out_R_r[1][2] , \out_R_r[1][1] , \out_R_r[1][0] , \out_R_r[2][11] , 
        \out_R_r[2][10] , \out_R_r[2][9] , \out_R_r[2][8] , \out_R_r[2][7] , 
        \out_R_r[2][6] , \out_R_r[2][5] , \out_R_r[2][4] , \out_R_r[2][3] , 
        \out_R_r[2][2] , \out_R_r[2][1] , \out_R_r[2][0] , \out_R_r[3][11] , 
        \out_R_r[3][10] , \out_R_r[3][9] , \out_R_r[3][8] , \out_R_r[3][7] , 
        \out_R_r[3][6] , \out_R_r[3][5] , \out_R_r[3][4] , \out_R_r[3][3] , 
        \out_R_r[3][2] , \out_R_r[3][1] , \out_R_r[3][0] }), .out_R_i({
        \out_R_i[0][11] , \out_R_i[0][10] , \out_R_i[0][9] , \out_R_i[0][8] , 
        \out_R_i[0][7] , \out_R_i[0][6] , \out_R_i[0][5] , \out_R_i[0][4] , 
        \out_R_i[0][3] , \out_R_i[0][2] , \out_R_i[0][1] , \out_R_i[0][0] , 
        \out_R_i[1][11] , \out_R_i[1][10] , \out_R_i[1][9] , \out_R_i[1][8] , 
        \out_R_i[1][7] , \out_R_i[1][6] , \out_R_i[1][5] , \out_R_i[1][4] , 
        \out_R_i[1][3] , \out_R_i[1][2] , \out_R_i[1][1] , \out_R_i[1][0] , 
        \out_R_i[2][11] , \out_R_i[2][10] , \out_R_i[2][9] , \out_R_i[2][8] , 
        \out_R_i[2][7] , \out_R_i[2][6] , \out_R_i[2][5] , \out_R_i[2][4] , 
        \out_R_i[2][3] , \out_R_i[2][2] , \out_R_i[2][1] , \out_R_i[2][0] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}), .wr_A(wr_A_QR), 
        .col_sel_AQ(col_sel_AQ), .col_sel_R(col_sel_R), .reduced_matrix(
        red_mat_reg), .clk(clk), .rst(rst), .start(start_QR), .done(done_QR)
         );
  INVX0 U3 ( .INP(n46), .ZN(n17) );
  NOR2X0 U4 ( .IN1(n29), .IN2(n32), .QN(n34) );
  NAND2X0 U5 ( .IN1(n34), .IN2(n25), .QN(n39) );
  INVX0 U6 ( .INP(n25), .ZN(n18) );
  NOR2X0 U7 ( .IN1(n18), .IN2(n29), .QN(n46) );
  INVX0 U8 ( .INP(n41), .ZN(n14) );
  NOR2X0 U9 ( .IN1(n19), .IN2(state[0]), .QN(n32) );
  NAND2X0 U10 ( .IN1(n37), .IN2(n38), .QN(n53) );
  INVX0 U11 ( .INP(n34), .ZN(n20) );
  NAND2X0 U12 ( .IN1(state[1]), .IN2(state[0]), .QN(n25) );
  NOR2X0 U13 ( .IN1(n25), .IN2(col_sel_R[0]), .QN(n27) );
  OR2X1 U14 ( .IN1(n27), .IN2(n12), .Q(n49) );
  AND3X1 U15 ( .IN1(n26), .IN2(n25), .IN3(col_sel_R[0]), .Q(n12) );
  NAND2X0 U16 ( .IN1(n31), .IN2(n18), .QN(n33) );
  INVX0 U17 ( .INP(n26), .ZN(n22) );
  NOR2X0 U18 ( .IN1(state[0]), .IN2(state[1]), .QN(n35) );
  NOR2X0 U19 ( .IN1(col_sel_R[1]), .IN2(n25), .QN(n24) );
  OA21X1 U20 ( .IN1(red_mat_reg), .IN2(col_sel_AQ[1]), .IN3(col_sel_AQ[0]), 
        .Q(n31) );
  INVX0 U21 ( .INP(n30), .ZN(n16) );
  INVX0 U22 ( .INP(n36), .ZN(n15) );
  INVX0 U23 ( .INP(start), .ZN(n28) );
  INVX0 U24 ( .INP(rst), .ZN(n1) );
  INVX0 U25 ( .INP(rst), .ZN(n2) );
  INVX0 U26 ( .INP(rst), .ZN(n3) );
  INVX0 U27 ( .INP(rst), .ZN(n4) );
  INVX0 U28 ( .INP(rst), .ZN(n5) );
  INVX0 U29 ( .INP(rst), .ZN(n6) );
  INVX0 U30 ( .INP(rst), .ZN(n7) );
  INVX0 U31 ( .INP(rst), .ZN(n8) );
  INVX0 U32 ( .INP(rst), .ZN(n9) );
  INVX0 U33 ( .INP(rst), .ZN(n10) );
  INVX0 U34 ( .INP(rst), .ZN(n11) );
endmodule


module qr_wrapper_wrapper ( CLK, RST, REDUCED0MATRIX, START, REQUEST0OUT, 
        VALID0OUT, READY, IN0A0R, IN0A0I, SIGMA0IN, OUT0Q0R, OUT0Q0I, OUT0R0R, 
        OUT0R0I, PERMUT );
  input [47:0] IN0A0R;
  input [47:0] IN0A0I;
  input [11:0] SIGMA0IN;
  output [47:0] OUT0Q0R;
  output [47:0] OUT0Q0I;
  output [47:0] OUT0R0R;
  output [47:0] OUT0R0I;
  output [7:0] PERMUT;
  input CLK, RST, REDUCED0MATRIX, START, REQUEST0OUT;
  output VALID0OUT, READY;

  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11;
  assign PERMUT[0] = 1'b0;
  assign PERMUT[1] = 1'b0;
  assign PERMUT[2] = 1'b0;
  assign PERMUT[3] = 1'b0;
  assign PERMUT[4] = 1'b0;
  assign PERMUT[5] = 1'b0;
  assign PERMUT[6] = 1'b0;
  assign PERMUT[7] = 1'b0;
  assign OUT0R0I[11] = 1'b0;
  assign OUT0R0I[10] = 1'b0;
  assign OUT0R0I[9] = 1'b0;
  assign OUT0R0I[8] = 1'b0;
  assign OUT0R0I[7] = 1'b0;
  assign OUT0R0I[6] = 1'b0;
  assign OUT0R0I[5] = 1'b0;
  assign OUT0R0I[4] = 1'b0;
  assign OUT0R0I[3] = 1'b0;
  assign OUT0R0I[2] = 1'b0;
  assign OUT0R0I[1] = 1'b0;
  assign OUT0R0I[0] = 1'b0;

  qr_wrapper_1 QR0WRAPPER0INST ( .clk(CLK), .rst(RST), .reduced_matrix(
        REDUCED0MATRIX), .start(START), .request_out(REQUEST0OUT), .valid_out(
        VALID0OUT), .ready(READY), .in_A_r(IN0A0R), .in_A_i(IN0A0I), .out_Q_r(
        OUT0Q0R), .out_Q_i(OUT0Q0I), .out_R_r(OUT0R0R), .out_R_i({
        OUT0R0I[47:12], SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11}) );
endmodule

