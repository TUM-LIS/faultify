
module c432 ( N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, 
        N43, N47, N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, 
        N89, N92, N95, N99, N102, N105, N108, N112, N115, N223, N329, N370, 
        N421, N430, N431, N432 );
  input N1, N4, N8, N11, N14, N17, N21, N24, N27, N30, N34, N37, N40, N43, N47,
         N50, N53, N56, N60, N63, N66, N69, N73, N76, N79, N82, N86, N89, N92,
         N95, N99, N102, N105, N108, N112, N115;
  output N223, N329, N370, N421, N430, N431, N432;
  wire   n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204;

  AO21X1 U111 ( .IN1(n110), .IN2(n111), .IN3(n112), .Q(N432) );
  INVX0 U112 ( .INP(n113), .ZN(n112) );
  AO221X1 U113 ( .IN1(n114), .IN2(n115), .IN3(n116), .IN4(n117), .IN5(n118), 
        .Q(n110) );
  INVX0 U114 ( .INP(n119), .ZN(n118) );
  INVX0 U115 ( .INP(n120), .ZN(n116) );
  NAND3X0 U116 ( .IN1(n113), .IN2(n111), .IN3(n121), .QN(N431) );
  NAND3X0 U117 ( .IN1(n119), .IN2(n117), .IN3(n122), .QN(n121) );
  NOR2X0 U118 ( .IN1(n123), .IN2(n124), .QN(N421) );
  OA221X1 U119 ( .IN1(n125), .IN2(n126), .IN3(n127), .IN4(n128), .IN5(n129), 
        .Q(n124) );
  INVX0 U120 ( .INP(N370), .ZN(n125) );
  NOR4X0 U121 ( .IN1(N108), .IN2(N430), .IN3(n114), .IN4(n122), .QN(n123) );
  NAND2X0 U122 ( .IN1(n120), .IN2(n115), .QN(n122) );
  AO222X1 U123 ( .IN1(N86), .IN2(N329), .IN3(n130), .IN4(n131), .IN5(N92), 
        .IN6(N370), .Q(n115) );
  NAND2X0 U124 ( .IN1(N82), .IN2(n132), .QN(n130) );
  AO221X1 U125 ( .IN1(N73), .IN2(N329), .IN3(N79), .IN4(N370), .IN5(n133), .Q(
        n120) );
  AOI222X1 U126 ( .IN1(n134), .IN2(n135), .IN3(N99), .IN4(N329), .IN5(N105), 
        .IN6(N370), .QN(n114) );
  NAND2X0 U127 ( .IN1(N95), .IN2(n132), .QN(n135) );
  NAND4X0 U128 ( .IN1(n119), .IN2(n117), .IN3(n113), .IN4(n111), .QN(N430) );
  AO221X1 U129 ( .IN1(N34), .IN2(N329), .IN3(N40), .IN4(N370), .IN5(n136), .Q(
        n111) );
  AO222X1 U130 ( .IN1(N21), .IN2(N329), .IN3(n137), .IN4(n138), .IN5(N27), 
        .IN6(N370), .Q(n113) );
  NAND2X0 U131 ( .IN1(N17), .IN2(n132), .QN(n137) );
  AO221X1 U132 ( .IN1(N60), .IN2(N329), .IN3(N66), .IN4(N370), .IN5(n139), .Q(
        n117) );
  AO222X1 U133 ( .IN1(N47), .IN2(N329), .IN3(n140), .IN4(n141), .IN5(N53), 
        .IN6(N370), .Q(n119) );
  NAND2X0 U134 ( .IN1(N43), .IN2(n132), .QN(n140) );
  NAND4X0 U135 ( .IN1(n142), .IN2(n143), .IN3(n144), .IN4(n145), .QN(N370) );
  AND4X1 U136 ( .IN1(n146), .IN2(n147), .IN3(n148), .IN4(n149), .Q(n145) );
  OR4X1 U137 ( .IN1(n150), .IN2(n151), .IN3(N115), .IN4(n152), .Q(n149) );
  INVX0 U138 ( .INP(n153), .ZN(n152) );
  NOR2X0 U139 ( .IN1(n127), .IN2(n154), .QN(n150) );
  NAND3X0 U140 ( .IN1(n155), .IN2(n156), .IN3(n157), .QN(n148) );
  INVX0 U141 ( .INP(N105), .ZN(n156) );
  NAND2X0 U142 ( .IN1(N329), .IN2(n158), .QN(n155) );
  NAND3X0 U143 ( .IN1(n159), .IN2(n160), .IN3(n161), .QN(n147) );
  INVX0 U144 ( .INP(N92), .ZN(n160) );
  NAND2X0 U145 ( .IN1(N329), .IN2(n162), .QN(n159) );
  OR3X1 U146 ( .IN1(n163), .IN2(N40), .IN3(n136), .Q(n146) );
  NOR2X0 U147 ( .IN1(n127), .IN2(n164), .QN(n163) );
  AOI222X1 U148 ( .IN1(n165), .IN2(n166), .IN3(n167), .IN4(n168), .IN5(n169), 
        .IN6(n170), .QN(n144) );
  INVX0 U149 ( .INP(n139), .ZN(n170) );
  OA21X1 U150 ( .IN1(n171), .IN2(n127), .IN3(n172), .Q(n169) );
  INVX0 U151 ( .INP(N66), .ZN(n172) );
  INVX0 U152 ( .INP(n133), .ZN(n168) );
  AOI21X1 U153 ( .IN1(n173), .IN2(N329), .IN3(N79), .QN(n167) );
  OA21X1 U154 ( .IN1(n174), .IN2(n127), .IN3(n175), .Q(n165) );
  INVX0 U155 ( .INP(N27), .ZN(n175) );
  NAND3X0 U156 ( .IN1(n176), .IN2(n177), .IN3(n178), .QN(n143) );
  INVX0 U157 ( .INP(N53), .ZN(n177) );
  OR2X1 U158 ( .IN1(n127), .IN2(n179), .Q(n176) );
  NAND3X0 U159 ( .IN1(n180), .IN2(n126), .IN3(n129), .QN(n142) );
  INVX0 U160 ( .INP(N14), .ZN(n126) );
  NAND2X0 U161 ( .IN1(N329), .IN2(n181), .QN(n180) );
  INVX0 U162 ( .INP(n127), .ZN(N329) );
  NOR4X0 U163 ( .IN1(n182), .IN2(n164), .IN3(n183), .IN4(n184), .QN(n127) );
  NAND4X0 U164 ( .IN1(n185), .IN2(n173), .IN3(n162), .IN4(n158), .QN(n184) );
  NAND2X0 U165 ( .IN1(n157), .IN2(n186), .QN(n158) );
  INVX0 U166 ( .INP(N99), .ZN(n186) );
  OA21X1 U167 ( .IN1(n132), .IN2(n187), .IN3(N95), .Q(n157) );
  NAND2X0 U168 ( .IN1(n161), .IN2(n188), .QN(n162) );
  INVX0 U169 ( .INP(N86), .ZN(n188) );
  AOI21X1 U170 ( .IN1(N223), .IN2(n131), .IN3(n189), .QN(n161) );
  OR2X1 U171 ( .IN1(n133), .IN2(N73), .Q(n173) );
  AO21X1 U172 ( .IN1(N63), .IN2(N223), .IN3(n190), .Q(n133) );
  NAND3X0 U173 ( .IN1(n153), .IN2(n154), .IN3(N108), .QN(n185) );
  INVX0 U174 ( .INP(N112), .ZN(n154) );
  NAND2X0 U175 ( .IN1(N102), .IN2(N223), .QN(n153) );
  OR3X1 U176 ( .IN1(n171), .IN2(n179), .IN3(n174), .Q(n183) );
  NOR2X0 U177 ( .IN1(n191), .IN2(N21), .QN(n174) );
  INVX0 U178 ( .INP(n166), .ZN(n191) );
  OA21X1 U179 ( .IN1(n132), .IN2(n192), .IN3(N17), .Q(n166) );
  NOR2X0 U180 ( .IN1(n193), .IN2(N47), .QN(n179) );
  INVX0 U181 ( .INP(n178), .ZN(n193) );
  OA21X1 U182 ( .IN1(n132), .IN2(n194), .IN3(N43), .Q(n178) );
  INVX0 U183 ( .INP(N223), .ZN(n132) );
  NOR2X0 U184 ( .IN1(n139), .IN2(N60), .QN(n171) );
  AO21X1 U185 ( .IN1(N50), .IN2(N223), .IN3(n195), .Q(n139) );
  NOR2X0 U186 ( .IN1(n136), .IN2(N34), .QN(n164) );
  AO21X1 U187 ( .IN1(N24), .IN2(N223), .IN3(n196), .Q(n136) );
  INVX0 U188 ( .INP(n181), .ZN(n182) );
  NAND2X0 U189 ( .IN1(n129), .IN2(n128), .QN(n181) );
  INVX0 U190 ( .INP(N8), .ZN(n128) );
  AOI21X1 U191 ( .IN1(N1), .IN2(N223), .IN3(n197), .QN(n129) );
  NAND4X0 U192 ( .IN1(n198), .IN2(n131), .IN3(n199), .IN4(n200), .QN(N223) );
  OA221X1 U193 ( .IN1(N24), .IN2(n196), .IN3(N102), .IN4(n151), .IN5(n201), 
        .Q(n200) );
  OA22X1 U194 ( .IN1(N50), .IN2(n195), .IN3(N63), .IN4(n190), .Q(n201) );
  INVX0 U195 ( .INP(N69), .ZN(n190) );
  INVX0 U196 ( .INP(N56), .ZN(n195) );
  INVX0 U197 ( .INP(N108), .ZN(n151) );
  INVX0 U198 ( .INP(N30), .ZN(n196) );
  NOR3X0 U199 ( .IN1(n187), .IN2(n192), .IN3(n194), .QN(n199) );
  INVX0 U200 ( .INP(n141), .ZN(n194) );
  NAND2X0 U201 ( .IN1(n202), .IN2(N43), .QN(n141) );
  INVX0 U202 ( .INP(N37), .ZN(n202) );
  INVX0 U203 ( .INP(n138), .ZN(n192) );
  NAND2X0 U204 ( .IN1(n203), .IN2(N17), .QN(n138) );
  INVX0 U205 ( .INP(N11), .ZN(n203) );
  INVX0 U206 ( .INP(n134), .ZN(n187) );
  NAND2X0 U207 ( .IN1(n204), .IN2(N95), .QN(n134) );
  INVX0 U208 ( .INP(N89), .ZN(n204) );
  OR2X1 U209 ( .IN1(N76), .IN2(n189), .Q(n131) );
  INVX0 U210 ( .INP(N82), .ZN(n189) );
  OR2X1 U211 ( .IN1(n197), .IN2(N1), .Q(n198) );
  INVX0 U212 ( .INP(N4), .ZN(n197) );
endmodule

