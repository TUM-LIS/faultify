`timescale 100 ps/100 ps
module circuit_under_test (
clk,
rst,
testVector,
resultVector,
injectionVector
);
input clk;
input rst;
input[69:0] testVector;
output[40:0] resultVector;
input[620:0] injectionVector;
fpu_inj toplevel_instance (
.opa_i(testVector [31:0]),
.opb_i(testVector [63:32]),
.fpu_op_i(testVector [66:64]),
.rmode_i(testVector [68:67]),
.output_o(resultVector [31:0]),
.clk_i(clk),
.start_i(testVector[69]),
.ready_o(resultVector[32]),
.ine_o(resultVector[33]),
.overflow_o(resultVector[34]),
.underflow_o(resultVector[35]),
.div_zero_o(resultVector[36]),
.inf_o(resultVector[37]),
.zero_o(resultVector[38]),
.qnan_o(resultVector[39]),
.snan_o(resultVector[40]),
.p_desc364_p_O_DFFX1pre_norm_mul_(injectionVector[0]),
.p_desc365_p_O_DFFX1pre_norm_mul_(injectionVector[1]),
.p_desc366_p_O_DFFX1pre_norm_mul_(injectionVector[2]),
.p_desc367_p_O_DFFX1pre_norm_mul_(injectionVector[3]),
.p_desc368_p_O_DFFX1pre_norm_mul_(injectionVector[4]),
.p_desc369_p_O_DFFX1pre_norm_mul_(injectionVector[5]),
.p_desc370_p_O_DFFX1pre_norm_mul_(injectionVector[6]),
.p_desc371_p_O_DFFX1pre_norm_mul_(injectionVector[7]),
.p_desc372_p_O_DFFX1pre_norm_mul_(injectionVector[8]),
.p_desc373_p_O_DFFX1pre_norm_mul_(injectionVector[9]),
.p_desc375_p_O_DFFX1mul_24_(injectionVector[10]),
.p_desc376_p_O_DFFX1mul_24_(injectionVector[11]),
.p_desc377_p_O_DFFX1mul_24_(injectionVector[12]),
.p_desc378_p_O_DFFX1mul_24_(injectionVector[13]),
.p_desc379_p_O_DFFX1mul_24_(injectionVector[14]),
.p_desc380_p_O_DFFX1mul_24_(injectionVector[15]),
.p_desc381_p_O_DFFX1mul_24_(injectionVector[16]),
.p_desc382_p_O_DFFX1mul_24_(injectionVector[17]),
.p_desc383_p_O_DFFX1mul_24_(injectionVector[18]),
.p_desc384_p_O_DFFX1mul_24_(injectionVector[19]),
.p_desc385_p_O_DFFX1mul_24_(injectionVector[20]),
.p_desc386_p_O_DFFX1mul_24_(injectionVector[21]),
.p_desc387_p_O_DFFX1mul_24_(injectionVector[22]),
.p_desc388_p_O_DFFX1mul_24_(injectionVector[23]),
.p_desc389_p_O_DFFX1mul_24_(injectionVector[24]),
.p_desc390_p_O_DFFX1mul_24_(injectionVector[25]),
.p_desc391_p_O_DFFX1mul_24_(injectionVector[26]),
.p_desc392_p_O_DFFX1mul_24_(injectionVector[27]),
.p_desc393_p_O_DFFX1mul_24_(injectionVector[28]),
.p_desc394_p_O_DFFX1mul_24_(injectionVector[29]),
.p_desc395_p_O_DFFX1mul_24_(injectionVector[30]),
.p_desc396_p_O_DFFX1mul_24_(injectionVector[31]),
.p_desc397_p_O_DFFX1mul_24_(injectionVector[32]),
.p_desc398_p_O_DFFX1mul_24_(injectionVector[33]),
.p_desc399_p_O_DFFX1mul_24_(injectionVector[34]),
.p_desc400_p_O_DFFX1mul_24_(injectionVector[35]),
.p_desc401_p_O_DFFX1mul_24_(injectionVector[36]),
.p_desc402_p_O_DFFX1mul_24_(injectionVector[37]),
.p_desc403_p_O_DFFX1mul_24_(injectionVector[38]),
.p_desc404_p_O_DFFX1mul_24_(injectionVector[39]),
.p_desc405_p_O_DFFX1mul_24_(injectionVector[40]),
.p_desc406_p_O_DFFX1mul_24_(injectionVector[41]),
.p_desc407_p_O_DFFX1mul_24_(injectionVector[42]),
.p_desc408_p_O_DFFX1mul_24_(injectionVector[43]),
.p_desc409_p_O_DFFX1mul_24_(injectionVector[44]),
.p_desc410_p_O_DFFX1mul_24_(injectionVector[45]),
.p_desc411_p_O_DFFX1mul_24_(injectionVector[46]),
.p_desc412_p_O_DFFX1mul_24_(injectionVector[47]),
.p_desc413_p_O_DFFX1mul_24_(injectionVector[48]),
.p_desc414_p_O_DFFX1mul_24_(injectionVector[49]),
.p_desc415_p_O_DFFX1mul_24_(injectionVector[50]),
.p_desc416_p_O_DFFX1mul_24_(injectionVector[51]),
.p_desc417_p_O_DFFX1mul_24_(injectionVector[52]),
.p_desc418_p_O_DFFX1mul_24_(injectionVector[53]),
.p_desc419_p_O_DFFX1mul_24_(injectionVector[54]),
.p_desc420_p_O_DFFX1mul_24_(injectionVector[55]),
.p_desc421_p_O_DFFX1mul_24_(injectionVector[56]),
.p_desc422_p_O_DFFX1mul_24_(injectionVector[57]),
.p_s_signa_i_reg_p_O_DFFX1mul_24_(injectionVector[58]),
.p_s_signb_i_reg_p_O_DFFX1mul_24_(injectionVector[59]),
.p_s_start_i_reg_p_O_DFFX1mul_24_(injectionVector[60]),
.p_desc423_p_O_DFFX1mul_24_(injectionVector[61]),
.p_s_state_reg_p_O_DFFX1mul_24_(injectionVector[62]),
.p_s_ready_o_reg_p_O_DFFX1mul_24_(injectionVector[63]),
.p_desc424_p_O_DFFX1mul_24_(injectionVector[64]),
.p_desc425_p_O_DFFX1mul_24_(injectionVector[65]),
.p_desc426_p_O_DFFX1mul_24_(injectionVector[66]),
.p_desc427_p_O_DFFX1mul_24_(injectionVector[67]),
.p_desc428_p_O_DFFX1mul_24_(injectionVector[68]),
.p_desc429_p_O_DFFX1mul_24_(injectionVector[69]),
.p_desc430_p_O_DFFX1mul_24_(injectionVector[70]),
.p_desc431_p_O_DFFX1mul_24_(injectionVector[71]),
.p_desc432_p_O_DFFX1mul_24_(injectionVector[72]),
.p_desc433_p_O_DFFX1mul_24_(injectionVector[73]),
.p_desc434_p_O_DFFX1mul_24_(injectionVector[74]),
.p_desc435_p_O_DFFX1mul_24_(injectionVector[75]),
.p_desc436_p_O_DFFX1mul_24_(injectionVector[76]),
.p_desc437_p_O_DFFX1mul_24_(injectionVector[77]),
.p_desc438_p_O_DFFX1mul_24_(injectionVector[78]),
.p_desc439_p_O_DFFX1mul_24_(injectionVector[79]),
.p_desc440_p_O_DFFX1mul_24_(injectionVector[80]),
.p_desc441_p_O_DFFX1mul_24_(injectionVector[81]),
.p_desc442_p_O_DFFX1mul_24_(injectionVector[82]),
.p_desc443_p_O_DFFX1mul_24_(injectionVector[83]),
.p_desc444_p_O_DFFX1mul_24_(injectionVector[84]),
.p_desc445_p_O_DFFX1mul_24_(injectionVector[85]),
.p_desc446_p_O_DFFX1mul_24_(injectionVector[86]),
.p_desc447_p_O_DFFX1mul_24_(injectionVector[87]),
.p_desc448_p_O_DFFX1mul_24_(injectionVector[88]),
.p_desc449_p_O_DFFX1mul_24_(injectionVector[89]),
.p_desc450_p_O_DFFX1mul_24_(injectionVector[90]),
.p_desc451_p_O_DFFX1mul_24_(injectionVector[91]),
.p_desc452_p_O_DFFX1mul_24_(injectionVector[92]),
.p_desc453_p_O_DFFX1mul_24_(injectionVector[93]),
.p_desc454_p_O_DFFX1mul_24_(injectionVector[94]),
.p_desc455_p_O_DFFX1mul_24_(injectionVector[95]),
.p_desc456_p_O_DFFX1mul_24_(injectionVector[96]),
.p_desc457_p_O_DFFX1mul_24_(injectionVector[97]),
.p_desc458_p_O_DFFX1mul_24_(injectionVector[98]),
.p_desc459_p_O_DFFX1mul_24_(injectionVector[99]),
.p_desc460_p_O_DFFX1mul_24_(injectionVector[100]),
.p_desc461_p_O_DFFX1mul_24_(injectionVector[101]),
.p_desc462_p_O_DFFX1mul_24_(injectionVector[102]),
.p_desc463_p_O_DFFX1mul_24_(injectionVector[103]),
.p_desc464_p_O_DFFX1mul_24_(injectionVector[104]),
.p_desc465_p_O_DFFX1mul_24_(injectionVector[105]),
.p_desc466_p_O_DFFX1mul_24_(injectionVector[106]),
.p_desc467_p_O_DFFX1mul_24_(injectionVector[107]),
.p_desc468_p_O_DFFX1mul_24_(injectionVector[108]),
.p_desc469_p_O_DFFX1mul_24_(injectionVector[109]),
.p_desc470_p_O_DFFX1mul_24_(injectionVector[110]),
.p_desc471_p_O_DFFX1mul_24_(injectionVector[111]),
.p_desc472_p_O_DFFX1mul_24_(injectionVector[112]),
.p_desc473_p_O_DFFX1mul_24_(injectionVector[113]),
.p_desc474_p_O_DFFX1mul_24_(injectionVector[114]),
.p_desc475_p_O_DFFX1mul_24_(injectionVector[115]),
.p_desc476_p_O_DFFX1mul_24_(injectionVector[116]),
.p_desc477_p_O_DFFX1mul_24_(injectionVector[117]),
.p_desc478_p_O_DFFX1mul_24_(injectionVector[118]),
.p_desc479_p_O_DFFX1mul_24_(injectionVector[119]),
.p_desc480_p_O_DFFX1mul_24_(injectionVector[120]),
.p_desc481_p_O_DFFX1mul_24_(injectionVector[121]),
.p_desc482_p_O_DFFX1mul_24_(injectionVector[122]),
.p_desc483_p_O_DFFX1mul_24_(injectionVector[123]),
.p_desc484_p_O_DFFX1mul_24_(injectionVector[124]),
.p_desc485_p_O_DFFX1mul_24_(injectionVector[125]),
.p_desc486_p_O_DFFX1mul_24_(injectionVector[126]),
.p_desc487_p_O_DFFX1mul_24_(injectionVector[127]),
.p_desc488_p_O_DFFX1mul_24_(injectionVector[128]),
.p_desc489_p_O_DFFX1mul_24_(injectionVector[129]),
.p_desc490_p_O_DFFX1mul_24_(injectionVector[130]),
.p_desc491_p_O_DFFX1mul_24_(injectionVector[131]),
.p_desc492_p_O_DFFX1mul_24_(injectionVector[132]),
.p_desc493_p_O_DFFX1mul_24_(injectionVector[133]),
.p_desc494_p_O_DFFX1mul_24_(injectionVector[134]),
.p_desc495_p_O_DFFX1mul_24_(injectionVector[135]),
.p_desc496_p_O_DFFX1mul_24_(injectionVector[136]),
.p_desc497_p_O_DFFX1mul_24_(injectionVector[137]),
.p_desc498_p_O_DFFX1mul_24_(injectionVector[138]),
.p_desc499_p_O_DFFX1mul_24_(injectionVector[139]),
.p_desc500_p_O_DFFX1mul_24_(injectionVector[140]),
.p_desc501_p_O_DFFX1mul_24_(injectionVector[141]),
.p_desc502_p_O_DFFX1mul_24_(injectionVector[142]),
.p_desc503_p_O_DFFX1mul_24_(injectionVector[143]),
.p_desc504_p_O_DFFX1mul_24_(injectionVector[144]),
.p_desc505_p_O_DFFX1mul_24_(injectionVector[145]),
.p_desc506_p_O_DFFX1mul_24_(injectionVector[146]),
.p_desc507_p_O_DFFX1mul_24_(injectionVector[147]),
.p_desc508_p_O_DFFX1mul_24_(injectionVector[148]),
.p_desc509_p_O_DFFX1mul_24_(injectionVector[149]),
.p_desc510_p_O_DFFX1mul_24_(injectionVector[150]),
.p_desc511_p_O_DFFX1mul_24_(injectionVector[151]),
.p_desc512_p_O_DFFX1mul_24_(injectionVector[152]),
.p_desc513_p_O_DFFX1mul_24_(injectionVector[153]),
.p_desc514_p_O_DFFX1mul_24_(injectionVector[154]),
.p_desc515_p_O_DFFX1mul_24_(injectionVector[155]),
.p_desc516_p_O_DFFX1mul_24_(injectionVector[156]),
.p_desc517_p_O_DFFX1mul_24_(injectionVector[157]),
.p_desc518_p_O_DFFX1mul_24_(injectionVector[158]),
.p_desc519_p_O_DFFX1mul_24_(injectionVector[159]),
.p_desc520_p_O_DFFX1mul_24_(injectionVector[160]),
.p_desc521_p_O_DFFX1mul_24_(injectionVector[161]),
.p_desc522_p_O_DFFX1mul_24_(injectionVector[162]),
.p_desc523_p_O_DFFX1mul_24_(injectionVector[163]),
.p_desc524_p_O_DFFX1mul_24_(injectionVector[164]),
.p_desc525_p_O_DFFX1mul_24_(injectionVector[165]),
.p_desc526_p_O_DFFX1mul_24_(injectionVector[166]),
.p_desc527_p_O_DFFX1mul_24_(injectionVector[167]),
.p_desc528_p_O_DFFX1mul_24_(injectionVector[168]),
.p_desc529_p_O_DFFX1mul_24_(injectionVector[169]),
.p_desc530_p_O_DFFX1mul_24_(injectionVector[170]),
.p_desc531_p_O_DFFX1mul_24_(injectionVector[171]),
.p_desc532_p_O_DFFX1mul_24_(injectionVector[172]),
.p_desc533_p_O_DFFX1mul_24_(injectionVector[173]),
.p_desc534_p_O_DFFX1mul_24_(injectionVector[174]),
.p_desc535_p_O_DFFX1mul_24_(injectionVector[175]),
.p_desc536_p_O_DFFX1mul_24_(injectionVector[176]),
.p_desc537_p_O_DFFX1mul_24_(injectionVector[177]),
.p_desc538_p_O_DFFX1mul_24_(injectionVector[178]),
.p_desc539_p_O_DFFX1mul_24_(injectionVector[179]),
.p_desc540_p_O_DFFX1mul_24_(injectionVector[180]),
.p_desc541_p_O_DFFX1mul_24_(injectionVector[181]),
.p_desc542_p_O_DFFX1mul_24_(injectionVector[182]),
.p_desc543_p_O_DFFX1mul_24_(injectionVector[183]),
.p_desc544_p_O_DFFX1mul_24_(injectionVector[184]),
.p_desc545_p_O_DFFX1mul_24_(injectionVector[185]),
.p_desc546_p_O_DFFX1mul_24_(injectionVector[186]),
.p_desc547_p_O_DFFX1mul_24_(injectionVector[187]),
.p_desc548_p_O_DFFX1mul_24_(injectionVector[188]),
.p_desc549_p_O_DFFX1mul_24_(injectionVector[189]),
.p_desc550_p_O_DFFX1mul_24_(injectionVector[190]),
.p_desc551_p_O_DFFX1mul_24_(injectionVector[191]),
.p_desc552_p_O_DFFX1mul_24_(injectionVector[192]),
.p_desc553_p_O_DFFX1mul_24_(injectionVector[193]),
.p_desc554_p_O_DFFX1mul_24_(injectionVector[194]),
.p_desc555_p_O_DFFX1mul_24_(injectionVector[195]),
.p_desc556_p_O_DFFX1mul_24_(injectionVector[196]),
.p_desc557_p_O_DFFX1mul_24_(injectionVector[197]),
.p_desc558_p_O_DFFX1mul_24_(injectionVector[198]),
.p_desc559_p_O_DFFX1mul_24_(injectionVector[199]),
.p_desc560_p_O_DFFX1mul_24_(injectionVector[200]),
.p_desc561_p_O_DFFX1mul_24_(injectionVector[201]),
.p_desc562_p_O_DFFX1mul_24_(injectionVector[202]),
.p_desc563_p_O_DFFX1mul_24_(injectionVector[203]),
.p_desc564_p_O_DFFX1mul_24_(injectionVector[204]),
.p_desc565_p_O_DFFX1mul_24_(injectionVector[205]),
.p_desc566_p_O_DFFX1mul_24_(injectionVector[206]),
.p_desc567_p_O_DFFX1mul_24_(injectionVector[207]),
.p_desc568_p_O_DFFX1mul_24_(injectionVector[208]),
.p_desc569_p_O_DFFX1mul_24_(injectionVector[209]),
.p_desc570_p_O_DFFX1mul_24_(injectionVector[210]),
.p_desc571_p_O_DFFX1mul_24_(injectionVector[211]),
.p_desc572_p_O_DFFX1mul_24_(injectionVector[212]),
.p_desc573_p_O_DFFX1mul_24_(injectionVector[213]),
.p_desc574_p_O_DFFX1mul_24_(injectionVector[214]),
.p_desc575_p_O_DFFX1mul_24_(injectionVector[215]),
.p_desc576_p_O_DFFX1mul_24_(injectionVector[216]),
.p_desc577_p_O_DFFX1mul_24_(injectionVector[217]),
.p_desc578_p_O_DFFX1mul_24_(injectionVector[218]),
.p_desc579_p_O_DFFX1mul_24_(injectionVector[219]),
.p_desc580_p_O_DFFX1mul_24_(injectionVector[220]),
.p_desc581_p_O_DFFX1mul_24_(injectionVector[221]),
.p_desc582_p_O_DFFX1mul_24_(injectionVector[222]),
.p_desc583_p_O_DFFX1mul_24_(injectionVector[223]),
.p_desc584_p_O_DFFX1mul_24_(injectionVector[224]),
.p_desc585_p_O_DFFX1mul_24_(injectionVector[225]),
.p_desc586_p_O_DFFX1mul_24_(injectionVector[226]),
.p_desc587_p_O_DFFX1mul_24_(injectionVector[227]),
.p_desc588_p_O_DFFX1mul_24_(injectionVector[228]),
.p_desc589_p_O_DFFX1mul_24_(injectionVector[229]),
.p_desc590_p_O_DFFX1mul_24_(injectionVector[230]),
.p_desc591_p_O_DFFX1mul_24_(injectionVector[231]),
.p_desc592_p_O_DFFX1mul_24_(injectionVector[232]),
.p_desc593_p_O_DFFX1mul_24_(injectionVector[233]),
.p_desc594_p_O_DFFX1mul_24_(injectionVector[234]),
.p_desc595_p_O_DFFX1mul_24_(injectionVector[235]),
.p_desc596_p_O_DFFX1mul_24_(injectionVector[236]),
.p_desc597_p_O_DFFX1mul_24_(injectionVector[237]),
.p_desc598_p_O_DFFX1mul_24_(injectionVector[238]),
.p_desc599_p_O_DFFX1mul_24_(injectionVector[239]),
.p_desc600_p_O_DFFX1mul_24_(injectionVector[240]),
.p_desc601_p_O_DFFX1mul_24_(injectionVector[241]),
.p_desc602_p_O_DFFX1mul_24_(injectionVector[242]),
.p_desc603_p_O_DFFX1mul_24_(injectionVector[243]),
.p_desc604_p_O_DFFX1mul_24_(injectionVector[244]),
.p_desc605_p_O_DFFX1mul_24_(injectionVector[245]),
.p_desc606_p_O_DFFX1mul_24_(injectionVector[246]),
.p_desc607_p_O_DFFX1mul_24_(injectionVector[247]),
.p_desc608_p_O_DFFX1mul_24_(injectionVector[248]),
.p_desc609_p_O_DFFX1mul_24_(injectionVector[249]),
.p_desc610_p_O_DFFX1mul_24_(injectionVector[250]),
.p_desc611_p_O_DFFX1mul_24_(injectionVector[251]),
.p_desc612_p_O_DFFX1mul_24_(injectionVector[252]),
.p_desc613_p_O_DFFX1mul_24_(injectionVector[253]),
.p_desc614_p_O_DFFX1mul_24_(injectionVector[254]),
.p_desc615_p_O_DFFX1mul_24_(injectionVector[255]),
.p_desc616_p_O_DFFX1mul_24_(injectionVector[256]),
.p_desc617_p_O_DFFX1mul_24_(injectionVector[257]),
.p_desc618_p_O_DFFX1mul_24_(injectionVector[258]),
.p_desc619_p_O_DFFX1mul_24_(injectionVector[259]),
.p_desc620_p_O_DFFX1mul_24_(injectionVector[260]),
.p_desc621_p_O_DFFX1mul_24_(injectionVector[261]),
.p_desc622_p_O_DFFX1mul_24_(injectionVector[262]),
.p_desc623_p_O_DFFX1mul_24_(injectionVector[263]),
.p_desc624_p_O_DFFX1mul_24_(injectionVector[264]),
.p_desc625_p_O_DFFX1mul_24_(injectionVector[265]),
.p_desc626_p_O_DFFX1mul_24_(injectionVector[266]),
.p_desc627_p_O_DFFX1mul_24_(injectionVector[267]),
.p_desc628_p_O_DFFX1mul_24_(injectionVector[268]),
.p_desc629_p_O_DFFX1mul_24_(injectionVector[269]),
.p_desc630_p_O_DFFX1mul_24_(injectionVector[270]),
.p_desc631_p_O_DFFX1mul_24_(injectionVector[271]),
.p_desc632_p_O_DFFX1mul_24_(injectionVector[272]),
.p_desc633_p_O_DFFX1mul_24_(injectionVector[273]),
.p_desc634_p_O_DFFX1mul_24_(injectionVector[274]),
.p_desc635_p_O_DFFX1mul_24_(injectionVector[275]),
.p_desc636_p_O_DFFX1mul_24_(injectionVector[276]),
.p_desc637_p_O_DFFX1mul_24_(injectionVector[277]),
.p_desc638_p_O_DFFX1mul_24_(injectionVector[278]),
.p_desc639_p_O_DFFX1mul_24_(injectionVector[279]),
.p_desc640_p_O_DFFX1mul_24_(injectionVector[280]),
.p_desc641_p_O_DFFX1mul_24_(injectionVector[281]),
.p_desc642_p_O_DFFX1mul_24_(injectionVector[282]),
.p_desc643_p_O_DFFX1mul_24_(injectionVector[283]),
.p_desc644_p_O_DFFX1mul_24_(injectionVector[284]),
.p_desc645_p_O_DFFX1mul_24_(injectionVector[285]),
.p_desc646_p_O_DFFX1mul_24_(injectionVector[286]),
.p_desc647_p_O_DFFX1mul_24_(injectionVector[287]),
.p_desc648_p_O_DFFX1mul_24_(injectionVector[288]),
.p_desc649_p_O_DFFX1mul_24_(injectionVector[289]),
.p_desc650_p_O_DFFX1mul_24_(injectionVector[290]),
.p_desc651_p_O_DFFX1mul_24_(injectionVector[291]),
.p_desc652_p_O_DFFX1mul_24_(injectionVector[292]),
.p_desc653_p_O_DFFX1mul_24_(injectionVector[293]),
.p_desc654_p_O_DFFX1mul_24_(injectionVector[294]),
.p_desc655_p_O_DFFX1mul_24_(injectionVector[295]),
.p_desc656_p_O_DFFX1mul_24_(injectionVector[296]),
.p_desc657_p_O_DFFX1mul_24_(injectionVector[297]),
.p_desc658_p_O_DFFX1mul_24_(injectionVector[298]),
.p_desc659_p_O_DFFX1mul_24_(injectionVector[299]),
.p_desc660_p_O_DFFX1mul_24_(injectionVector[300]),
.p_desc661_p_O_DFFX1mul_24_(injectionVector[301]),
.p_desc662_p_O_DFFX1mul_24_(injectionVector[302]),
.p_desc663_p_O_DFFX1mul_24_(injectionVector[303]),
.p_desc664_p_O_DFFX1mul_24_(injectionVector[304]),
.p_desc665_p_O_DFFX1mul_24_(injectionVector[305]),
.p_desc666_p_O_DFFX1mul_24_(injectionVector[306]),
.p_desc667_p_O_DFFX1mul_24_(injectionVector[307]),
.p_desc668_p_O_DFFX1mul_24_(injectionVector[308]),
.p_desc669_p_O_DFFX1mul_24_(injectionVector[309]),
.p_desc670_p_O_DFFX1mul_24_(injectionVector[310]),
.p_desc671_p_O_DFFX1mul_24_(injectionVector[311]),
.p_desc672_p_O_DFFX1mul_24_(injectionVector[312]),
.p_desc673_p_O_DFFX1mul_24_(injectionVector[313]),
.p_desc674_p_O_DFFX1mul_24_(injectionVector[314]),
.p_desc675_p_O_DFFX1mul_24_(injectionVector[315]),
.p_desc676_p_O_DFFX1mul_24_(injectionVector[316]),
.p_desc677_p_O_DFFX1mul_24_(injectionVector[317]),
.p_desc678_p_O_DFFX1mul_24_(injectionVector[318]),
.p_desc679_p_O_DFFX1mul_24_(injectionVector[319]),
.p_desc680_p_O_DFFX1mul_24_(injectionVector[320]),
.p_desc681_p_O_DFFX1mul_24_(injectionVector[321]),
.p_desc682_p_O_DFFX1mul_24_(injectionVector[322]),
.p_desc683_p_O_DFFX1mul_24_(injectionVector[323]),
.p_desc684_p_O_DFFX1mul_24_(injectionVector[324]),
.p_desc685_p_O_DFFX1mul_24_(injectionVector[325]),
.p_desc686_p_O_DFFX1mul_24_(injectionVector[326]),
.p_desc687_p_O_DFFX1mul_24_(injectionVector[327]),
.p_desc688_p_O_DFFX1mul_24_(injectionVector[328]),
.p_desc689_p_O_DFFX1mul_24_(injectionVector[329]),
.p_desc690_p_O_DFFX1mul_24_(injectionVector[330]),
.p_desc691_p_O_DFFX1mul_24_(injectionVector[331]),
.p_desc692_p_O_DFFX1mul_24_(injectionVector[332]),
.p_desc693_p_O_DFFX1mul_24_(injectionVector[333]),
.p_desc694_p_O_DFFX1mul_24_(injectionVector[334]),
.p_desc695_p_O_DFFX1mul_24_(injectionVector[335]),
.p_desc696_p_O_DFFX1mul_24_(injectionVector[336]),
.p_desc697_p_O_DFFX1mul_24_(injectionVector[337]),
.p_desc698_p_O_DFFX1mul_24_(injectionVector[338]),
.p_desc699_p_O_DFFX1mul_24_(injectionVector[339]),
.p_desc700_p_O_DFFX1mul_24_(injectionVector[340]),
.p_desc701_p_O_DFFX1mul_24_(injectionVector[341]),
.p_desc702_p_O_DFFX1mul_24_(injectionVector[342]),
.p_desc703_p_O_DFFX1mul_24_(injectionVector[343]),
.p_desc704_p_O_DFFX1mul_24_(injectionVector[344]),
.p_desc705_p_O_DFFX1mul_24_(injectionVector[345]),
.p_desc706_p_O_DFFX1mul_24_(injectionVector[346]),
.p_desc707_p_O_DFFX1mul_24_(injectionVector[347]),
.p_desc708_p_O_DFFX1mul_24_(injectionVector[348]),
.p_desc709_p_O_DFFX1mul_24_(injectionVector[349]),
.p_desc710_p_O_DFFX1mul_24_(injectionVector[350]),
.p_desc711_p_O_DFFX1mul_24_(injectionVector[351]),
.p_desc712_p_O_DFFX1mul_24_(injectionVector[352]),
.p_desc713_p_O_DFFX1mul_24_(injectionVector[353]),
.p_desc876_p_O_DFFX1post_norm_mul_(injectionVector[354]),
.p_desc877_p_O_DFFX1post_norm_mul_(injectionVector[355]),
.p_desc878_p_O_DFFX1post_norm_mul_(injectionVector[356]),
.p_desc879_p_O_DFFX1post_norm_mul_(injectionVector[357]),
.p_desc880_p_O_DFFX1post_norm_mul_(injectionVector[358]),
.p_desc881_p_O_DFFX1post_norm_mul_(injectionVector[359]),
.p_desc882_p_O_DFFX1post_norm_mul_(injectionVector[360]),
.p_desc883_p_O_DFFX1post_norm_mul_(injectionVector[361]),
.p_desc884_p_O_DFFX1post_norm_mul_(injectionVector[362]),
.p_desc885_p_O_DFFX1post_norm_mul_(injectionVector[363]),
.p_desc886_p_O_DFFX1post_norm_mul_(injectionVector[364]),
.p_desc887_p_O_DFFX1post_norm_mul_(injectionVector[365]),
.p_desc888_p_O_DFFX1post_norm_mul_(injectionVector[366]),
.p_desc889_p_O_DFFX1post_norm_mul_(injectionVector[367]),
.p_desc890_p_O_DFFX1post_norm_mul_(injectionVector[368]),
.p_desc891_p_O_DFFX1post_norm_mul_(injectionVector[369]),
.p_desc892_p_O_DFFX1post_norm_mul_(injectionVector[370]),
.p_desc893_p_O_DFFX1post_norm_mul_(injectionVector[371]),
.p_desc894_p_O_DFFX1post_norm_mul_(injectionVector[372]),
.p_desc895_p_O_DFFX1post_norm_mul_(injectionVector[373]),
.p_desc896_p_O_DFFX1post_norm_mul_(injectionVector[374]),
.p_desc897_p_O_DFFX1post_norm_mul_(injectionVector[375]),
.p_desc898_p_O_DFFX1post_norm_mul_(injectionVector[376]),
.p_desc899_p_O_DFFX1post_norm_mul_(injectionVector[377]),
.p_desc900_p_O_DFFX1post_norm_mul_(injectionVector[378]),
.p_desc901_p_O_DFFX1post_norm_mul_(injectionVector[379]),
.p_desc902_p_O_DFFX1post_norm_mul_(injectionVector[380]),
.p_desc903_p_O_DFFX1post_norm_mul_(injectionVector[381]),
.p_desc904_p_O_DFFX1post_norm_mul_(injectionVector[382]),
.p_desc905_p_O_DFFX1post_norm_mul_(injectionVector[383]),
.p_desc906_p_O_DFFX1post_norm_mul_(injectionVector[384]),
.p_desc907_p_O_DFFX1post_norm_mul_(injectionVector[385]),
.p_desc908_p_O_DFFX1post_norm_mul_(injectionVector[386]),
.p_desc909_p_O_DFFX1post_norm_mul_(injectionVector[387]),
.p_desc910_p_O_DFFX1post_norm_mul_(injectionVector[388]),
.p_desc911_p_O_DFFX1post_norm_mul_(injectionVector[389]),
.p_desc912_p_O_DFFX1post_norm_mul_(injectionVector[390]),
.p_desc913_p_O_DFFX1post_norm_mul_(injectionVector[391]),
.p_desc914_p_O_DFFX1post_norm_mul_(injectionVector[392]),
.p_desc915_p_O_DFFX1post_norm_mul_(injectionVector[393]),
.p_desc916_p_O_DFFX1post_norm_mul_(injectionVector[394]),
.p_desc917_p_O_DFFX1post_norm_mul_(injectionVector[395]),
.p_desc918_p_O_DFFX1post_norm_mul_(injectionVector[396]),
.p_desc919_p_O_DFFX1post_norm_mul_(injectionVector[397]),
.p_desc920_p_O_DFFX1post_norm_mul_(injectionVector[398]),
.p_desc921_p_O_DFFX1post_norm_mul_(injectionVector[399]),
.p_desc922_p_O_DFFX1post_norm_mul_(injectionVector[400]),
.p_desc923_p_O_DFFX1post_norm_mul_(injectionVector[401]),
.p_desc924_p_O_DFFX1post_norm_mul_(injectionVector[402]),
.p_desc925_p_O_DFFX1post_norm_mul_(injectionVector[403]),
.p_desc926_p_O_DFFX1post_norm_mul_(injectionVector[404]),
.p_desc927_p_O_DFFX1post_norm_mul_(injectionVector[405]),
.p_desc928_p_O_DFFX1post_norm_mul_(injectionVector[406]),
.p_desc929_p_O_DFFX1post_norm_mul_(injectionVector[407]),
.p_desc930_p_O_DFFX1post_norm_mul_(injectionVector[408]),
.p_desc931_p_O_DFFX1post_norm_mul_(injectionVector[409]),
.p_desc932_p_O_DFFX1post_norm_mul_(injectionVector[410]),
.p_desc933_p_O_DFFX1post_norm_mul_(injectionVector[411]),
.p_desc934_p_O_DFFX1post_norm_mul_(injectionVector[412]),
.p_desc935_p_O_DFFX1post_norm_mul_(injectionVector[413]),
.p_desc936_p_O_DFFX1post_norm_mul_(injectionVector[414]),
.p_desc937_p_O_DFFX1post_norm_mul_(injectionVector[415]),
.p_desc938_p_O_DFFX1post_norm_mul_(injectionVector[416]),
.p_desc939_p_O_DFFX1post_norm_mul_(injectionVector[417]),
.p_desc940_p_O_DFFX1post_norm_mul_(injectionVector[418]),
.p_desc941_p_O_DFFX1post_norm_mul_(injectionVector[419]),
.p_desc942_p_O_DFFX1post_norm_mul_(injectionVector[420]),
.p_desc943_p_O_DFFX1post_norm_mul_(injectionVector[421]),
.p_desc944_p_O_DFFX1post_norm_mul_(injectionVector[422]),
.p_desc945_p_O_DFFX1post_norm_mul_(injectionVector[423]),
.p_desc946_p_O_DFFX1post_norm_mul_(injectionVector[424]),
.p_desc947_p_O_DFFX1post_norm_mul_(injectionVector[425]),
.p_desc948_p_O_DFFX1post_norm_mul_(injectionVector[426]),
.p_desc949_p_O_DFFX1post_norm_mul_(injectionVector[427]),
.p_desc950_p_O_DFFX1post_norm_mul_(injectionVector[428]),
.p_desc951_p_O_DFFX1post_norm_mul_(injectionVector[429]),
.p_desc952_p_O_DFFX1post_norm_mul_(injectionVector[430]),
.p_desc953_p_O_DFFX1post_norm_mul_(injectionVector[431]),
.p_desc954_p_O_DFFX1post_norm_mul_(injectionVector[432]),
.p_desc955_p_O_DFFX1post_norm_mul_(injectionVector[433]),
.p_desc956_p_O_DFFX1post_norm_mul_(injectionVector[434]),
.p_desc957_p_O_DFFX1post_norm_mul_(injectionVector[435]),
.p_desc958_p_O_DFFX1post_norm_mul_(injectionVector[436]),
.p_desc959_p_O_DFFX1post_norm_mul_(injectionVector[437]),
.p_desc960_p_O_DFFX1post_norm_mul_(injectionVector[438]),
.p_desc961_p_O_DFFX1post_norm_mul_(injectionVector[439]),
.p_desc962_p_O_DFFX1post_norm_mul_(injectionVector[440]),
.p_desc963_p_O_DFFX1post_norm_mul_(injectionVector[441]),
.p_desc964_p_O_DFFX1post_norm_mul_(injectionVector[442]),
.p_desc965_p_O_DFFX1post_norm_mul_(injectionVector[443]),
.p_desc966_p_O_DFFX1post_norm_mul_(injectionVector[444]),
.p_desc967_p_O_DFFX1post_norm_mul_(injectionVector[445]),
.p_desc968_p_O_DFFX1post_norm_mul_(injectionVector[446]),
.p_desc969_p_O_DFFX1post_norm_mul_(injectionVector[447]),
.p_desc970_p_O_DFFX1post_norm_mul_(injectionVector[448]),
.p_desc971_p_O_DFFX1post_norm_mul_(injectionVector[449]),
.p_desc972_p_O_DFFX1post_norm_mul_(injectionVector[450]),
.p_desc973_p_O_DFFX1post_norm_mul_(injectionVector[451]),
.p_desc974_p_O_DFFX1post_norm_mul_(injectionVector[452]),
.p_desc975_p_O_DFFX1post_norm_mul_(injectionVector[453]),
.p_desc976_p_O_DFFX1post_norm_mul_(injectionVector[454]),
.p_desc977_p_O_DFFX1post_norm_mul_(injectionVector[455]),
.p_desc978_p_O_DFFX1post_norm_mul_(injectionVector[456]),
.p_desc979_p_O_DFFX1post_norm_mul_(injectionVector[457]),
.p_desc980_p_O_DFFX1post_norm_mul_(injectionVector[458]),
.p_desc981_p_O_DFFX1post_norm_mul_(injectionVector[459]),
.p_desc982_p_O_DFFX1post_norm_mul_(injectionVector[460]),
.p_desc983_p_O_DFFX1post_norm_mul_(injectionVector[461]),
.p_desc984_p_O_DFFX1post_norm_mul_(injectionVector[462]),
.p_desc985_p_O_DFFX1post_norm_mul_(injectionVector[463]),
.p_desc986_p_O_DFFX1post_norm_mul_(injectionVector[464]),
.p_desc987_p_O_DFFX1post_norm_mul_(injectionVector[465]),
.p_desc988_p_O_DFFX1post_norm_mul_(injectionVector[466]),
.p_desc989_p_O_DFFX1post_norm_mul_(injectionVector[467]),
.p_desc990_p_O_DFFX1post_norm_mul_(injectionVector[468]),
.p_desc991_p_O_DFFX1post_norm_mul_(injectionVector[469]),
.p_desc992_p_O_DFFX1post_norm_mul_(injectionVector[470]),
.p_desc993_p_O_DFFX1post_norm_mul_(injectionVector[471]),
.p_desc994_p_O_DFFX1post_norm_mul_(injectionVector[472]),
.p_desc995_p_O_DFFX1post_norm_mul_(injectionVector[473]),
.p_desc996_p_O_DFFX1post_norm_mul_(injectionVector[474]),
.p_desc997_p_O_DFFX1post_norm_mul_(injectionVector[475]),
.p_desc998_p_O_DFFX1post_norm_mul_(injectionVector[476]),
.p_desc999_p_O_DFFX1post_norm_mul_(injectionVector[477]),
.p_desc1000_p_O_DFFX1post_norm_mul_(injectionVector[478]),
.p_s_sign_i_reg_p_O_DFFX1post_norm_mul_(injectionVector[479]),
.p_desc1001_p_O_DFFX1post_norm_mul_(injectionVector[480]),
.p_desc1002_p_O_DFFX1post_norm_mul_(injectionVector[481]),
.p_desc1003_p_O_DFFX1post_norm_mul_(injectionVector[482]),
.p_desc1004_p_O_DFFX1post_norm_mul_(injectionVector[483]),
.p_desc1005_p_O_DFFX1post_norm_mul_(injectionVector[484]),
.p_desc1006_p_O_DFFX1post_norm_mul_(injectionVector[485]),
.p_desc1007_p_O_DFFX1post_norm_mul_(injectionVector[486]),
.p_desc1008_p_O_DFFX1post_norm_mul_(injectionVector[487]),
.p_desc1009_p_O_DFFX1post_norm_mul_(injectionVector[488]),
.p_desc1010_p_O_DFFX1post_norm_mul_(injectionVector[489]),
.p_desc1011_p_O_DFFX1post_norm_mul_(injectionVector[490]),
.p_desc1012_p_O_DFFX1post_norm_mul_(injectionVector[491]),
.p_desc1013_p_O_DFFX1post_norm_mul_(injectionVector[492]),
.p_desc1014_p_O_DFFX1post_norm_mul_(injectionVector[493]),
.p_desc1015_p_O_DFFX1post_norm_mul_(injectionVector[494]),
.p_desc1016_p_O_DFFX1post_norm_mul_(injectionVector[495]),
.p_desc1017_p_O_DFFX1post_norm_mul_(injectionVector[496]),
.p_desc1018_p_O_DFFX1post_norm_mul_(injectionVector[497]),
.p_desc1019_p_O_DFFX1post_norm_mul_(injectionVector[498]),
.p_desc1020_p_O_DFFX1post_norm_mul_(injectionVector[499]),
.p_desc1021_p_O_DFFX1post_norm_mul_(injectionVector[500]),
.p_desc1022_p_O_DFFX1post_norm_mul_(injectionVector[501]),
.p_desc1024_p_O_DFFX1post_norm_mul_(injectionVector[502]),
.p_desc1025_p_O_DFFX1post_norm_mul_(injectionVector[503]),
.p_desc1026_p_O_DFFX1post_norm_mul_(injectionVector[504]),
.p_desc1027_p_O_DFFX1post_norm_mul_(injectionVector[505]),
.p_desc1028_p_O_DFFX1post_norm_mul_(injectionVector[506]),
.p_desc1029_p_O_DFFX1post_norm_mul_(injectionVector[507]),
.p_desc1030_p_O_DFFX1post_norm_mul_(injectionVector[508]),
.p_desc1031_p_O_DFFX1post_norm_mul_(injectionVector[509]),
.p_desc1032_p_O_DFFX1post_norm_mul_(injectionVector[510]),
.p_desc1033_p_O_DFFX1post_norm_mul_(injectionVector[511]),
.p_desc1034_p_O_DFFX1post_norm_mul_(injectionVector[512]),
.p_desc1035_p_O_DFFX1post_norm_mul_(injectionVector[513]),
.p_desc1036_p_O_DFFX1post_norm_mul_(injectionVector[514]),
.p_desc1037_p_O_DFFX1post_norm_mul_(injectionVector[515]),
.p_desc1038_p_O_DFFX1post_norm_mul_(injectionVector[516]),
.p_desc1039_p_O_DFFX1post_norm_mul_(injectionVector[517]),
.p_desc1040_p_O_DFFX1post_norm_mul_(injectionVector[518]),
.p_desc1041_p_O_DFFX1post_norm_mul_(injectionVector[519]),
.p_desc1042_p_O_DFFX1post_norm_mul_(injectionVector[520]),
.p_desc1043_p_O_DFFX1post_norm_mul_(injectionVector[521]),
.p_desc1044_p_O_DFFX1post_norm_mul_(injectionVector[522]),
.p_desc1045_p_O_DFFX1post_norm_mul_(injectionVector[523]),
.p_desc1046_p_O_DFFX1post_norm_mul_(injectionVector[524]),
.p_desc1047_p_O_DFFX1post_norm_mul_(injectionVector[525]),
.p_desc1048_p_O_DFFX1post_norm_mul_(injectionVector[526]),
.p_desc1049_p_O_DFFX1post_norm_mul_(injectionVector[527]),
.p_desc1050_p_O_DFFX1post_norm_mul_(injectionVector[528]),
.p_desc1051_p_O_DFFX1post_norm_mul_(injectionVector[529]),
.p_desc1052_p_O_DFFX1post_norm_mul_(injectionVector[530]),
.p_desc1053_p_O_DFFX1post_norm_mul_(injectionVector[531]),
.p_desc1054_p_O_DFFX1post_norm_mul_(injectionVector[532]),
.p_desc1055_p_O_DFFX1post_norm_mul_(injectionVector[533]),
.p_desc1056_p_O_DFFX1post_norm_mul_(injectionVector[534]),
.p_desc1057_p_O_DFFX1post_norm_mul_(injectionVector[535]),
.p_desc1058_p_O_DFFX1post_norm_mul_(injectionVector[536]),
.p_desc1059_p_O_DFFX1post_norm_mul_(injectionVector[537]),
.p_desc1060_p_O_DFFX1post_norm_mul_(injectionVector[538]),
.p_desc1061_p_O_DFFX1post_norm_mul_(injectionVector[539]),
.p_desc1062_p_O_DFFX1post_norm_mul_(injectionVector[540]),
.p_desc1063_p_O_DFFX1post_norm_mul_(injectionVector[541]),
.p_desc1064_p_O_DFFX1post_norm_mul_(injectionVector[542]),
.p_desc1065_p_O_DFFX1post_norm_mul_(injectionVector[543]),
.p_desc1066_p_O_DFFX1post_norm_mul_(injectionVector[544]),
.p_desc1067_p_O_DFFX1post_norm_mul_(injectionVector[545]),
.p_desc1068_p_O_DFFX1post_norm_mul_(injectionVector[546]),
.p_desc1069_p_O_DFFX1post_norm_mul_(injectionVector[547]),
.p_desc1070_p_O_DFFX1post_norm_mul_(injectionVector[548]),
.p_desc1071_p_O_DFFX1post_norm_mul_(injectionVector[549]),
.p_desc1072_p_O_DFFX1post_norm_mul_(injectionVector[550]),
.p_desc1073_p_O_DFFX1post_norm_mul_(injectionVector[551]),
.p_desc1074_p_O_DFFX1post_norm_mul_(injectionVector[552]),
.p_desc1075_p_O_DFFX1post_norm_mul_(injectionVector[553]),
.p_desc1076_p_O_DFFX1post_norm_mul_(injectionVector[554]),
.p_desc1077_p_O_DFFX1post_norm_mul_(injectionVector[555]),
.p_desc1078_p_O_DFFX1post_norm_mul_(injectionVector[556]),
.p_desc1079_p_O_DFFX1post_norm_mul_(injectionVector[557]),
.p_desc1080_p_O_DFFX1post_norm_mul_(injectionVector[558]),
.p_desc1081_p_O_DFFX1post_norm_mul_(injectionVector[559]),
.p_desc1082_p_O_DFFX1post_norm_mul_(injectionVector[560]),
.p_desc1083_p_O_DFFX1post_norm_mul_(injectionVector[561]),
.p_ine_o_reg_p_O_DFFX1post_norm_mul_(injectionVector[562]),
.p_desc1084_p_O_DFFX1post_norm_mul_(injectionVector[563]),
.p_desc1085_p_O_DFFX1post_norm_mul_(injectionVector[564]),
.p_desc1086_p_O_DFFX1post_norm_mul_(injectionVector[565]),
.p_desc1087_p_O_DFFX1post_norm_mul_(injectionVector[566]),
.p_desc1088_p_O_DFFX1post_norm_mul_(injectionVector[567]),
.p_desc1089_p_O_DFFX1post_norm_mul_(injectionVector[568]),
.p_desc1090_p_O_DFFX1post_norm_mul_(injectionVector[569]),
.p_desc1091_p_O_DFFX1post_norm_mul_(injectionVector[570]),
.p_desc1092_p_O_DFFX1post_norm_mul_(injectionVector[571]),
.p_desc1093_p_O_DFFX1post_norm_mul_(injectionVector[572]),
.p_desc1094_p_O_DFFX1post_norm_mul_(injectionVector[573]),
.p_desc1095_p_O_DFFX1post_norm_mul_(injectionVector[574]),
.p_desc1096_p_O_DFFX1post_norm_mul_(injectionVector[575]),
.p_desc1097_p_O_DFFX1post_norm_mul_(injectionVector[576]),
.p_desc1098_p_O_DFFX1post_norm_mul_(injectionVector[577]),
.p_desc1099_p_O_DFFX1post_norm_mul_(injectionVector[578]),
.p_desc1100_p_O_DFFX1post_norm_mul_(injectionVector[579]),
.p_desc1101_p_O_DFFX1post_norm_mul_(injectionVector[580]),
.p_desc1102_p_O_DFFX1post_norm_mul_(injectionVector[581]),
.p_desc1103_p_O_DFFX1post_norm_mul_(injectionVector[582]),
.p_desc1104_p_O_DFFX1post_norm_mul_(injectionVector[583]),
.p_desc1105_p_O_DFFX1post_norm_mul_(injectionVector[584]),
.p_desc1106_p_O_DFFX1post_norm_mul_(injectionVector[585]),
.p_desc1107_p_O_DFFX1post_norm_mul_(injectionVector[586]),
.p_desc1108_p_O_DFFX1post_norm_mul_(injectionVector[587]),
.p_desc1109_p_O_DFFX1post_norm_mul_(injectionVector[588]),
.p_desc1110_p_O_DFFX1post_norm_mul_(injectionVector[589]),
.p_desc1111_p_O_DFFX1post_norm_mul_(injectionVector[590]),
.p_desc1112_p_O_DFFX1post_norm_mul_(injectionVector[591]),
.p_desc1113_p_O_DFFX1post_norm_mul_(injectionVector[592]),
.p_desc1114_p_O_DFFX1post_norm_mul_(injectionVector[593]),
.p_desc1115_p_O_DFFX1post_norm_mul_(injectionVector[594]),
.p_desc1116_p_O_DFFX1post_norm_mul_(injectionVector[595]),
.p_desc1117_p_O_DFFX1post_norm_mul_(injectionVector[596]),
.p_desc1118_p_O_DFFX1post_norm_mul_(injectionVector[597]),
.p_desc1119_p_O_DFFX1post_norm_mul_(injectionVector[598]),
.p_desc1120_p_O_DFFX1post_norm_mul_(injectionVector[599]),
.p_desc1121_p_O_DFFX1post_norm_mul_(injectionVector[600]),
.p_desc1122_p_O_DFFX1post_norm_mul_(injectionVector[601]),
.p_desc1123_p_O_DFFX1post_norm_mul_(injectionVector[602]),
.p_desc1124_p_O_DFFX1post_norm_mul_(injectionVector[603]),
.p_desc1125_p_O_DFFX1post_norm_mul_(injectionVector[604]),
.p_desc1126_p_O_DFFX1post_norm_mul_(injectionVector[605]),
.p_desc1127_p_O_DFFX1post_norm_mul_(injectionVector[606]),
.p_desc1128_p_O_DFFX1post_norm_mul_(injectionVector[607]),
.p_desc1129_p_O_DFFX1post_norm_mul_(injectionVector[608]),
.p_desc1130_p_O_DFFX1post_norm_mul_(injectionVector[609]),
.p_desc1131_p_O_DFFX1post_norm_mul_(injectionVector[610]),
.p_desc1132_p_O_DFFX1post_norm_mul_(injectionVector[611]),
.p_desc1133_p_O_DFFX1post_norm_mul_(injectionVector[612]),
.p_desc1134_p_O_DFFX1post_norm_mul_(injectionVector[613]),
.p_desc1135_p_O_DFFX1post_norm_mul_(injectionVector[614]),
.p_desc1136_p_O_DFFX1post_norm_mul_(injectionVector[615]),
.p_desc1137_p_O_DFFX1post_norm_mul_(injectionVector[616]),
.p_desc1138_p_O_DFFX1post_norm_mul_(injectionVector[617]),
.p_desc1171_p_O_DFFX1post_norm_mul_(injectionVector[618]),
.p_desc1172_p_O_DFFX1post_norm_mul_(injectionVector[619]),
.p_desc1174_p_O_DFFX1post_norm_mul_(injectionVector[620]));
endmodule